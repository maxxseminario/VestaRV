

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO MCU 
  PIN resetn_in 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 25.842 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 113.749 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6 ; 
    ANTENNAMAXAREACAR 974.013 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4292.32 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.32103 LAYER VIA6 ;
  END resetn_in
  PIN resetn_out 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.474 LAYER M2 ;
  END resetn_out
  PIN resetn_dir 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6365 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8446 LAYER M2 ;
  END resetn_dir
  PIN resetn_ren 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5895 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6378 LAYER M2 ;
  END resetn_ren
  PIN prt1_in[7] 
    ANTENNAPARTIALMETALAREA 15.4155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 67.9162 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2 ; 
    ANTENNAMAXAREACAR 570.452 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2511.78 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.369004 LAYER VIA2 ;
  END prt1_in[7]
  PIN prt1_in[6] 
    ANTENNAPARTIALMETALAREA 22.6125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 99.495 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.962 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.2768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 112.492 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 485.766 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.08401 LAYER VIA3 ;
  END prt1_in[6]
  PIN prt1_in[5] 
    ANTENNAPARTIALMETALAREA 14.0905 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 62.0422 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.706 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.5504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1305 LAYER M3 ; 
    ANTENNAMAXAREACAR 98.311 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 432.269 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.782188 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M4 ;
    ANTENNAGATEAREA 0.2577 LAYER M4 ; 
    ANTENNAMAXAREACAR 99.1725 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 436.23 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.782188 LAYER VIA4 ;
  END prt1_in[5]
  PIN prt1_in[4] 
    ANTENNAPARTIALMETALAREA 4.8725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.439 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.59 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.04 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1305 LAYER M3 ; 
    ANTENNAMAXAREACAR 97.1232 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 427.042 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.782188 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.178 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M4 ;
    ANTENNAGATEAREA 0.1305 LAYER M4 ; 
    ANTENNAMAXAREACAR 98.4872 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 433.381 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAMAXCUTCAR 0.935444 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 6.006 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 26.4704 LAYER M5 ;
    ANTENNAGATEAREA 0.2577 LAYER M5 ; 
    ANTENNAMAXAREACAR 121.793 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 536.099 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.935444 LAYER VIA5 ;
  END prt1_in[4]
  PIN prt1_in[3] 
    ANTENNAPARTIALMETALAREA 0.176 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1936 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4982 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.242 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8422 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 LAYER M4 ; 
    ANTENNAMAXAREACAR 19.556 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 25.0566 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAMAXCUTCAR 0.314465 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.52 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER M5 ;
    ANTENNAGATEAREA 0.318 LAYER M5 ; 
    ANTENNAMAXAREACAR 30.6252 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 45.1069 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.25786 LAYER VIA5 ;
  END prt1_in[3]
  PIN prt1_in[2] 
    ANTENNAPARTIALMETALAREA 2.1135 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3434 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 12.418 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.7712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1931 LAYER M3 ; 
    ANTENNAMAXAREACAR 122.456 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 540.411 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3 ;
  END prt1_in[2]
  PIN prt1_in[1] 
    ANTENNAPARTIALMETALAREA 13.1575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 57.937 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.782 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.0848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3 ; 
    ANTENNAMAXAREACAR 112.431 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 494.435 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3 ;
  END prt1_in[1]
  PIN prt1_in[0] 
    ANTENNAPARTIALMETALAREA 22.0995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 97.2378 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.418 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.4832 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3 ; 
    ANTENNAMAXAREACAR 52.3228 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 229.855 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3 ;
  END prt1_in[0]
  PIN prt1_out[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2 ;
  END prt1_out[7]
  PIN prt1_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.499 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 55.0836 LAYER M2 ;
  END prt1_out[6]
  PIN prt1_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[5]
  PIN prt1_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[4]
  PIN prt1_out[3] 
    ANTENNAPARTIALMETALAREA 1.796 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9024 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.186 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.0624 LAYER M3 ;
  END prt1_out[3]
  PIN prt1_out[2] 
    ANTENNAPARTIALMETALAREA 0.092 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.804 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.8256 LAYER M3 ;
  END prt1_out[2]
  PIN prt1_out[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 64.042 LAYER M2 ;
  END prt1_out[1]
  PIN prt1_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 51.018 LAYER M2 ;
  END prt1_out[0]
  PIN prt1_dir[7] 
    ANTENNAPARTIALMETALAREA 3.0115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.2506 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.782 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.6848 LAYER M3 ;
  END prt1_dir[7]
  PIN prt1_dir[6] 
    ANTENNAPARTIALMETALAREA 0.2165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9526 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.266 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2144 LAYER M3 ;
  END prt1_dir[6]
  PIN prt1_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2 ;
  END prt1_dir[5]
  PIN prt1_dir[4] 
    ANTENNAPARTIALMETALAREA 3.3585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.098 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.0752 LAYER M3 ;
  END prt1_dir[4]
  PIN prt1_dir[3] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.064 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.1696 LAYER M3 ;
  END prt1_dir[3]
  PIN prt1_dir[2] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0855 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4202 LAYER M2 ;
  END prt1_dir[2]
  PIN prt1_dir[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[1]
  PIN prt1_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.2345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 53.9198 LAYER M2 ;
  END prt1_dir[0]
  PIN prt1_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0855 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4202 LAYER M2 ;
  END prt1_ren[7]
  PIN prt1_ren[6] 
    ANTENNAPARTIALMETALAREA 1.1805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1942 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.466 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4944 LAYER M3 ;
  END prt1_ren[6]
  PIN prt1_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M2 ;
  END prt1_ren[5]
  PIN prt1_ren[4] 
    ANTENNAPARTIALMETALAREA 3.2985 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.5574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.2368 LAYER M3 ;
  END prt1_ren[4]
  PIN prt1_ren[3] 
    ANTENNAPARTIALMETALAREA 0.2475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.089 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.566 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.7344 LAYER M3 ;
  END prt1_ren[3]
  PIN prt1_ren[2] 
    ANTENNAPARTIALMETALAREA 1.5295 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7738 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.702 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5328 LAYER M3 ;
  END prt1_ren[2]
  PIN prt1_ren[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
  END prt1_ren[1]
  PIN prt1_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.3905 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 54.6062 LAYER M2 ;
  END prt1_ren[0]
  PIN prt2_in[7] 
    ANTENNAPARTIALMETALAREA 0.7785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5134 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0595 LAYER M2 ; 
    ANTENNAMAXAREACAR 18.0714 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 78.4706 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.336134 LAYER VIA2 ;
  END prt2_in[7]
  PIN prt2_in[6] 
    ANTENNAPARTIALMETALAREA 0.7555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4122 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2 ; 
    ANTENNAMAXAREACAR 27.7954 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 121.522 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2 ;
  END prt2_in[6]
  PIN prt2_in[5] 
    ANTENNAPARTIALMETALAREA 0.7125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.135 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 LAYER M2 ; 
    ANTENNAMAXAREACAR 7.72407 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 32.9611 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.185185 LAYER VIA2 ;
  END prt2_in[5]
  PIN prt2_in[4] 
    ANTENNAPARTIALMETALAREA 0.5555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.2368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 146.784 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 630.772 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt2_in[4]
  PIN prt2_in[3] 
    ANTENNAPARTIALMETALAREA 1.234 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5334 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M2 ; 
    ANTENNAMAXAREACAR 6.88784 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 9.43291 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.104822 LAYER VIA2 ;
  END prt2_in[3]
  PIN prt2_in[2] 
    ANTENNAPARTIALMETALAREA 0.6785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9854 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0893 LAYER M2 ; 
    ANTENNAMAXAREACAR 11.5812 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 48.6697 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.223964 LAYER VIA2 ;
  END prt2_in[2]
  PIN prt2_in[1] 
    ANTENNAPARTIALMETALAREA 0.7155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1482 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0893 LAYER M2 ; 
    ANTENNAMAXAREACAR 11.3908 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 48.0739 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.223964 LAYER VIA2 ;
  END prt2_in[1]
  PIN prt2_in[0] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 30.982 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 136.365 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0381 LAYER M3 ; 
    ANTENNAMAXAREACAR 850.332 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3731.77 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.04987 LAYER VIA3 ;
  END prt2_in[0]
  PIN prt2_out[7] 
    ANTENNAPARTIALMETALAREA 0.471 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0724 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.4368 LAYER M3 ;
  END prt2_out[7]
  PIN prt2_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.681 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2 ;
  END prt2_out[6]
  PIN prt2_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.577 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6708 LAYER M2 ;
  END prt2_out[5]
  PIN prt2_out[4] 
    ANTENNAPARTIALMETALAREA 0.679 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9876 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.038 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.2112 LAYER M3 ;
  END prt2_out[4]
  PIN prt2_out[3] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2 ;
  END prt2_out[3]
  PIN prt2_out[2] 
    ANTENNAPARTIALMETALAREA 0.152 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.586 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 59.8224 LAYER M3 ;
  END prt2_out[2]
  PIN prt2_out[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.279 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2276 LAYER M2 ;
  END prt2_out[1]
  PIN prt2_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.512 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M2 ;
  END prt2_out[0]
  PIN prt2_dir[7] 
    ANTENNAPARTIALMETALAREA 0.711 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1284 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.8928 LAYER M3 ;
  END prt2_dir[7]
  PIN prt2_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6554 LAYER M2 ;
  END prt2_dir[6]
  PIN prt2_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6815 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0426 LAYER M2 ;
  END prt2_dir[5]
  PIN prt2_dir[4] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1946 LAYER M2 ;
  END prt2_dir[4]
  PIN prt2_dir[3] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1946 LAYER M2 ;
  END prt2_dir[3]
  PIN prt2_dir[2] 
    ANTENNAPARTIALMETALAREA 0.531 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3364 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.2368 LAYER M3 ;
  END prt2_dir[2]
  PIN prt2_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9018 LAYER M2 ;
  END prt2_dir[1]
  PIN prt2_dir[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2254 LAYER M2 ;
  END prt2_dir[0]
  PIN prt2_ren[7] 
    ANTENNAPARTIALMETALAREA 0.6435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8314 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.878 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.1072 LAYER M3 ;
  END prt2_ren[7]
  PIN prt2_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2714 LAYER M2 ;
  END prt2_ren[6]
  PIN prt2_ren[5] 
    ANTENNAPARTIALMETALAREA 0.7345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2318 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.758 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7792 LAYER M3 ;
  END prt2_ren[5]
  PIN prt2_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.519 LAYER M2 ;
  END prt2_ren[4]
  PIN prt2_ren[3] 
    ANTENNAPARTIALMETALAREA 0.8875 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.905 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.146 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.8864 LAYER M3 ;
  END prt2_ren[3]
  PIN prt2_ren[2] 
    ANTENNAPARTIALMETALAREA 0.667 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9348 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.2095 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.7658 LAYER M3 ;
  END prt2_ren[2]
  PIN prt2_ren[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2855 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3002 LAYER M2 ;
  END prt2_ren[1]
  PIN prt2_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6855 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0602 LAYER M2 ;
  END prt2_ren[0]
  PIN prt3_in[7] 
    ANTENNAPARTIALMETALAREA 18.7995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 82.8058 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2 ; 
    ANTENNAMAXAREACAR 698.801 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3074.69 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.738007 LAYER VIA2 ;
  END prt3_in[7]
  PIN prt3_in[6] 
    ANTENNAPARTIALMETALAREA 15.9905 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 70.4022 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 16.178 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.2272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 610.052 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2670.41 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[6]
  PIN prt3_in[5] 
    ANTENNAPARTIALMETALAREA 7.9325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.903 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 15.938 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 70.1712 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.258 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9792 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 39.3685 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 175.57 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA4 ;
  END prt3_in[5]
  PIN prt3_in[4] 
    ANTENNAPARTIALMETALAREA 0.6325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.783 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.9248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.278 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.622 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.9808 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M5 ; 
    ANTENNAMAXAREACAR 47.4781 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 209.971 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.876988 LAYER VIA5 ;
  END prt3_in[4]
  PIN prt3_in[3] 
    ANTENNAPARTIALMETALAREA 4.7355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.8362 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 18.226 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.2384 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1707 LAYER M3 ; 
    ANTENNAMAXAREACAR 119.268 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 524.402 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA3 ;
  END prt3_in[3]
  PIN prt3_in[2] 
    ANTENNAPARTIALMETALAREA 0.5755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5322 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 16.952 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 74.7648 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 644.59 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2824.86 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[2]
  PIN prt3_in[1] 
    ANTENNAPARTIALMETALAREA 14.5355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 63.9562 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.722 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.8208 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 285.009 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1255.83 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3 ;
  END prt3_in[1]
  PIN prt3_in[0] 
    ANTENNAPARTIALMETALAREA 1.9105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.4502 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.438 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.5712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 294.622 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1280.64 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt3_in[0]
  PIN prt3_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.743 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 64.9572 LAYER M2 ;
  END prt3_out[7]
  PIN prt3_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 6.423 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.3492 LAYER M2 ;
  END prt3_out[6]
  PIN prt3_out[5] 
    ANTENNAPARTIALMETALAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5584 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.766 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.8144 LAYER M3 ;
  END prt3_out[5]
  PIN prt3_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.379 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1556 LAYER M2 ;
  END prt3_out[4]
  PIN prt3_out[3] 
    ANTENNAPARTIALMETALAREA 1.792 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.8848 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.806 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9904 LAYER M3 ;
  END prt3_out[3]
  PIN prt3_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.175 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.458 LAYER M2 ;
  END prt3_out[2]
  PIN prt3_out[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.855 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 56.65 LAYER M2 ;
  END prt3_out[1]
  PIN prt3_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.901 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.2084 LAYER M2 ;
  END prt3_out[0]
  PIN prt3_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.2415 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 62.7066 LAYER M2 ;
  END prt3_dir[7]
  PIN prt3_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.0055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.1562 LAYER M2 ;
  END prt3_dir[6]
  PIN prt3_dir[5] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.186 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M3 ;
  END prt3_dir[5]
  PIN prt3_dir[4] 
    ANTENNAPARTIALMETALAREA 0.4165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8326 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.842 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.3488 LAYER M3 ;
  END prt3_dir[4]
  PIN prt3_dir[3] 
    ANTENNAPARTIALMETALAREA 0.1515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.646 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.4864 LAYER M3 ;
  END prt3_dir[3]
  PIN prt3_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.7345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 60.5198 LAYER M2 ;
  END prt3_dir[2]
  PIN prt3_dir[1] 
    ANTENNAPARTIALMETALAREA 14.0495 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.8618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.646 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8864 LAYER M3 ;
  END prt3_dir[1]
  PIN prt3_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.1345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.8798 LAYER M2 ;
  END prt3_dir[0]
  PIN prt3_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.3255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.7642 LAYER M2 ;
  END prt3_ren[7]
  PIN prt3_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.1075 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.561 LAYER M2 ;
  END prt3_ren[6]
  PIN prt3_ren[5] 
    ANTENNAPARTIALMETALAREA 0.2605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1462 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3 ;
  END prt3_ren[5]
  PIN prt3_ren[4] 
    ANTENNAPARTIALMETALAREA 0.6605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9062 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.77 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0582 LAYER M3 ; 
    ANTENNAMAXAREACAR 258.459 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1136.85 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.687285 LAYER VIA3 ;
  END prt3_ren[4]
  PIN prt3_ren[3] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.9872 LAYER M3 ;
  END prt3_ren[3]
  PIN prt3_ren[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 9.6885 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 42.7614 LAYER M2 ;
  END prt3_ren[2]
  PIN prt3_ren[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.3125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 63.107 LAYER M2 ;
  END prt3_ren[1]
  PIN prt3_ren[0] 
    ANTENNAPARTIALMETALAREA 0.5805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5542 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.118 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M3 ;
  END prt3_ren[0]
  PIN prt4_in[7] 
    ANTENNAPARTIALMETALAREA 1.9555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6042 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 26.828 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 118.131 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 389.192 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1708.37 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3 ;
  END prt4_in[7]
  PIN prt4_in[6] 
    ANTENNAPARTIALMETALAREA 1.8555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1642 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 19.838 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 87.4192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 198.371 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 873.831 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.08401 LAYER VIA3 ;
  END prt4_in[6]
  PIN prt4_in[5] 
    ANTENNAPARTIALMETALAREA 1.6785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3854 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.9056 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 251.47 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1102.34 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.16802 LAYER VIA3 ;
  END prt4_in[5]
  PIN prt4_in[4] 
    ANTENNAPARTIALMETALAREA 1.9755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6922 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.858 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.4192 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1204 LAYER M4 ; 
    ANTENNAMAXAREACAR 63.5979 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 279.093 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.25012 LAYER VIA4 ;
  END prt4_in[4]
  PIN prt4_in[3] 
    ANTENNAPARTIALMETALAREA 6.4505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.4262 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.246 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1456 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.2257 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 66.8666 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.08401 LAYER VIA3 ;
  END prt4_in[3]
  PIN prt4_in[2] 
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.998 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 52.8352 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 6.818 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 30.0432 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 96.3583 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 423.219 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.81869 LAYER VIA4 ;
  END prt4_in[2]
  PIN prt4_in[1] 
    ANTENNAPARTIALMETALAREA 0.731 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 20.818 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.6432 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 6.556 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 28.9344 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0636 LAYER M4 ; 
    ANTENNAMAXAREACAR 126.222 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 557.921 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAMAXCUTCAR 1.41509 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.506 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2704 LAYER M5 ;
    ANTENNAGATEAREA 0.1305 LAYER M5 ; 
    ANTENNAMAXAREACAR 130.099 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 575.319 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.41509 LAYER VIA5 ;
  END prt4_in[1]
  PIN prt4_in[0] 
    ANTENNAPARTIALMETALAREA 0.2725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 27.886 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 122.742 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 1080.52 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4736.44 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt4_in[0]
  PIN prt4_out[7] 
    ANTENNAPARTIALMETALAREA 5.292 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8806 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 82.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.256 LAYER M3 ;
  END prt4_out[7]
  PIN prt4_out[6] 
    ANTENNAPARTIALMETALAREA 10.332 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4246 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.736 LAYER M3 ;
  END prt4_out[6]
  PIN prt4_out[5] 
    ANTENNAPARTIALMETALAREA 0.43 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.473 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 19.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22 LAYER M3 ;
  END prt4_out[5]
  PIN prt4_out[4] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.8902 LAYER M3 ;
  END prt4_out[4]
  PIN prt4_out[3] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.998 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.4352 LAYER M3 ;
  END prt4_out[3]
  PIN prt4_out[2] 
    ANTENNAPARTIALMETALAREA 0.331 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.278 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.8672 LAYER M3 ;
  END prt4_out[2]
  PIN prt4_out[1] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.922 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 74.5008 LAYER M6 ;
  END prt4_out[1]
  PIN prt4_out[0] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
  END prt4_out[0]
  PIN prt4_dir[7] 
    ANTENNAPARTIALMETALAREA 0.2915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.6704 LAYER M3 ;
  END prt4_dir[7]
  PIN prt4_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.3785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5534 LAYER M2 ;
  END prt4_dir[6]
  PIN prt4_dir[5] 
    ANTENNADIFFAREA 1.968 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.5785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4334 LAYER M2 ;
  END prt4_dir[5]
  PIN prt4_dir[4] 
    ANTENNADIFFAREA 1.968 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.6385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0974 LAYER M2 ;
  END prt4_dir[4]
  PIN prt4_dir[3] 
    ANTENNAPARTIALMETALAREA 0.871 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.1088 LAYER M3 ;
  END prt4_dir[3]
  PIN prt4_dir[2] 
    ANTENNAPARTIALMETALAREA 0.511 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2484 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.278 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.4672 LAYER M3 ;
  END prt4_dir[2]
  PIN prt4_dir[1] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 17.122 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 75.3808 LAYER M6 ;
  END prt4_dir[1]
  PIN prt4_dir[0] 
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.386 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 72.1424 LAYER M6 ;
  END prt4_dir[0]
  PIN prt4_ren[7] 
    ANTENNAPARTIALMETALAREA 0.5075 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.233 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 59.4528 LAYER M3 ;
  END prt4_ren[7]
  PIN prt4_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.9475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.257 LAYER M2 ;
  END prt4_ren[6]
  PIN prt4_ren[5] 
    ANTENNAPARTIALMETALAREA 1.2105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3262 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.066 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.1344 LAYER M3 ;
  END prt4_ren[5]
  PIN prt4_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.7055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5482 LAYER M2 ;
  END prt4_ren[4]
  PIN prt4_ren[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.1625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.159 LAYER M2 ;
  END prt4_ren[3]
  PIN prt4_ren[2] 
    ANTENNAPARTIALMETALAREA 0.4435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9514 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.1328 LAYER M3 ;
  END prt4_ren[2]
  PIN prt4_ren[1] 
    ANTENNAPARTIALMETALAREA 0.8035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.342 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 71.9488 LAYER M6 ;
  END prt4_ren[1]
  PIN prt4_ren[0] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 17.146 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 75.4864 LAYER M6 ;
  END prt4_ren[0]
  PIN use_dac_glb_bias 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
  END use_dac_glb_bias
  PIN en_bias_buf 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.246 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M3 ;
  END en_bias_buf
  PIN en_bias_gen 
    ANTENNAPARTIALMETALAREA 0.041 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1804 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.566 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.096 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 26.9104 LAYER M4 ;
  END en_bias_gen
  PIN BIAS_ADJ[5] 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.358 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M3 ;
  END BIAS_ADJ[5]
  PIN BIAS_ADJ[4] 
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.438 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7712 LAYER M4 ;
  END BIAS_ADJ[4]
  PIN BIAS_ADJ[3] 
    ANTENNAPARTIALMETALAREA 0.019 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0836 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.178 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M3 ;
  END BIAS_ADJ[3]
  PIN BIAS_ADJ[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.344 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6016 LAYER M2 ;
  END BIAS_ADJ[2]
  PIN BIAS_ADJ[1] 
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.282 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M4 ;
  END BIAS_ADJ[1]
  PIN BIAS_ADJ[0] 
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.278 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M4 ;
  END BIAS_ADJ[0]
  PIN BIAS_DBP[13] 
    ANTENNAPARTIALMETALAREA 0.031 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1364 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.446 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.718 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2032 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.426 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3184 LAYER M6 ;
  END BIAS_DBP[13]
  PIN BIAS_DBP[12] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.7985 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.4014 LAYER M2 ;
  END BIAS_DBP[12]
  PIN BIAS_DBP[11] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3 ;
  END BIAS_DBP[11]
  PIN BIAS_DBP[10] 
    ANTENNAPARTIALMETALAREA 0.1185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5654 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3888 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.642 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2688 LAYER M4 ;
  END BIAS_DBP[10]
  PIN BIAS_DBP[9] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.278 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.6672 LAYER M4 ;
  END BIAS_DBP[9]
  PIN BIAS_DBP[8] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8288 LAYER M3 ;
  END BIAS_DBP[8]
  PIN BIAS_DBP[7] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
  END BIAS_DBP[7]
  PIN BIAS_DBP[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0675 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.341 LAYER M2 ;
  END BIAS_DBP[6]
  PIN BIAS_DBP[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.064 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3256 LAYER M2 ;
  END BIAS_DBP[5]
  PIN BIAS_DBP[4] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.4255 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9162 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.178 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0544 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.158 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 18.3392 LAYER M6 ;
  END BIAS_DBP[4]
  PIN BIAS_DBP[3] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4352 LAYER M3 ;
  END BIAS_DBP[3]
  PIN BIAS_DBP[2] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.122 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9808 LAYER M4 ;
  END BIAS_DBP[2]
  PIN BIAS_DBP[1] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.782 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M4 ;
  END BIAS_DBP[1]
  PIN BIAS_DBP[0] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.566 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.098 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2752 LAYER M4 ;
  END BIAS_DBP[0]
  PIN BIAS_DBN[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.613 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7412 LAYER M2 ;
  END BIAS_DBN[13]
  PIN BIAS_DBN[12] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.626 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1984 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.258 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.7792 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.918 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.2832 LAYER M6 ;
  END BIAS_DBN[12]
  PIN BIAS_DBN[11] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_DBN[11]
  PIN BIAS_DBN[10] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.3935 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7754 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.998 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 26.4352 LAYER M4 ;
  END BIAS_DBN[10]
  PIN BIAS_DBN[9] 
    ANTENNAPARTIALMETALAREA 0.05 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.422 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.186 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.4624 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.978 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 39.5472 LAYER M6 ;
  END BIAS_DBN[9]
  PIN BIAS_DBN[8] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.702 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1328 LAYER M3 ;
  END BIAS_DBN[8]
  PIN BIAS_DBN[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.236 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M2 ;
  END BIAS_DBN[7]
  PIN BIAS_DBN[6] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.658 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.5392 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 6.302 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.7728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.098 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 13.6752 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 162.882 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 719.276 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA6 ;
  END BIAS_DBN[6]
  PIN BIAS_DBN[5] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.458 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0512 LAYER M4 ;
  END BIAS_DBN[5]
  PIN BIAS_DBN[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.964 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.3296 LAYER M2 ;
  END BIAS_DBN[4]
  PIN BIAS_DBN[3] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.158 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1392 LAYER M4 ;
  END BIAS_DBN[3]
  PIN BIAS_DBN[2] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.6275 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.249 LAYER M3 ;
  END BIAS_DBN[2]
  PIN BIAS_DBN[1] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.418 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 37.0832 LAYER M4 ;
  END BIAS_DBN[1]
  PIN BIAS_DBN[0] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.978 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3472 LAYER M4 ;
  END BIAS_DBN[0]
  PIN BIAS_DBPC[13] 
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.858 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8192 LAYER M3 ;
  END BIAS_DBPC[13]
  PIN BIAS_DBPC[12] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.243 LAYER M2 ;
  END BIAS_DBPC[12]
  PIN BIAS_DBPC[11] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.018 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.1232 LAYER M4 ;
  END BIAS_DBPC[11]
  PIN BIAS_DBPC[10] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.476 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.3824 LAYER M2 ;
  END BIAS_DBPC[10]
  PIN BIAS_DBPC[9] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
  END BIAS_DBPC[9]
  PIN BIAS_DBPC[8] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_DBPC[8]
  PIN BIAS_DBPC[7] 
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.008 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5232 LAYER M3 ;
  END BIAS_DBPC[7]
  PIN BIAS_DBPC[6] 
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.338 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.898 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1952 LAYER M4 ;
  END BIAS_DBPC[6]
  PIN BIAS_DBPC[5] 
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7728 LAYER M3 ;
  END BIAS_DBPC[5]
  PIN BIAS_DBPC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.7105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.4142 LAYER M2 ;
  END BIAS_DBPC[4]
  PIN BIAS_DBPC[3] 
    ANTENNAPARTIALMETALAREA 0.019 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0836 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
  END BIAS_DBPC[3]
  PIN BIAS_DBPC[2] 
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6528 LAYER M3 ;
  END BIAS_DBPC[2]
  PIN BIAS_DBPC[1] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.422 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7008 LAYER M4 ;
  END BIAS_DBPC[1]
  PIN BIAS_DBPC[0] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.278 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6672 LAYER M4 ;
  END BIAS_DBPC[0]
  PIN BIAS_DBNC[13] 
    ANTENNAPARTIALMETALAREA 0.173 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8052 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8368 LAYER M3 ;
  END BIAS_DBNC[13]
  PIN BIAS_DBNC[12] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.426 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3184 LAYER M3 ;
  END BIAS_DBNC[12]
  PIN BIAS_DBNC[11] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.706 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5504 LAYER M3 ;
  END BIAS_DBNC[11]
  PIN BIAS_DBNC[10] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.744 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7616 LAYER M3 ;
  END BIAS_DBNC[10]
  PIN BIAS_DBNC[9] 
    ANTENNAPARTIALMETALAREA 0.019 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0836 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.878 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.3072 LAYER M3 ;
  END BIAS_DBNC[9]
  PIN BIAS_DBNC[8] 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.618 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7632 LAYER M3 ;
  END BIAS_DBNC[8]
  PIN BIAS_DBNC[7] 
    ANTENNAPARTIALMETALAREA 0.03 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.132 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3 ;
  END BIAS_DBNC[7]
  PIN BIAS_DBNC[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0615 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3146 LAYER M2 ;
  END BIAS_DBNC[6]
  PIN BIAS_DBNC[5] 
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.038 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6112 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.226 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4384 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.418 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 32.6832 LAYER M6 ;
  END BIAS_DBNC[5]
  PIN BIAS_DBNC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_DBNC[4]
  PIN BIAS_DBNC[3] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6528 LAYER M3 ;
  END BIAS_DBNC[3]
  PIN BIAS_DBNC[2] 
    ANTENNAPARTIALMETALAREA 0.1105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5302 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.918 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0832 LAYER M3 ;
  END BIAS_DBNC[2]
  PIN BIAS_DBNC[1] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.104 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9456 LAYER M3 ;
  END BIAS_DBNC[1]
  PIN BIAS_DBNC[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0245 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1518 LAYER M2 ;
  END BIAS_DBNC[0]
  PIN BIAS_TC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.5305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3782 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2 ; 
    ANTENNAMAXAREACAR 8.27742 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 36.8629 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.0379 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 45.2439 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.922 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1008 LAYER M4 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 23.3424 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 104.418 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA4 ;
  END BIAS_TC_POT[5]
  PIN BIAS_TC_POT[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.442 LAYER M2 ;
  END BIAS_TC_POT[4]
  PIN BIAS_TC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.2135 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9394 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.586 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6224 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.618 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7632 LAYER M4 ;
  END BIAS_TC_POT[3]
  PIN BIAS_TC_POT[2] 
    ANTENNAPARTIALMETALAREA 0.302 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3288 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.498 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2352 LAYER M3 ;
  END BIAS_TC_POT[2]
  PIN BIAS_TC_POT[1] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.2665 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2166 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.062 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.1168 LAYER M4 ;
  END BIAS_TC_POT[1]
  PIN BIAS_TC_POT[0] 
    ANTENNAPARTIALMETALAREA 0.207 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9108 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M5 ;
  END BIAS_TC_POT[0]
  PIN BIAS_LC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.1325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.583 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.69 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.7482 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 126.309 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_LC_POT[5]
  PIN BIAS_LC_POT[4] 
    ANTENNAPARTIALMETALAREA 0.091 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.139 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6556 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.32 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.296 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ; 
    ANTENNAMAXAREACAR 85.1298 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 376.552 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.63934 LAYER VIA4 ;
  END BIAS_LC_POT[4]
  PIN BIAS_LC_POT[3] 
    ANTENNAPARTIALMETALAREA 1.11 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.928 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.7583 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 108.713 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_LC_POT[3]
  PIN BIAS_LC_POT[2] 
    ANTENNAPARTIALMETALAREA 0.767 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3748 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M2 ; 
    ANTENNAMAXAREACAR 18.357 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 78.2922 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.823045 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.858 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8192 LAYER M3 ;
    ANTENNAGATEAREA 0.0486 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.0113 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 156.877 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.823045 LAYER VIA3 ;
  END BIAS_LC_POT[2]
  PIN BIAS_LC_POT[1] 
    ANTENNAPARTIALMETALAREA 0.6805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9942 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.318 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4432 LAYER M3 ;
  END BIAS_LC_POT[1]
  PIN BIAS_LC_POT[0] 
    ANTENNAPARTIALMETALAREA 0.386 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6984 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3 ;
  END BIAS_LC_POT[0]
  PIN BIAS_TIA_G_POT[16] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3112 LAYER M2 ;
  END BIAS_TIA_G_POT[16]
  PIN BIAS_TIA_G_POT[15] 
    ANTENNAPARTIALMETALAREA 0.9965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3846 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.886 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.7424 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 6.678 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 29.4272 LAYER M5 ;
  END BIAS_TIA_G_POT[15]
  PIN BIAS_TIA_G_POT[14] 
    ANTENNAPARTIALMETALAREA 0.087 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3828 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.726 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2384 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.562 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5168 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.946 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.4064 LAYER M5 ;
  END BIAS_TIA_G_POT[14]
  PIN BIAS_TIA_G_POT[13] 
    ANTENNAPARTIALMETALAREA 0.2455 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0802 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.802 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.878 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1072 LAYER M5 ;
  END BIAS_TIA_G_POT[13]
  PIN BIAS_TIA_G_POT[12] 
    ANTENNAPARTIALMETALAREA 1.214 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3416 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.8288 LAYER M3 ;
  END BIAS_TIA_G_POT[12]
  PIN BIAS_TIA_G_POT[11] 
    ANTENNAPARTIALMETALAREA 0.171 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7524 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.418 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8832 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.062 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.9168 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.402 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M6 ;
  END BIAS_TIA_G_POT[11]
  PIN BIAS_TIA_G_POT[10] 
    ANTENNAPARTIALMETALAREA 1.109 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8796 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.678 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.4272 LAYER M3 ;
  END BIAS_TIA_G_POT[10]
  PIN BIAS_TIA_G_POT[9] 
    ANTENNAPARTIALMETALAREA 0.3475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.529 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.782 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M3 ;
  END BIAS_TIA_G_POT[9]
  PIN BIAS_TIA_G_POT[8] 
    ANTENNAPARTIALMETALAREA 0.301 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.1328 LAYER M3 ;
  END BIAS_TIA_G_POT[8]
  PIN BIAS_TIA_G_POT[7] 
    ANTENNAPARTIALMETALAREA 0.0695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3058 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.566 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.838 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7312 LAYER M4 ;
  END BIAS_TIA_G_POT[7]
  PIN BIAS_TIA_G_POT[6] 
    ANTENNAPARTIALMETALAREA 0.347 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5268 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.466 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0944 LAYER M3 ;
  END BIAS_TIA_G_POT[6]
  PIN BIAS_TIA_G_POT[5] 
    ANTENNAPARTIALMETALAREA 0.1585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6974 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.446 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0064 LAYER M3 ;
  END BIAS_TIA_G_POT[5]
  PIN BIAS_TIA_G_POT[4] 
    ANTENNAPARTIALMETALAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1132 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.526 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M3 ;
  END BIAS_TIA_G_POT[4]
  PIN BIAS_TIA_G_POT[3] 
    ANTENNAPARTIALMETALAREA 0.087 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3828 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.766 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4144 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 17.7363 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 79.7518 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA4 ;
  END BIAS_TIA_G_POT[3]
  PIN BIAS_TIA_G_POT[2] 
    ANTENNAPARTIALMETALAREA 0.615 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.75 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.49675 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 42.228 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.2886 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.2471 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 46.1645 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.742 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3088 LAYER M4 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 20.9542 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 93.9105 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA4 ;
  END BIAS_TIA_G_POT[2]
  PIN BIAS_TIA_G_POT[1] 
    ANTENNAPARTIALMETALAREA 0.0765 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3366 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.146 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.318 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.2432 LAYER M4 ;
  END BIAS_TIA_G_POT[1]
  PIN BIAS_TIA_G_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.278 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7112 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2 ; 
    ANTENNAMAXAREACAR 19.0639 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 84.9582 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.1443 LAYER VIA2 ;
  END BIAS_TIA_G_POT[0]
  PIN BIAS_REV_POT[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.318 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.6432 LAYER M2 ;
  END BIAS_REV_POT[13]
  PIN BIAS_REV_POT[12] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.868 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9072 LAYER M3 ;
  END BIAS_REV_POT[12]
  PIN BIAS_REV_POT[11] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.818 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6432 LAYER M4 ;
  END BIAS_REV_POT[11]
  PIN BIAS_REV_POT[10] 
    ANTENNAPARTIALMETALAREA 0.7465 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2846 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.606 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7104 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.938 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5712 LAYER M4 ;
  END BIAS_REV_POT[10]
  PIN BIAS_REV_POT[9] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.398 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.4392 LAYER M2 ;
  END BIAS_REV_POT[9]
  PIN BIAS_REV_POT[8] 
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0512 LAYER M4 ;
  END BIAS_REV_POT[8]
  PIN BIAS_REV_POT[7] 
    ANTENNAPARTIALMETALAREA 0.11 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.484 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.722 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2208 LAYER M3 ;
  END BIAS_REV_POT[7]
  PIN BIAS_REV_POT[6] 
    ANTENNAPARTIALMETALAREA 0.0215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0946 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.678 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0272 LAYER M3 ;
  END BIAS_REV_POT[6]
  PIN BIAS_REV_POT[5] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.141 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6644 LAYER M2 ;
  END BIAS_REV_POT[5]
  PIN BIAS_REV_POT[4] 
    ANTENNAPARTIALMETALAREA 0.0705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3102 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9568 LAYER M3 ;
  END BIAS_REV_POT[4]
  PIN BIAS_REV_POT[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.528 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3672 LAYER M2 ;
  END BIAS_REV_POT[3]
  PIN BIAS_REV_POT[2] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0245 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1518 LAYER M2 ;
  END BIAS_REV_POT[2]
  PIN BIAS_REV_POT[1] 
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.718 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2032 LAYER M3 ;
  END BIAS_REV_POT[1]
  PIN BIAS_REV_POT[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4158 LAYER M2 ;
  END BIAS_REV_POT[0]
  PIN BIAS_TC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.4585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0174 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.738 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2912 LAYER M3 ;
  END BIAS_TC_DSADC[5]
  PIN BIAS_TC_DSADC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.65 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.904 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.478 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.45 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.297 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.333333 LAYER VIA3 ;
  END BIAS_TC_DSADC[4]
  PIN BIAS_TC_DSADC[3] 
    ANTENNAPARTIALMETALAREA 1.0735 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7234 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.838 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1312 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.539 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 147.388 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_TC_DSADC[3]
  PIN BIAS_TC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.671 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9524 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.715 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 108.257 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_TC_DSADC[2]
  PIN BIAS_TC_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.6105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6862 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7904 LAYER M3 ;
  END BIAS_TC_DSADC[1]
  PIN BIAS_TC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 1.045 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.642 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2448 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.8737 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.221 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_TC_DSADC[0]
  PIN BIAS_LC_DSADC[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.1165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0006 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.616 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.0332 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 264.524 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA3 ;
  END BIAS_LC_DSADC[5]
  PIN BIAS_LC_DSADC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.029 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.0596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 55.6448 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 241.042 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA3 ;
  END BIAS_LC_DSADC[4]
  PIN BIAS_LC_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.0215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5386 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.822 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0608 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 68.5121 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 300.175 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA3 ;
  END BIAS_LC_DSADC[3]
  PIN BIAS_LC_DSADC[2] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.49 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER M2 ;
  END BIAS_LC_DSADC[2]
  PIN BIAS_LC_DSADC[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.1155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9522 LAYER M2 ;
  END BIAS_LC_DSADC[1]
  PIN BIAS_LC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 1.132 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9808 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.566 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.9488 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 134.231 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_LC_DSADC[0]
  PIN BIAS_RIN_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.1855 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8162 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.542 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4288 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.618 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1632 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M5 ; 
    ANTENNAMAXAREACAR 102.165 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 453.592 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.26537 LAYER VIA5 ;
  END BIAS_RIN_DSADC[5]
  PIN BIAS_RIN_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.775 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.41 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 54.4628 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 240.854 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3 ;
  END BIAS_RIN_DSADC[4]
  PIN BIAS_RIN_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.402 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M2 ; 
    ANTENNAMAXAREACAR 48.3463 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 213.942 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.323625 LAYER VIA2 ;
  END BIAS_RIN_DSADC[3]
  PIN BIAS_RIN_DSADC[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.118 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9632 LAYER M2 ;
  END BIAS_RIN_DSADC[2]
  PIN BIAS_RIN_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.8305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6542 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.684 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 63.4595 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 281.864 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3 ;
  END BIAS_RIN_DSADC[1]
  PIN BIAS_RIN_DSADC[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.613 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1852 LAYER M2 ;
  END BIAS_RIN_DSADC[0]
  PIN BIAS_RFB_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5346 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.962 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 LAYER M3 ; 
    ANTENNAMAXAREACAR 51.7748 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 227.908 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VIA3 ;
  END BIAS_RFB_DSADC[5]
  PIN BIAS_RFB_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.153 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6732 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.502 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 21.28 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 93.72 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.082 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8048 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 3.588 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8752 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M7 ; 
    ANTENNAMAXAREACAR 288.189 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 1260.12 LAYER M7 ;
    ANTENNAMAXCUTCAR 3.8835 LAYER VIA7 ;
  END BIAS_RFB_DSADC[4]
  PIN BIAS_RFB_DSADC[3] 
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.4415 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9866 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.762 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3968 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 LAYER M4 ; 
    ANTENNAMAXAREACAR 41.6223 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 184.461 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VIA4 ;
  END BIAS_RFB_DSADC[3]
  PIN BIAS_RFB_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.085 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.374 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.958 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.246 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.598 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0752 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M5 ; 
    ANTENNAMAXAREACAR 277.204 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1225.4 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.589 LAYER VIA5 ;
  END BIAS_RFB_DSADC[2]
  PIN BIAS_RFB_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.3755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6522 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.802 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5728 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 103.852 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 457.327 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA4 ;
  END BIAS_RFB_DSADC[1]
  PIN BIAS_RFB_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.137 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6028 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.766 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4144 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.898 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9952 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.226 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 441.294 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1949.05 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.23625 LAYER VIA6 ;
  END BIAS_RFB_DSADC[0]
  PIN BIAS_DSADC_VCM[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.19 LAYER M2 ;
  END BIAS_DSADC_VCM[13]
  PIN BIAS_DSADC_VCM[12] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.942 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1888 LAYER M4 ;
  END BIAS_DSADC_VCM[12]
  PIN BIAS_DSADC_VCM[11] 
    ANTENNAPARTIALMETALAREA 2.529 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.1276 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.426 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9184 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.778 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.8672 LAYER M4 ;
  END BIAS_DSADC_VCM[11]
  PIN BIAS_DSADC_VCM[10] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
  END BIAS_DSADC_VCM[10]
  PIN BIAS_DSADC_VCM[9] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.411 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.4964 LAYER M2 ;
  END BIAS_DSADC_VCM[9]
  PIN BIAS_DSADC_VCM[8] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.158 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1392 LAYER M4 ;
  END BIAS_DSADC_VCM[8]
  PIN BIAS_DSADC_VCM[7] 
    ANTENNAPARTIALMETALAREA 0.158 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7392 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9568 LAYER M3 ;
  END BIAS_DSADC_VCM[7]
  PIN BIAS_DSADC_VCM[6] 
    ANTENNAPARTIALMETALAREA 0.0625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
  END BIAS_DSADC_VCM[6]
  PIN BIAS_DSADC_VCM[5] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.758 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3792 LAYER M3 ;
  END BIAS_DSADC_VCM[5]
  PIN BIAS_DSADC_VCM[4] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
  END BIAS_DSADC_VCM[4]
  PIN BIAS_DSADC_VCM[3] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.008 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 6.802 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 29.9728 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 102.543 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 452.277 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA5 ;
  END BIAS_DSADC_VCM[3]
  PIN BIAS_DSADC_VCM[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0655 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3322 LAYER M2 ;
  END BIAS_DSADC_VCM[2]
  PIN BIAS_DSADC_VCM[1] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3 ;
  END BIAS_DSADC_VCM[1]
  PIN BIAS_DSADC_VCM[0] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.546 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4464 LAYER M3 ;
  END BIAS_DSADC_VCM[0]
  PIN dsadc_conv_done 
    ANTENNAPARTIALMETALAREA 0.042 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1848 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.278 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.402 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2128 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 12.446 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 54.8944 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0381 LAYER M5 ; 
    ANTENNAMAXAREACAR 384.411 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1684.27 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.09974 LAYER VIA5 ;
  END dsadc_conv_done
  PIN dsadc_en 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.288 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3112 LAYER M2 ;
  END dsadc_en
  PIN dsadc_clk 
    ANTENNAPARTIALMETALAREA 0.196 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2156 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 61.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.4982 LAYER M3 ;
  END dsadc_clk
  PIN dsadc_switch[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1858 LAYER M2 ;
  END dsadc_switch[2]
  PIN dsadc_switch[1] 
    ANTENNAPARTIALMETALAREA 0.244 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0736 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.938 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5712 LAYER M3 ;
  END dsadc_switch[1]
  PIN dsadc_switch[0] 
    ANTENNAPARTIALMETALAREA 0.6225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.739 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8368 LAYER M3 ;
  END dsadc_switch[0]
  PIN dac_en_pot 
    ANTENNAPARTIALMETALAREA 0.8065 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.026 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.5584 LAYER M3 ;
  END dac_en_pot
  PIN adc_ext_in 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.342 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M2 ;
  END adc_ext_in
  PIN atp_en 
    ANTENNAPARTIALMETALAREA 0.4445 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9558 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.002 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.8528 LAYER M3 ;
  END atp_en
  PIN atp_sel 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.738 LAYER M2 ;
  END atp_sel
  PIN adc_sel 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8546 LAYER M2 ;
  END adc_sel
  PIN saradc_clk 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.8042 LAYER M3 ;
  END saradc_clk
  PIN saradc_rdy 
    ANTENNAPARTIALMETALAREA 0.131 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5764 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.484 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.618 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7632 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M5 ; 
    ANTENNAMAXAREACAR 278.703 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1227.84 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.30548 LAYER VIA5 ;
  END saradc_rdy
  PIN saradc_rst 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2682 LAYER M2 ;
  END saradc_rst
  PIN saradc_data[9] 
    ANTENNAPARTIALMETALAREA 0.087 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3828 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.8215 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6586 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.404 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2656 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.778 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.0672 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.606 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7104 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6 ; 
    ANTENNAMAXAREACAR 195.333 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 865.486 LAYER M6 ;
    ANTENNAMAXCUTCAR 4.08163 LAYER VIA6 ;
  END saradc_data[9]
  PIN saradc_data[8] 
    ANTENNAPARTIALMETALAREA 0.1515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 6.844 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.2016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 6.678 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 29.4272 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 0.946 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2064 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M7 ; 
    ANTENNAMAXAREACAR 174.435 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 759.135 LAYER M7 ;
    ANTENNAMAXCUTCAR 4.89796 LAYER VIA7 ;
  END saradc_data[8]
  PIN saradc_data[7] 
    ANTENNAPARTIALMETALAREA 0.3515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5466 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.642 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8688 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.946 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2064 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 16.424 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 72.3536 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 723.796 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 3192.06 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.85714 LAYER VIA5 ;
  END saradc_data[7]
  PIN saradc_data[6] 
    ANTENNAPARTIALMETALAREA 0.1915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8426 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.782 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 15.778 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 69.4672 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 1.418 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2832 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6 ; 
    ANTENNAMAXAREACAR 78.0265 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 349.306 LAYER M6 ;
    ANTENNAMAXCUTCAR 4.08163 LAYER VIA6 ;
  END saradc_data[6]
  PIN saradc_data[5] 
    ANTENNAPARTIALMETALAREA 0.2315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0186 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.026 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.9584 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.222 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.6208 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M5 ; 
    ANTENNAMAXAREACAR 140.579 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 617.929 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.01511 LAYER VIA5 ;
  END saradc_data[5]
  PIN saradc_data[4] 
    ANTENNAPARTIALMETALAREA 0.7425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.267 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.978 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3472 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 12.378 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 54.5072 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 683.186 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2995.25 LAYER M5 ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5 ;
  END saradc_data[4]
  PIN saradc_data[3] 
    ANTENNAPARTIALMETALAREA 0.5845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6158 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.558 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6992 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.146 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 9.196 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 40.5504 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 399.659 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1761.26 LAYER M5 ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5 ;
  END saradc_data[3]
  PIN saradc_data[2] 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.62972 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 43.6625 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.251889 LAYER VIA2 ;
  END saradc_data[2]
  PIN saradc_data[1] 
    ANTENNAPARTIALMETALAREA 0.9025 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.971 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 5.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.3968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 7.818 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 34.4432 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.622 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7808 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6 ; 
    ANTENNAMAXAREACAR 206.859 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 901.796 LAYER M6 ;
    ANTENNAMAXCUTCAR 4.08163 LAYER VIA6 ;
  END saradc_data[1]
  PIN saradc_data[0] 
    ANTENNAPARTIALMETALAREA 0.3595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5818 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.9088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 266.826 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1167.91 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END saradc_data[0]
END MCU

END LIBRARY
