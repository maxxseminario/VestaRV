

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO MCU 
  PIN resetn_in 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3408 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 25.822 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 113.661 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6 ; 
    ANTENNAMAXAREACAR 974.972 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4296.54 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.32103 LAYER VIA6 ;
  END resetn_in
  PIN resetn_out 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.474 LAYER M2 ;
  END resetn_out
  PIN resetn_dir 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6365 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8446 LAYER M2 ;
  END resetn_dir
  PIN resetn_ren 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5895 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6378 LAYER M2 ;
  END resetn_ren
  PIN prt1_in[7] 
    ANTENNAPARTIALMETALAREA 3.9755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.4922 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 25.778 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 113.467 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 771.741 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3377.47 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt1_in[7]
  PIN prt1_in[6] 
    ANTENNAPARTIALMETALAREA 20.6525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 90.871 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 5.918 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.0832 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0269 LAYER M3 ; 
    ANTENNAMAXAREACAR 313.729 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1381.81 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.48699 LAYER VIA3 ;
  END prt1_in[6]
  PIN prt1_in[5] 
    ANTENNAPARTIALMETALAREA 3.6505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.1062 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 24.162 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 106.357 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0381 LAYER M3 ; 
    ANTENNAMAXAREACAR 649.03 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2856.09 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.04987 LAYER VIA3 ;
  END prt1_in[5]
  PIN prt1_in[4] 
    ANTENNAPARTIALMETALAREA 0.2725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.882 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.5248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 8.578 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 37.7872 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0893 LAYER M5 ; 
    ANTENNAMAXAREACAR 102.572 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 451.807 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.895857 LAYER VIA5 ;
  END prt1_in[4]
  PIN prt1_in[3] 
    ANTENNAPARTIALMETALAREA 0.176 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1936 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6182 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.344 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3816 LAYER M4 ; 
    ANTENNAMAXAREACAR 18.8268 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 24.2175 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.366876 LAYER VIA4 ;
  END prt1_in[3]
  PIN prt1_in[2] 
    ANTENNAPARTIALMETALAREA 4.3395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.0938 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.642 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.8688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 LAYER M3 ; 
    ANTENNAMAXAREACAR 157.444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 688.959 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.542005 LAYER VIA3 ;
  END prt1_in[2]
  PIN prt1_in[1] 
    ANTENNAPARTIALMETALAREA 1.2935 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.982 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.7648 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 350.151 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1541.07 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END prt1_in[1]
  PIN prt1_in[0] 
    ANTENNAPARTIALMETALAREA 10.9995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 48.3978 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.9056 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0893 LAYER M3 ; 
    ANTENNAMAXAREACAR 52.8511 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 233.2 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.335946 LAYER VIA3 ;
  END prt1_in[0]
  PIN prt1_out[7] 
    ANTENNAPARTIALMETALAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5584 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.532 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8288 LAYER M3 ;
  END prt1_out[7]
  PIN prt1_out[6] 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.426 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7184 LAYER M3 ;
  END prt1_out[6]
  PIN prt1_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.376 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M2 ;
  END prt1_out[5]
  PIN prt1_out[4] 
    ANTENNAPARTIALMETALAREA 0.176 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.186 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M3 ;
  END prt1_out[4]
  PIN prt1_out[3] 
    ANTENNAPARTIALMETALAREA 0.956 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2064 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.526 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7584 LAYER M3 ;
  END prt1_out[3]
  PIN prt1_out[2] 
    ANTENNAPARTIALMETALAREA 1.712 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5328 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3 ;
  END prt1_out[2]
  PIN prt1_out[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2 ;
  END prt1_out[1]
  PIN prt1_out[0] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2 ;
  END prt1_out[0]
  PIN prt1_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.8395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1818 LAYER M2 ;
  END prt1_dir[7]
  PIN prt1_dir[6] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.426 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7184 LAYER M3 ;
  END prt1_dir[6]
  PIN prt1_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5126 LAYER M2 ;
  END prt1_dir[5]
  PIN prt1_dir[4] 
    ANTENNAPARTIALMETALAREA 0.0965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4246 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.626 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.3984 LAYER M3 ;
  END prt1_dir[4]
  PIN prt1_dir[3] 
    ANTENNAPARTIALMETALAREA 0.2365 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0406 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.706 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.7504 LAYER M3 ;
  END prt1_dir[3]
  PIN prt1_dir[2] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1946 LAYER M2 ;
  END prt1_dir[2]
  PIN prt1_dir[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2 ;
  END prt1_dir[1]
  PIN prt1_dir[0] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2 ;
  END prt1_dir[0]
  PIN prt1_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M2 ;
  END prt1_ren[7]
  PIN prt1_ren[6] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.266 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2144 LAYER M3 ;
  END prt1_ren[6]
  PIN prt1_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5302 LAYER M2 ;
  END prt1_ren[5]
  PIN prt1_ren[4] 
    ANTENNAPARTIALMETALAREA 0.5205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.406 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8304 LAYER M3 ;
  END prt1_ren[4]
  PIN prt1_ren[3] 
    ANTENNAPARTIALMETALAREA 0.9005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9622 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.606 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.7104 LAYER M3 ;
  END prt1_ren[3]
  PIN prt1_ren[2] 
    ANTENNAPARTIALMETALAREA 4.4675 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.657 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8368 LAYER M3 ;
  END prt1_ren[2]
  PIN prt1_ren[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.1495 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.7018 LAYER M2 ;
  END prt1_ren[1]
  PIN prt1_ren[0] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
  END prt1_ren[0]
  PIN prt2_in[7] 
    ANTENNAPARTIALMETALAREA 0.5505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4662 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2 ; 
    ANTENNAMAXAREACAR 7.12421 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 30.0865 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA2 ;
  END prt2_in[7]
  PIN prt2_in[6] 
    ANTENNAPARTIALMETALAREA 0.7555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4122 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2 ; 
    ANTENNAMAXAREACAR 24.683 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 109.072 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2 ;
  END prt2_in[6]
  PIN prt2_in[5] 
    ANTENNAPARTIALMETALAREA 0.7325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.223 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 LAYER M2 ; 
    ANTENNAMAXAREACAR 7.31574 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 31.5093 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VIA2 ;
  END prt2_in[5]
  PIN prt2_in[4] 
    ANTENNAPARTIALMETALAREA 0.331 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 5.702 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.1328 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 180.086 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 789.527 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt2_in[4]
  PIN prt2_in[3] 
    ANTENNAPARTIALMETALAREA 1.328 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.28166 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 5.07296 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0419287 LAYER VIA2 ;
  END prt2_in[3]
  PIN prt2_in[2] 
    ANTENNAPARTIALMETALAREA 0.2995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3178 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.03459 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 8.46331 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.104822 LAYER VIA2 ;
  END prt2_in[2]
  PIN prt2_in[1] 
    ANTENNAPARTIALMETALAREA 0.4785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1054 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M2 ; 
    ANTENNAMAXAREACAR 4.13417 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 17.2138 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.104822 LAYER VIA2 ;
  END prt2_in[1]
  PIN prt2_in[0] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 23.782 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 104.685 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1476 LAYER M3 ; 
    ANTENNAMAXAREACAR 176.163 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 770.575 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.271003 LAYER VIA3 ;
  END prt2_in[0]
  PIN prt2_out[7] 
    ANTENNAPARTIALMETALAREA 0.711 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1284 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.0928 LAYER M3 ;
  END prt2_out[7]
  PIN prt2_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.681 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2 ;
  END prt2_out[6]
  PIN prt2_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.234 LAYER M2 ;
  END prt2_out[5]
  PIN prt2_out[4] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2 ;
  END prt2_out[4]
  PIN prt2_out[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.317 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4388 LAYER M2 ;
  END prt2_out[3]
  PIN prt2_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.579 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6356 LAYER M2 ;
  END prt2_out[2]
  PIN prt2_out[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.279 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2276 LAYER M2 ;
  END prt2_out[1]
  PIN prt2_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.292 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M2 ;
  END prt2_out[0]
  PIN prt2_dir[7] 
    ANTENNAPARTIALMETALAREA 0.6565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8886 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.106 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.9104 LAYER M3 ;
  END prt2_dir[7]
  PIN prt2_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2186 LAYER M2 ;
  END prt2_dir[6]
  PIN prt2_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2186 LAYER M2 ;
  END prt2_dir[5]
  PIN prt2_dir[4] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.4448 LAYER M3 ;
  END prt2_dir[4]
  PIN prt2_dir[3] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M2 ;
  END prt2_dir[3]
  PIN prt2_dir[2] 
    ANTENNAPARTIALMETALAREA 0.431 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8964 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 59.8928 LAYER M3 ;
  END prt2_dir[2]
  PIN prt2_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9018 LAYER M2 ;
  END prt2_dir[1]
  PIN prt2_dir[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3046 LAYER M2 ;
  END prt2_dir[0]
  PIN prt2_ren[7] 
    ANTENNAPARTIALMETALAREA 0.4835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1274 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.7248 LAYER M3 ;
  END prt2_ren[7]
  PIN prt2_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3562 LAYER M2 ;
  END prt2_ren[6]
  PIN prt2_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2362 LAYER M2 ;
  END prt2_ren[5]
  PIN prt2_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.519 LAYER M2 ;
  END prt2_ren[4]
  PIN prt2_ren[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2154 LAYER M2 ;
  END prt2_ren[3]
  PIN prt2_ren[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8622 LAYER M2 ;
  END prt2_ren[2]
  PIN prt2_ren[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3222 LAYER M2 ;
  END prt2_ren[1]
  PIN prt2_ren[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4895 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1978 LAYER M2 ;
  END prt2_ren[0]
  PIN prt3_in[7] 
    ANTENNAPARTIALMETALAREA 18.7995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 82.8058 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2 ; 
    ANTENNAMAXAREACAR 545.72 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2401.22 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2 ;
  END prt3_in[7]
  PIN prt3_in[6] 
    ANTENNAPARTIALMETALAREA 16.1105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 70.9302 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 14.798 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.1552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 562.952 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2474.57 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[6]
  PIN prt3_in[5] 
    ANTENNAPARTIALMETALAREA 6.6925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.447 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 15.026 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.1584 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.62 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.616 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 53.3072 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 237.512 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.71003 LAYER VIA4 ;
  END prt3_in[5]
  PIN prt3_in[4] 
    ANTENNAPARTIALMETALAREA 0.6925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.047 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 14.586 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.2224 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.526 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M5 ; 
    ANTENNAMAXAREACAR 17.5911 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 77.4752 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.927362 LAYER VIA5 ;
  END prt3_in[4]
  PIN prt3_in[3] 
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 22.168 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 97.6272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1707 LAYER M3 ; 
    ANTENNAMAXAREACAR 166.842 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 733.458 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.734684 LAYER VIA3 ;
  END prt3_in[3]
  PIN prt3_in[2] 
    ANTENNAPARTIALMETALAREA 12.2535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 53.9594 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 14.638 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.4512 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 563.852 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2462.88 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[2]
  PIN prt3_in[1] 
    ANTENNAPARTIALMETALAREA 19.1205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 84.1742 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2 ; 
    ANTENNAMAXAREACAR 710.646 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3125.19 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.738007 LAYER VIA2 ;
  END prt3_in[1]
  PIN prt3_in[0] 
    ANTENNAPARTIALMETALAREA 1.8725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.239 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.518 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.9232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 294.334 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1280.41 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt3_in[0]
  PIN prt3_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 15.203 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 66.9812 LAYER M2 ;
  END prt3_out[7]
  PIN prt3_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 6.001 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.5364 LAYER M2 ;
  END prt3_out[6]
  PIN prt3_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.241 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1044 LAYER M2 ;
  END prt3_out[5]
  PIN prt3_out[4] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.157 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7348 LAYER M2 ;
  END prt3_out[4]
  PIN prt3_out[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.157 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7348 LAYER M2 ;
  END prt3_out[3]
  PIN prt3_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.257 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.5748 LAYER M2 ;
  END prt3_out[2]
  PIN prt3_out[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.683 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 60.2932 LAYER M2 ;
  END prt3_out[1]
  PIN prt3_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.943 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.4372 LAYER M2 ;
  END prt3_out[0]
  PIN prt3_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.9215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.2986 LAYER M2 ;
  END prt3_dir[7]
  PIN prt3_dir[6] 
    ANTENNAPARTIALMETALAREA 5.0785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.586 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6224 LAYER M3 ;
  END prt3_dir[6]
  PIN prt3_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt3_dir[5]
  PIN prt3_dir[4] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2 ;
  END prt3_dir[4]
  PIN prt3_dir[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END prt3_dir[3]
  PIN prt3_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.2725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.331 LAYER M2 ;
  END prt3_dir[2]
  PIN prt3_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.9165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.3646 LAYER M2 ;
  END prt3_dir[1]
  PIN prt3_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.8835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.7754 LAYER M2 ;
  END prt3_dir[0]
  PIN prt3_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.5435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.6794 LAYER M2 ;
  END prt3_ren[7]
  PIN prt3_ren[6] 
    ANTENNAPARTIALMETALAREA 4.7585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.9814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.106 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3104 LAYER M3 ;
  END prt3_ren[6]
  PIN prt3_ren[5] 
    ANTENNAPARTIALMETALAREA 6.5785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.9894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.2448 LAYER M3 ;
  END prt3_ren[5]
  PIN prt3_ren[4] 
    ANTENNAPARTIALMETALAREA 0.2605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1462 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.738 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.0912 LAYER M3 ;
  END prt3_ren[4]
  PIN prt3_ren[3] 
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.162 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M3 ;
  END prt3_ren[3]
  PIN prt3_ren[2] 
    ANTENNAPARTIALMETALAREA 8.8055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 38.7882 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.766 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4144 LAYER M3 ;
  END prt3_ren[2]
  PIN prt3_ren[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.8905 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.6062 LAYER M2 ;
  END prt3_ren[1]
  PIN prt3_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.5255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2442 LAYER M2 ;
  END prt3_ren[0]
  PIN prt4_in[7] 
    ANTENNAPARTIALMETALAREA 1.9555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6042 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 27.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 119.821 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.438 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7712 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1456 LAYER M4 ; 
    ANTENNAMAXAREACAR 73.3885 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 321.007 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.76338 LAYER VIA4 ;
  END prt4_in[7]
  PIN prt4_in[6] 
    ANTENNAPARTIALMETALAREA 2.1155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3082 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 17.864 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 78.6896 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 268.215 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1176.6 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.16802 LAYER VIA3 ;
  END prt4_in[6]
  PIN prt4_in[5] 
    ANTENNAPARTIALMETALAREA 1.3185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8014 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.062 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.3168 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 5.198 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.9152 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1456 LAYER M4 ; 
    ANTENNAMAXAREACAR 52.3306 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 231.477 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA4 ;
  END prt4_in[5]
  PIN prt4_in[4] 
    ANTENNAPARTIALMETALAREA 6.2955 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.7002 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.224 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.8736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.9176 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.877 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA3 ;
  END prt4_in[4]
  PIN prt4_in[3] 
    ANTENNAPARTIALMETALAREA 6.5305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.7782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.766 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4144 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1204 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.725 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 62.6902 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.708118 LAYER VIA3 ;
  END prt4_in[3]
  PIN prt4_in[2] 
    ANTENNAPARTIALMETALAREA 7.5505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.746 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.865 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 64.0081 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.734684 LAYER VIA3 ;
  END prt4_in[2]
  PIN prt4_in[1] 
    ANTENNAPARTIALMETALAREA 0.2725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 19.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.9904 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 761.255 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3332.75 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt4_in[1]
  PIN prt4_in[0] 
    ANTENNAPARTIALMETALAREA 0.491 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1604 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 28.578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 125.787 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 1084.22 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4750.11 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt4_in[0]
  PIN prt4_out[7] 
    ANTENNAPARTIALMETALAREA 5.292 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8806 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 46.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.48 LAYER M3 ;
  END prt4_out[7]
  PIN prt4_out[6] 
    ANTENNAPARTIALMETALAREA 0.172 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 18.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.0662 LAYER M3 ;
  END prt4_out[6]
  PIN prt4_out[5] 
    ANTENNAPARTIALMETALAREA 0.172 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 12.882 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.3462 LAYER M3 ;
  END prt4_out[5]
  PIN prt4_out[4] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.8902 LAYER M3 ;
  END prt4_out[4]
  PIN prt4_out[3] 
    ANTENNAPARTIALMETALAREA 0.939 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1316 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.142 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.0688 LAYER M3 ;
  END prt4_out[3]
  PIN prt4_out[2] 
    ANTENNAPARTIALMETALAREA 0.639 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8116 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.0784 LAYER M3 ;
  END prt4_out[2]
  PIN prt4_out[1] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.946 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 74.6064 LAYER M6 ;
  END prt4_out[1]
  PIN prt4_out[0] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
  END prt4_out[0]
  PIN prt4_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.2965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1486 LAYER M2 ;
  END prt4_dir[7]
  PIN prt4_dir[6] 
    ANTENNAPARTIALMETALAREA 1.231 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4164 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 12.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.8912 LAYER M3 ;
  END prt4_dir[6]
  PIN prt4_dir[5] 
    ANTENNADIFFAREA 1.968 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.7945 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3838 LAYER M2 ;
  END prt4_dir[5]
  PIN prt4_dir[4] 
    ANTENNADIFFAREA 1.968 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.9585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.5054 LAYER M2 ;
  END prt4_dir[4]
  PIN prt4_dir[3] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.5808 LAYER M3 ;
  END prt4_dir[3]
  PIN prt4_dir[2] 
    ANTENNAPARTIALMETALAREA 0.3565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5686 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.106 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.7104 LAYER M3 ;
  END prt4_dir[2]
  PIN prt4_dir[1] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 17.122 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 75.3808 LAYER M6 ;
  END prt4_dir[1]
  PIN prt4_dir[0] 
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.362 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 72.0368 LAYER M6 ;
  END prt4_dir[0]
  PIN prt4_ren[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2286 LAYER M2 ;
  END prt4_ren[7]
  PIN prt4_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.431 LAYER M2 ;
  END prt4_ren[6]
  PIN prt4_ren[5] 
    ANTENNAPARTIALMETALAREA 0.4945 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1758 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.962 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.0768 LAYER M3 ;
  END prt4_ren[5]
  PIN prt4_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.2095 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3658 LAYER M2 ;
  END prt4_ren[4]
  PIN prt4_ren[3] 
    ANTENNAPARTIALMETALAREA 0.9035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9754 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.9408 LAYER M3 ;
  END prt4_ren[3]
  PIN prt4_ren[2] 
    ANTENNAPARTIALMETALAREA 0.7435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2714 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 12.962 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.0768 LAYER M3 ;
  END prt4_ren[2]
  PIN prt4_ren[1] 
    ANTENNAPARTIALMETALAREA 0.8035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.342 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 71.9488 LAYER M6 ;
  END prt4_ren[1]
  PIN prt4_ren[0] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 17.122 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 75.3808 LAYER M6 ;
  END prt4_ren[0]
  PIN use_dac_glb_bias 
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.478 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 41.7472 LAYER M6 ;
  END use_dac_glb_bias
  PIN en_bias_buf 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.979 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.5956 LAYER M2 ;
  END en_bias_buf
  PIN en_bias_gen 
    ANTENNAPARTIALMETALAREA 0.081 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.226 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M3 ;
  END en_bias_gen
  PIN BIAS_ADJ[5] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M3 ;
  END BIAS_ADJ[5]
  PIN BIAS_ADJ[4] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
  END BIAS_ADJ[4]
  PIN BIAS_ADJ[3] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.378 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7072 LAYER M3 ;
  END BIAS_ADJ[3]
  PIN BIAS_ADJ[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2665 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2606 LAYER M2 ;
  END BIAS_ADJ[2]
  PIN BIAS_ADJ[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.872 LAYER M2 ;
  END BIAS_ADJ[1]
  PIN BIAS_ADJ[0] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.418 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8832 LAYER M3 ;
  END BIAS_ADJ[0]
  PIN BIAS_DBP[13] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
  END BIAS_DBP[13]
  PIN BIAS_DBP[12] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3088 LAYER M3 ;
  END BIAS_DBP[12]
  PIN BIAS_DBP[11] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.265 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.254 LAYER M2 ;
  END BIAS_DBP[11]
  PIN BIAS_DBP[10] 
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.562 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5168 LAYER M3 ;
  END BIAS_DBP[10]
  PIN BIAS_DBP[9] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.664 LAYER M3 ;
  END BIAS_DBP[9]
  PIN BIAS_DBP[8] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1474 LAYER M2 ;
  END BIAS_DBP[8]
  PIN BIAS_DBP[7] 
    ANTENNAPARTIALMETALAREA 0.024 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1056 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3608 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.366 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M5 ;
  END BIAS_DBP[7]
  PIN BIAS_DBP[6] 
    ANTENNAPARTIALMETALAREA 0.0185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.458 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.178 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 42.7768 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 1.242 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5088 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 221.356 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 972.227 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.77994 LAYER VIA7 ;
  END BIAS_DBP[6]
  PIN BIAS_DBP[5] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.178 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.4272 LAYER M4 ;
  END BIAS_DBP[5]
  PIN BIAS_DBP[4] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.5655 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9322 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.938 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1712 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.482 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5648 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.078 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 44.3872 LAYER M6 ;
  END BIAS_DBP[4]
  PIN BIAS_DBP[3] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6528 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.426 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7184 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.698 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 51.5152 LAYER M6 ;
  END BIAS_DBP[3]
  PIN BIAS_DBP[2] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.878 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9072 LAYER M3 ;
  END BIAS_DBP[2]
  PIN BIAS_DBP[1] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.158 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7392 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.366 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8544 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.338 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 45.5312 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 586.489 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2587.24 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6 ;
  END BIAS_DBP[1]
  PIN BIAS_DBP[0] 
    ANTENNAPARTIALMETALAREA 0.0225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.099 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.002 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6528 LAYER M4 ;
  END BIAS_DBP[0]
  PIN BIAS_DBN[13] 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5648 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.898 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.5952 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.412 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3008 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.662 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9568 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 36.9517 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 164.638 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.2987 LAYER VIA6 ;
  END BIAS_DBN[13]
  PIN BIAS_DBN[12] 
    ANTENNAPARTIALMETALAREA 2.434 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7536 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.078 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.9872 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.938 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7712 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.608 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.9632 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 73.3369 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 324.404 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA5 ;
  END BIAS_DBN[12]
  PIN BIAS_DBN[11] 
    ANTENNAPARTIALMETALAREA 0.157 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7348 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.018 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.7232 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.146 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.478 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 19.7472 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 244.766 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1082.65 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.26537 LAYER VIA6 ;
  END BIAS_DBN[11]
  PIN BIAS_DBN[10] 
    ANTENNAPARTIALMETALAREA 0.0315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1386 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 8.296 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 36.5904 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 0.126 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M7 ; 
    ANTENNAMAXAREACAR 86.9372 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 384.574 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.7316 LAYER VIA7 ;
  END BIAS_DBN[10]
  PIN BIAS_DBN[9] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.748 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.158 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7392 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 8.21 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 36.256 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 133.157 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 588.482 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA5 ;
  END BIAS_DBN[9]
  PIN BIAS_DBN[8] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.558 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.0992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.106 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.078 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.9872 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 297.82 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1317.91 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.23625 LAYER VIA6 ;
  END BIAS_DBN[8]
  PIN BIAS_DBN[7] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.324 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5136 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.358 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.2192 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 167.938 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 740.337 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA4 ;
  END BIAS_DBN[7]
  PIN BIAS_DBN[6] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.384 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M3 ; 
    ANTENNAMAXAREACAR 53.7582 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 230.082 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.823045 LAYER VIA3 ;
  END BIAS_DBN[6]
  PIN BIAS_DBN[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.608 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.7632 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.262 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9968 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.95 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 26.312 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ; 
    ANTENNAMAXAREACAR 201.807 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 896 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.18579 LAYER VIA6 ;
  END BIAS_DBN[5]
  PIN BIAS_DBN[4] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.566 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.242 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 23.1088 LAYER M4 ;
  END BIAS_DBN[4]
  PIN BIAS_DBN[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.932 LAYER M2 ;
  END BIAS_DBN[3]
  PIN BIAS_DBN[2] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.6255 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M3 ; 
    ANTENNAMAXAREACAR 133.04 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 586.021 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.823045 LAYER VIA3 ;
  END BIAS_DBN[2]
  PIN BIAS_DBN[1] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.398 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1952 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.018 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 26.5232 LAYER M4 ;
  END BIAS_DBN[1]
  PIN BIAS_DBN[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.1235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4314 LAYER M2 ;
  END BIAS_DBN[0]
  PIN BIAS_DBPC[13] 
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4912 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.046 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.4464 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 10.18 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 44.88 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 1.326 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8784 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 79.6262 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 355.197 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.77994 LAYER VIA7 ;
  END BIAS_DBPC[13]
  PIN BIAS_DBPC[12] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.155 LAYER M2 ;
  END BIAS_DBPC[12]
  PIN BIAS_DBPC[11] 
    ANTENNAPARTIALMETALAREA 0.023 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1012 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.992 LAYER M3 ;
  END BIAS_DBPC[11]
  PIN BIAS_DBPC[10] 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.778 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4672 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.846 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7664 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.358 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 41.2192 LAYER M6 ;
  END BIAS_DBPC[10]
  PIN BIAS_DBPC[9] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5872 LAYER M3 ;
  END BIAS_DBPC[9]
  PIN BIAS_DBPC[8] 
    ANTENNAPARTIALMETALAREA 0.0215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0946 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.438 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9712 LAYER M3 ;
  END BIAS_DBPC[8]
  PIN BIAS_DBPC[7] 
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3056 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.6833 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.39 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3 ;
  END BIAS_DBPC[7]
  PIN BIAS_DBPC[6] 
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.788 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9552 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.626 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 11.5984 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.56 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 20.152 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 219.838 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 969.336 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_DBPC[6]
  PIN BIAS_DBPC[5] 
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.478 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.3472 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 LAYER M4 ; 
    ANTENNAMAXAREACAR 42.1301 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 186.866 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.514403 LAYER VIA4 ;
  END BIAS_DBPC[5]
  PIN BIAS_DBPC[4] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.5065 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3166 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.438 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3712 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ; 
    ANTENNAMAXAREACAR 47.5717 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 212.557 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.0929 LAYER VIA4 ;
  END BIAS_DBPC[4]
  PIN BIAS_DBPC[3] 
    ANTENNAPARTIALMETALAREA 0.019 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0836 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6528 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.998 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4352 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.484 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 50.6176 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 314.239 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1384.7 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_DBPC[3]
  PIN BIAS_DBPC[2] 
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.682 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.158 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.3392 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ; 
    ANTENNAMAXAREACAR 340.717 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1502.42 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.73224 LAYER VIA6 ;
  END BIAS_DBPC[2]
  PIN BIAS_DBPC[1] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.926 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1184 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.178 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.202 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 9.7328 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.58 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 46.64 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 578.04 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2534.76 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.23625 LAYER VIA6 ;
  END BIAS_DBPC[1]
  PIN BIAS_DBPC[0] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.3795 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7138 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.562 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 37.7168 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.104 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 18.1456 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 194.297 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 856.332 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_DBPC[0]
  PIN BIAS_DBNC[13] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.968 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.778 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.0672 LAYER M4 ;
  END BIAS_DBNC[13]
  PIN BIAS_DBNC[12] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.7275 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.645 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.498 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 37.4352 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 159.208 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 704.133 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA6 ;
  END BIAS_DBNC[12]
  PIN BIAS_DBNC[11] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.3968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.222 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.6208 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 469.544 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2071.48 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6 ;
  END BIAS_DBNC[11]
  PIN BIAS_DBNC[10] 
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.638 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 38.0512 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 149.425 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 660.45 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA4 ;
  END BIAS_DBNC[10]
  PIN BIAS_DBNC[9] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 6.576 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.0224 LAYER M2 ;
  END BIAS_DBNC[9]
  PIN BIAS_DBNC[8] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.882 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.7248 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.078 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.0752 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 405.272 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1791.53 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.589 LAYER VIA6 ;
  END BIAS_DBNC[8]
  PIN BIAS_DBNC[7] 
    ANTENNAPARTIALMETALAREA 0.808 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5992 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.296 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.4784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 179.188 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 793.916 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3 ;
  END BIAS_DBNC[7]
  PIN BIAS_DBNC[6] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.864 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.1898 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 152.877 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.411523 LAYER VIA3 ;
  END BIAS_DBNC[6]
  PIN BIAS_DBNC[5] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.645 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.282 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.0512 LAYER M4 ;
  END BIAS_DBNC[5]
  PIN BIAS_DBNC[4] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.396 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.1184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ; 
    ANTENNAMAXAREACAR 97.862 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 434.301 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.819672 LAYER VIA3 ;
  END BIAS_DBNC[4]
  PIN BIAS_DBNC[3] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.618 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 24.7632 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 102.873 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 454.355 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA4 ;
  END BIAS_DBNC[3]
  PIN BIAS_DBNC[2] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.0215 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3826 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M3 ; 
    ANTENNAMAXAREACAR 135.075 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 597.675 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.617284 LAYER VIA3 ;
  END BIAS_DBNC[2]
  PIN BIAS_DBNC[1] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.503 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2572 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.326 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8784 LAYER M5 ;
  END BIAS_DBNC[1]
  PIN BIAS_DBNC[0] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4784 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4512 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 62.0653 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 275.434 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA4 ;
  END BIAS_DBNC[0]
  PIN BIAS_TC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.2055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9042 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3 ;
  END BIAS_TC_POT[5]
  PIN BIAS_TC_POT[4] 
    ANTENNAPARTIALMETALAREA 0.151 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6644 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
  END BIAS_TC_POT[4]
  PIN BIAS_TC_POT[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.891 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
  END BIAS_TC_POT[3]
  PIN BIAS_TC_POT[2] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.108 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.1632 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ; 
    ANTENNAMAXAREACAR 118.829 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 526.087 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.819672 LAYER VIA3 ;
  END BIAS_TC_POT[2]
  PIN BIAS_TC_POT[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.664 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0096 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.438 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9712 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.142 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0688 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 33.7767 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 151.036 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA5 ;
  END BIAS_TC_POT[1]
  PIN BIAS_TC_POT[0] 
    ANTENNAPARTIALMETALAREA 0.118 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5192 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.126 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.7984 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.578 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.7872 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 79.4679 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 352.006 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA5 ;
  END BIAS_TC_POT[0]
  PIN BIAS_LC_POT[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.9995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4858 LAYER M2 ;
  END BIAS_LC_POT[5]
  PIN BIAS_LC_POT[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.738 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2912 LAYER M2 ;
  END BIAS_LC_POT[4]
  PIN BIAS_LC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.9535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1954 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.658 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9392 LAYER M3 ;
  END BIAS_LC_POT[3]
  PIN BIAS_LC_POT[2] 
    ANTENNAPARTIALMETALAREA 0.575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.53 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.046 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6464 LAYER M3 ;
  END BIAS_LC_POT[2]
  PIN BIAS_LC_POT[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4034 LAYER M2 ;
  END BIAS_LC_POT[1]
  PIN BIAS_LC_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.468 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1032 LAYER M2 ;
  END BIAS_LC_POT[0]
  PIN BIAS_TIA_G_POT[16] 
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M3 ;
  END BIAS_TIA_G_POT[16]
  PIN BIAS_TIA_G_POT[15] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7015 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0866 LAYER M2 ;
  END BIAS_TIA_G_POT[15]
  PIN BIAS_TIA_G_POT[14] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.329 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4916 LAYER M2 ;
  END BIAS_TIA_G_POT[14]
  PIN BIAS_TIA_G_POT[13] 
    ANTENNAPARTIALMETALAREA 0.7495 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2978 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7728 LAYER M3 ;
  END BIAS_TIA_G_POT[13]
  PIN BIAS_TIA_G_POT[12] 
    ANTENNAPARTIALMETALAREA 0.117 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5148 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.338 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M5 ;
  END BIAS_TIA_G_POT[12]
  PIN BIAS_TIA_G_POT[11] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.691 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2 ;
  END BIAS_TIA_G_POT[11]
  PIN BIAS_TIA_G_POT[10] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.342 LAYER M2 ;
  END BIAS_TIA_G_POT[10]
  PIN BIAS_TIA_G_POT[9] 
    ANTENNAPARTIALMETALAREA 0.6345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7918 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.978 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3472 LAYER M3 ;
  END BIAS_TIA_G_POT[9]
  PIN BIAS_TIA_G_POT[8] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.471 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0724 LAYER M2 ;
  END BIAS_TIA_G_POT[8]
  PIN BIAS_TIA_G_POT[7] 
    ANTENNAPARTIALMETALAREA 0.3525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.551 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.226 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.2384 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.142 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 6.478 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 28.5472 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0447 LAYER M5 ; 
    ANTENNAMAXAREACAR 264.498 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1167.52 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.78971 LAYER VIA5 ;
  END BIAS_TIA_G_POT[7]
  PIN BIAS_TIA_G_POT[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.509 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6836 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.918 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.4832 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.538 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 28.8112 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 6.358 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 28.0192 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 28.024 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 123.482 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 441.914 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1949.31 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6 ;
  END BIAS_TIA_G_POT[6]
  PIN BIAS_TIA_G_POT[5] 
    ANTENNAPARTIALMETALAREA 0.1725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.759 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.902 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0128 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 21.964 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 96.7296 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ; 
    ANTENNAMAXAREACAR 734.195 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 3226.68 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.91257 LAYER VIA5 ;
  END BIAS_TIA_G_POT[5]
  PIN BIAS_TIA_G_POT[4] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.061 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3124 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.442 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7888 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 30.446 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 134.006 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.122 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 58.6815 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 261.815 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6 ;
  END BIAS_TIA_G_POT[4]
  PIN BIAS_TIA_G_POT[3] 
    ANTENNAPARTIALMETALAREA 1.3145 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7838 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.9728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.462 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.2768 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 90.4058 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 400.768 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA5 ;
  END BIAS_TIA_G_POT[3]
  PIN BIAS_TIA_G_POT[2] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.956 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6504 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.868 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.3072 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 140.651 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 621.847 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA4 ;
  END BIAS_TIA_G_POT[2]
  PIN BIAS_TIA_G_POT[1] 
    ANTENNAPARTIALMETALAREA 0.051 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2244 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.378 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5072 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.226 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4384 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 6.918 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 30.4832 LAYER M5 ;
  END BIAS_TIA_G_POT[1]
  PIN BIAS_TIA_G_POT[0] 
    ANTENNAPARTIALMETALAREA 0.151 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6644 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.698 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.9152 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.586 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6224 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 6.498 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 28.7232 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.646 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8864 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 18.4289 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 84.0693 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6 ;
  END BIAS_TIA_G_POT[0]
  PIN BIAS_REV_POT[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.563 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.0772 LAYER M2 ;
  END BIAS_REV_POT[13]
  PIN BIAS_REV_POT[12] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.318 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4432 LAYER M3 ;
  END BIAS_REV_POT[12]
  PIN BIAS_REV_POT[11] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
  END BIAS_REV_POT[11]
  PIN BIAS_REV_POT[10] 
    ANTENNAPARTIALMETALAREA 1.0455 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3 ;
  END BIAS_REV_POT[10]
  PIN BIAS_REV_POT[9] 
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.564 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5696 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.878 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9072 LAYER M4 ;
  END BIAS_REV_POT[9]
  PIN BIAS_REV_POT[8] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.428 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9712 LAYER M3 ;
  END BIAS_REV_POT[8]
  PIN BIAS_REV_POT[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
  END BIAS_REV_POT[7]
  PIN BIAS_REV_POT[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0265 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1606 LAYER M2 ;
  END BIAS_REV_POT[6]
  PIN BIAS_REV_POT[5] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.298 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3552 LAYER M3 ;
  END BIAS_REV_POT[5]
  PIN BIAS_REV_POT[4] 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.942 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1888 LAYER M4 ;
  END BIAS_REV_POT[4]
  PIN BIAS_REV_POT[3] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_REV_POT[3]
  PIN BIAS_REV_POT[2] 
    ANTENNAPARTIALMETALAREA 0.5225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.299 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3968 LAYER M3 ;
  END BIAS_REV_POT[2]
  PIN BIAS_REV_POT[1] 
    ANTENNAPARTIALMETALAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3256 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3408 LAYER M3 ;
  END BIAS_REV_POT[1]
  PIN BIAS_REV_POT[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3498 LAYER M2 ;
  END BIAS_REV_POT[0]
  PIN BIAS_TC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.771 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.162 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M4 ;
  END BIAS_TC_DSADC[5]
  PIN BIAS_TC_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.131 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5764 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.401 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8084 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.746 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3264 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.018 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5232 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.206 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 164.517 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 728.457 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_TC_DSADC[4]
  PIN BIAS_TC_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3506 LAYER M2 ;
  END BIAS_TC_DSADC[3]
  PIN BIAS_TC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.891 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9204 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.562 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5168 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 7.138 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 31.4512 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 140.429 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 619.212 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA5 ;
  END BIAS_TC_DSADC[2]
  PIN BIAS_TC_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.2105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9262 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.786 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5024 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 6.958 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 30.6592 LAYER M5 ;
  END BIAS_TC_DSADC[1]
  PIN BIAS_TC_DSADC[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.528 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3232 LAYER M2 ;
  END BIAS_TC_DSADC[0]
  PIN BIAS_LC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.6315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7786 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.378 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1072 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 8.662 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 38.1568 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.182 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 104.176 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 461.832 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.23625 LAYER VIA6 ;
  END BIAS_LC_DSADC[5]
  PIN BIAS_LC_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.131 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5764 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.678 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0272 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.698 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.7152 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.126 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 173.755 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 768.265 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.23625 LAYER VIA6 ;
  END BIAS_LC_DSADC[4]
  PIN BIAS_LC_DSADC[3] 
    ANTENNAPARTIALMETALAREA 1.1715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1546 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5648 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.522 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3408 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 8.656 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 38.1744 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 159.135 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 702.294 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA5 ;
  END BIAS_LC_DSADC[3]
  PIN BIAS_LC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 1.386 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0984 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 6.618 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 29.1632 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 150.285 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 661.838 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA5 ;
  END BIAS_LC_DSADC[2]
  PIN BIAS_LC_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.5405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.002 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6528 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.662 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 16.1568 LAYER M5 ;
  END BIAS_LC_DSADC[1]
  PIN BIAS_LC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.131 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6204 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.438 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9712 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.106 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9104 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 7.018 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 30.9232 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 133.604 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 588.857 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA5 ;
  END BIAS_LC_DSADC[0]
  PIN BIAS_RIN_DSADC[5] 
    ANTENNAPARTIALMETALAREA 1.0285 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5254 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.638 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.6512 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.186 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 6.678 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 29.4272 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M5 ; 
    ANTENNAMAXAREACAR 301.841 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1332.17 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.26537 LAYER VIA5 ;
  END BIAS_RIN_DSADC[5]
  PIN BIAS_RIN_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.383 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6852 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.866 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8544 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.264 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2496 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.202 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.5328 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.206 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 152.974 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 680 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6 ;
  END BIAS_RIN_DSADC[4]
  PIN BIAS_RIN_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.191 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8404 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0676 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.244 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9616 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 8.738 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 38.4912 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 175.919 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 771.592 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.13269 LAYER VIA5 ;
  END BIAS_RIN_DSADC[3]
  PIN BIAS_RIN_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.398 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.7952 LAYER M3 ;
  END BIAS_RIN_DSADC[2]
  PIN BIAS_RIN_DSADC[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1902 LAYER M2 ;
  END BIAS_RIN_DSADC[1]
  PIN BIAS_RIN_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.118 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5192 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.338 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.146 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0864 LAYER M5 ;
  END BIAS_RIN_DSADC[0]
  PIN BIAS_RFB_DSADC[5] 
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.3325 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.507 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.458 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.466 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0944 LAYER M4 ;
  END BIAS_RFB_DSADC[5]
  PIN BIAS_RFB_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.157 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6908 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5008 LAYER M3 ;
  END BIAS_RFB_DSADC[4]
  PIN BIAS_RFB_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.091 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1545 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7238 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.686 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0624 LAYER M4 ;
  END BIAS_RFB_DSADC[3]
  PIN BIAS_RFB_DSADC[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.649 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8996 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.802 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.866 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8544 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.22 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 5.456 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 2.866 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6544 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M7 ; 
    ANTENNAMAXAREACAR 581.1 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 2564.19 LAYER M7 ;
    ANTENNAMAXCUTCAR 3.8835 LAYER VIA7 ;
  END BIAS_RFB_DSADC[2]
  PIN BIAS_RFB_DSADC[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.9565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2526 LAYER M2 ;
  END BIAS_RFB_DSADC[1]
  PIN BIAS_RFB_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.937 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1228 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.162 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1568 LAYER M3 ;
  END BIAS_RFB_DSADC[0]
  PIN BIAS_DSADC_VCM[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.975 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.934 LAYER M2 ;
  END BIAS_DSADC_VCM[13]
  PIN BIAS_DSADC_VCM[12] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.598 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6752 LAYER M4 ;
  END BIAS_DSADC_VCM[12]
  PIN BIAS_DSADC_VCM[11] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.848 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7752 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.858 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8192 LAYER M4 ;
  END BIAS_DSADC_VCM[11]
  PIN BIAS_DSADC_VCM[10] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3408 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.006 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4704 LAYER M4 ;
  END BIAS_DSADC_VCM[10]
  PIN BIAS_DSADC_VCM[9] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.882 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9248 LAYER M4 ;
  END BIAS_DSADC_VCM[9]
  PIN BIAS_DSADC_VCM[8] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.2165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.1526 LAYER M2 ;
  END BIAS_DSADC_VCM[8]
  PIN BIAS_DSADC_VCM[7] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.558 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4992 LAYER M4 ;
  END BIAS_DSADC_VCM[7]
  PIN BIAS_DSADC_VCM[6] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8766 LAYER M2 ;
  END BIAS_DSADC_VCM[6]
  PIN BIAS_DSADC_VCM[5] 
    ANTENNAPARTIALMETALAREA 0.073 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3212 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3968 LAYER M3 ;
  END BIAS_DSADC_VCM[5]
  PIN BIAS_DSADC_VCM[4] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8048 LAYER M3 ;
  END BIAS_DSADC_VCM[4]
  PIN BIAS_DSADC_VCM[3] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.138 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6512 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.982 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3648 LAYER M4 ;
  END BIAS_DSADC_VCM[3]
  PIN BIAS_DSADC_VCM[2] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3968 LAYER M3 ;
  END BIAS_DSADC_VCM[2]
  PIN BIAS_DSADC_VCM[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.308 LAYER M2 ;
  END BIAS_DSADC_VCM[1]
  PIN BIAS_DSADC_VCM[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.099 LAYER M2 ;
  END BIAS_DSADC_VCM[0]
  PIN dsadc_conv_done 
    ANTENNAPARTIALMETALAREA 0.806 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.138 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0512 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 7.978 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 35.1472 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.718 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2032 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0269 LAYER M6 ; 
    ANTENNAMAXAREACAR 408.487 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1804.16 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.34572 LAYER VIA6 ;
  END dsadc_conv_done
  PIN dsadc_en 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.506 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2264 LAYER M2 ;
  END dsadc_en
  PIN dsadc_clk 
    ANTENNAPARTIALMETALAREA 0.196 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2156 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 30.002 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.1782 LAYER M3 ;
  END dsadc_clk
  PIN dsadc_switch[2] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1858 LAYER M2 ;
  END dsadc_switch[2]
  PIN dsadc_switch[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.474 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0856 LAYER M2 ;
  END dsadc_switch[1]
  PIN dsadc_switch[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3046 LAYER M2 ;
  END dsadc_switch[0]
  PIN dac_en_pot 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1902 LAYER M2 ;
  END dac_en_pot
  PIN adc_ext_in 
    ANTENNAPARTIALMETALAREA 0.151 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6644 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M3 ;
  END adc_ext_in
  PIN atp_en 
    ANTENNAPARTIALMETALAREA 0.3045 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.882 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9248 LAYER M3 ;
  END atp_en
  PIN atp_sel 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.381 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7204 LAYER M2 ;
  END atp_sel
  PIN adc_sel 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4002 LAYER M2 ;
  END adc_sel
  PIN saradc_clk 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 67.982 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 74.9562 LAYER M3 ;
  END saradc_clk
  PIN saradc_rdy 
    ANTENNAPARTIALMETALAREA 0.167 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7348 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.0015 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4506 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.702 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1328 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.538 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.0112 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M5 ; 
    ANTENNAMAXAREACAR 350.48 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1534.17 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.95203 LAYER VIA5 ;
  END saradc_rdy
  PIN saradc_rst 
    ANTENNAPARTIALMETALAREA 1.0825 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.763 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.0608 LAYER M3 ;
  END saradc_rst
  PIN saradc_data[9] 
    ANTENNAPARTIALMETALAREA 0.5485 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 8.638 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.0512 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 330.494 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1440.89 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[9]
  PIN saradc_data[8] 
    ANTENNAPARTIALMETALAREA 0.8825 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.883 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 8.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.2208 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 340.664 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1489.59 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[8]
  PIN saradc_data[7] 
    ANTENNAPARTIALMETALAREA 0.431 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8964 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.1335 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.2314 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 371.125 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1625.48 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[7]
  PIN saradc_data[6] 
    ANTENNAPARTIALMETALAREA 0.7665 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3726 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 8.178 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.0272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 351.587 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1532.34 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[6]
  PIN saradc_data[5] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0975 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.473 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.346 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9664 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M4 ; 
    ANTENNAMAXAREACAR 417.343 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1833.39 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.21402 LAYER VIA4 ;
  END saradc_data[5]
  PIN saradc_data[4] 
    ANTENNAPARTIALMETALAREA 0.3575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.178 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.6716 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.8561 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[4]
  PIN saradc_data[3] 
    ANTENNAPARTIALMETALAREA 0.9225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.059 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 8.186 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.0624 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 359.779 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1568.12 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[3]
  PIN saradc_data[2] 
    ANTENNAPARTIALMETALAREA 0.5825 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.563 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 8.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.5408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 332.399 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1458.54 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[2]
  PIN saradc_data[1] 
    ANTENNAPARTIALMETALAREA 0.6425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.827 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 7.898 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.7952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 325.107 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1408.41 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[1]
  PIN saradc_data[0] 
    ANTENNAPARTIALMETALAREA 0.8025 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.531 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.9968 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 370.554 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1630.94 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[0]
END MCU

END LIBRARY
