

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO MCU 
  PIN resetn_in 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 26.022 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 114.541 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6 ; 
    ANTENNAMAXAREACAR 974.013 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4292.32 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.32103 LAYER VIA6 ;
  END resetn_in
  PIN resetn_out 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.562 LAYER M2 ;
  END resetn_out
  PIN resetn_dir 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6654 LAYER M2 ;
  END resetn_dir
  PIN resetn_ren 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5895 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6378 LAYER M2 ;
  END resetn_ren
  PIN prt1_in[7] 
    ANTENNAPARTIALMETALAREA 21.3345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 93.9158 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.682 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.2448 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 198.303 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 858.686 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt1_in[7]
  PIN prt1_in[6] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.682 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.8448 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0269 LAYER M3 ; 
    ANTENNAMAXAREACAR 105.104 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 463.859 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.48699 LAYER VIA3 ;
  END prt1_in[6]
  PIN prt1_in[5] 
    ANTENNAPARTIALMETALAREA 9.9325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 43.703 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 6.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.6848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 248.892 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1095.53 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END prt1_in[5]
  PIN prt1_in[4] 
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.796 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3904 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2577 LAYER M4 ; 
    ANTENNAMAXAREACAR 223.702 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 986.113 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.09268 LAYER VIA4 ;
  END prt1_in[4]
  PIN prt1_in[3] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6182 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.402 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6182 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.68 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.424 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 LAYER M5 ; 
    ANTENNAMAXAREACAR 55.9025 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 65.8857 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.10063 LAYER VIA5 ;
  END prt1_in[3]
  PIN prt1_in[2] 
    ANTENNAPARTIALMETALAREA 0.5355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3562 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 15.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 69.872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1931 LAYER M3 ; 
    ANTENNAMAXAREACAR 111.068 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 488.742 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.895857 LAYER VIA3 ;
  END prt1_in[2]
  PIN prt1_in[1] 
    ANTENNAPARTIALMETALAREA 13.5175 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.521 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.1888 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3 ; 
    ANTENNAMAXAREACAR 65.9383 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 282.417 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3 ;
  END prt1_in[1]
  PIN prt1_in[0] 
    ANTENNAPARTIALMETALAREA 23.1955 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 102.06 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.3248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3 ; 
    ANTENNAMAXAREACAR 62.722 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 275.441 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3 ;
  END prt1_in[0]
  PIN prt1_out[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2 ;
  END prt1_out[7]
  PIN prt1_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.337 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.8148 LAYER M2 ;
  END prt1_out[6]
  PIN prt1_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[5]
  PIN prt1_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.041 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2244 LAYER M2 ;
  END prt1_out[4]
  PIN prt1_out[3] 
    ANTENNAPARTIALMETALAREA 1.336 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8784 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.062 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.5168 LAYER M3 ;
  END prt1_out[3]
  PIN prt1_out[2] 
    ANTENNAPARTIALMETALAREA 0.036 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1584 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3 ;
  END prt1_out[2]
  PIN prt1_out[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[1]
  PIN prt1_out[0] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2 ;
  END prt1_out[0]
  PIN prt1_dir[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[7]
  PIN prt1_dir[6] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
  END prt1_dir[6]
  PIN prt1_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2 ;
  END prt1_dir[5]
  PIN prt1_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1455 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6842 LAYER M2 ;
  END prt1_dir[4]
  PIN prt1_dir[3] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[3]
  PIN prt1_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2142 LAYER M2 ;
  END prt1_dir[2]
  PIN prt1_dir[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[1]
  PIN prt1_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.9345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 52.5998 LAYER M2 ;
  END prt1_dir[0]
  PIN prt1_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.1235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.0314 LAYER M2 ;
  END prt1_ren[7]
  PIN prt1_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.3835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.9754 LAYER M2 ;
  END prt1_ren[6]
  PIN prt1_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 15.8235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 69.7114 LAYER M2 ;
  END prt1_ren[5]
  PIN prt1_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M2 ;
  END prt1_ren[4]
  PIN prt1_ren[3] 
    ANTENNAPARTIALMETALAREA 0.3075 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.353 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.9488 LAYER M3 ;
  END prt1_ren[3]
  PIN prt1_ren[2] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.9136 LAYER M3 ;
  END prt1_ren[2]
  PIN prt1_ren[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.5505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 50.9102 LAYER M2 ;
  END prt1_ren[1]
  PIN prt1_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.2145 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 53.8318 LAYER M2 ;
  END prt1_ren[0]
  PIN prt2_in[7] 
    ANTENNAPARTIALMETALAREA 0.7775 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.465 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 LAYER M2 ; 
    ANTENNAMAXAREACAR 7.94537 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 34.5167 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.185185 LAYER VIA2 ;
  END prt2_in[7]
  PIN prt2_in[6] 
    ANTENNAPARTIALMETALAREA 0.4975 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.233 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2 ; 
    ANTENNAMAXAREACAR 17.7666 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 77.1643 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2 ;
  END prt2_in[6]
  PIN prt2_in[5] 
    ANTENNAPARTIALMETALAREA 0.7125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.135 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2 ; 
    ANTENNAMAXAREACAR 6.69969 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 28.5519 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA2 ;
  END prt2_in[5]
  PIN prt2_in[4] 
    ANTENNAPARTIALMETALAREA 0.7595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3418 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.3088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 329.539 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1444.21 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt2_in[4]
  PIN prt2_in[3] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3916 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.64 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 LAYER M4 ; 
    ANTENNAMAXAREACAR 14.9049 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 19.2925 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.235849 LAYER VIA4 ;
  END prt2_in[3]
  PIN prt2_in[2] 
    ANTENNAPARTIALMETALAREA 0.6599 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6026 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 31.158 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 137.139 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 926.784 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4059.66 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt2_in[2]
  PIN prt2_in[1] 
    ANTENNAPARTIALMETALAREA 0.3355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4762 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 27.346 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 120.366 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0381 LAYER M3 ; 
    ANTENNAMAXAREACAR 732.747 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3223.46 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.04987 LAYER VIA3 ;
  END prt2_in[1]
  PIN prt2_in[0] 
    ANTENNAPARTIALMETALAREA 0.3535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5994 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2 ; 
    ANTENNAMAXAREACAR 5.43396 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 22.706 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA2 ;
  END prt2_in[0]
  PIN prt2_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.701 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1284 LAYER M2 ;
  END prt2_out[7]
  PIN prt2_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.681 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2 ;
  END prt2_out[6]
  PIN prt2_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.234 LAYER M2 ;
  END prt2_out[5]
  PIN prt2_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.297 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3508 LAYER M2 ;
  END prt2_out[4]
  PIN prt2_out[3] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.914 LAYER M2 ;
  END prt2_out[3]
  PIN prt2_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.554 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4816 LAYER M2 ;
  END prt2_out[2]
  PIN prt2_out[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.279 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2276 LAYER M2 ;
  END prt2_out[1]
  PIN prt2_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.512 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M2 ;
  END prt2_out[0]
  PIN prt2_dir[7] 
    ANTENNAPARTIALMETALAREA 0.691 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5968 LAYER M3 ;
  END prt2_dir[7]
  PIN prt2_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.8005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5662 LAYER M2 ;
  END prt2_dir[6]
  PIN prt2_dir[5] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M2 ;
  END prt2_dir[5]
  PIN prt2_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6765 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0206 LAYER M2 ;
  END prt2_dir[4]
  PIN prt2_dir[3] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1946 LAYER M2 ;
  END prt2_dir[3]
  PIN prt2_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3706 LAYER M2 ;
  END prt2_dir[2]
  PIN prt2_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M2 ;
  END prt2_dir[1]
  PIN prt2_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3166 LAYER M2 ;
  END prt2_dir[0]
  PIN prt2_ren[7] 
    ANTENNAPARTIALMETALAREA 0.6435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8314 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.582 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8048 LAYER M3 ;
  END prt2_ren[7]
  PIN prt2_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.299 LAYER M2 ;
  END prt2_ren[6]
  PIN prt2_ren[5] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.639 LAYER M2 ;
  END prt2_ren[5]
  PIN prt2_ren[4] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5275 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.409 LAYER M2 ;
  END prt2_ren[4]
  PIN prt2_ren[3] 
    ANTENNAPARTIALMETALAREA 0.5305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3342 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.918 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.8832 LAYER M3 ;
  END prt2_ren[3]
  PIN prt2_ren[2] 
    ANTENNAPARTIALMETALAREA 0.887 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9028 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.0495 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.4618 LAYER M3 ;
  END prt2_ren[2]
  PIN prt2_ren[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2078 LAYER M2 ;
  END prt2_ren[1]
  PIN prt2_ren[0] 
    ANTENNAPARTIALMETALAREA 0.6875 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.025 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.4848 LAYER M3 ;
  END prt2_ren[0]
  PIN prt3_in[7] 
    ANTENNAPARTIALMETALAREA 24.9345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 109.756 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.078 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.5872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 507.616 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2214.91 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[7]
  PIN prt3_in[6] 
    ANTENNAPARTIALMETALAREA 16.1305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 71.0182 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2 ; 
    ANTENNAMAXAREACAR 596.836 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2626.24 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.369004 LAYER VIA2 ;
  END prt3_in[6]
  PIN prt3_in[5] 
    ANTENNAPARTIALMETALAREA 7.5705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.3542 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.71 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 151.946 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 669.018 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.08401 LAYER VIA3 ;
  END prt3_in[5]
  PIN prt3_in[4] 
    ANTENNAPARTIALMETALAREA 0.1155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5082 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 8.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.5904 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.378 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.7072 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M5 ; 
    ANTENNAMAXAREACAR 65.5619 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 285.971 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.12004 LAYER VIA5 ;
  END prt3_in[4]
  PIN prt3_in[3] 
    ANTENNAPARTIALMETALAREA 4.4395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.5338 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 18.864 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 83.0896 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1707 LAYER M3 ; 
    ANTENNAMAXAREACAR 143.68 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 633.441 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA3 ;
  END prt3_in[3]
  PIN prt3_in[2] 
    ANTENNAPARTIALMETALAREA 6.0735 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.7674 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.078 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.5872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 510.273 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2225.54 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[2]
  PIN prt3_in[1] 
    ANTENNAPARTIALMETALAREA 14.5735 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 64.1674 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.622 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.3808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 409.594 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1802.45 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[1]
  PIN prt3_in[0] 
    ANTENNAPARTIALMETALAREA 1.8905 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.3622 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 8.118 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.7632 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 265.401 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1148.54 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt3_in[0]
  PIN prt3_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 66.154 LAYER M2 ;
  END prt3_out[7]
  PIN prt3_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 6.359 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.0676 LAYER M2 ;
  END prt3_out[6]
  PIN prt3_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.137 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6468 LAYER M2 ;
  END prt3_out[5]
  PIN prt3_out[4] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.261 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1924 LAYER M2 ;
  END prt3_out[4]
  PIN prt3_out[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.137 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6468 LAYER M2 ;
  END prt3_out[3]
  PIN prt3_out[2] 
    ANTENNAPARTIALMETALAREA 3.69 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.28 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.162 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.3568 LAYER M3 ;
  END prt3_out[2]
  PIN prt3_out[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.202 LAYER M2 ;
  END prt3_out[1]
  PIN prt3_out[0] 
    ANTENNAPARTIALMETALAREA 1.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.664 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.086 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8224 LAYER M4 ;
  END prt3_out[0]
  PIN prt3_dir[7] 
    ANTENNAPARTIALMETALAREA 0.9995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3978 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.336 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6104 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.478 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1472 LAYER M4 ;
  END prt3_dir[7]
  PIN prt3_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 8.4095 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 37.1338 LAYER M2 ;
  END prt3_dir[6]
  PIN prt3_dir[5] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.686 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4624 LAYER M3 ;
  END prt3_dir[5]
  PIN prt3_dir[4] 
    ANTENNAPARTIALMETALAREA 0.3965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7446 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.898 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.9952 LAYER M3 ;
  END prt3_dir[4]
  PIN prt3_dir[3] 
    ANTENNAPARTIALMETALAREA 0.9915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3626 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.008 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.5232 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.698 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1152 LAYER M4 ;
  END prt3_dir[3]
  PIN prt3_dir[2] 
    ANTENNAPARTIALMETALAREA 1.0715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7146 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.118 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M3 ;
  END prt3_dir[2]
  PIN prt3_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.9325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.435 LAYER M2 ;
  END prt3_dir[1]
  PIN prt3_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.8875 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.793 LAYER M2 ;
  END prt3_dir[0]
  PIN prt3_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.3255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.7642 LAYER M2 ;
  END prt3_ren[7]
  PIN prt3_ren[6] 
    ANTENNAPARTIALMETALAREA 5.406 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.8304 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2368 LAYER M3 ;
  END prt3_ren[6]
  PIN prt3_ren[5] 
    ANTENNAPARTIALMETALAREA 0.5805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5542 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.184 LAYER M3 ;
  END prt3_ren[5]
  PIN prt3_ren[4] 
    ANTENNAPARTIALMETALAREA 0.5405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.144 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.1216 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0582 LAYER M3 ; 
    ANTENNAMAXAREACAR 198.304 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 871.869 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.687285 LAYER VIA3 ;
  END prt3_ren[4]
  PIN prt3_ren[3] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.548 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.8992 LAYER M3 ;
  END prt3_ren[3]
  PIN prt3_ren[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 8.9125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 39.347 LAYER M2 ;
  END prt3_ren[2]
  PIN prt3_ren[1] 
    ANTENNAPARTIALMETALAREA 11.3205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.8102 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.1568 LAYER M3 ;
  END prt3_ren[1]
  PIN prt3_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.5255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2442 LAYER M2 ;
  END prt3_ren[0]
  PIN prt4_in[7] 
    ANTENNAPARTIALMETALAREA 2.4955 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.9802 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 18.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 82.5088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 8.582 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 37.8048 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 4.558 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 20.0992 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M6 ; 
    ANTENNAMAXAREACAR 76.8125 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 332.355 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.71003 LAYER VIA6 ;
  END prt4_in[7]
  PIN prt4_in[6] 
    ANTENNAPARTIALMETALAREA 1.5355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7562 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 19.07 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.04 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 190.873 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 841.845 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA3 ;
  END prt4_in[6]
  PIN prt4_in[5] 
    ANTENNAPARTIALMETALAREA 2.8755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6522 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.0688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 115.758 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 509.971 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA3 ;
  END prt4_in[5]
  PIN prt4_in[4] 
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 6.398 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 28.1952 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1456 LAYER M4 ; 
    ANTENNAMAXAREACAR 63.4771 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 280.938 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.49238 LAYER VIA4 ;
  END prt4_in[4]
  PIN prt4_in[3] 
    ANTENNAPARTIALMETALAREA 7.5285 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.2134 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1456 LAYER M2 ; 
    ANTENNAMAXAREACAR 53.3995 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 234.539 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.271003 LAYER VIA2 ;
  END prt4_in[3]
  PIN prt4_in[2] 
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 12.432 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.7888 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 123.595 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 544.031 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA3 ;
  END prt4_in[2]
  PIN prt4_in[1] 
    ANTENNAPARTIALMETALAREA 0.731 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 21.664 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 95.4096 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 412.611 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1817.07 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA3 ;
  END prt4_in[1]
  PIN prt4_in[0] 
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.8528 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 15.802 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 69.5728 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M6 ; 
    ANTENNAMAXAREACAR 476.628 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2101.44 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.88184 LAYER VIA6 ;
  END prt4_in[0]
  PIN prt4_out[7] 
    ANTENNAPARTIALMETALAREA 10.652 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.7766 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 48.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.592 LAYER M3 ;
  END prt4_out[7]
  PIN prt4_out[6] 
    ANTENNAPARTIALMETALAREA 8.492 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4006 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 32.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.728 LAYER M3 ;
  END prt4_out[6]
  PIN prt4_out[5] 
    ANTENNAPARTIALMETALAREA 0.172 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 18.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.5062 LAYER M3 ;
  END prt4_out[5]
  PIN prt4_out[4] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7382 LAYER M3 ;
  END prt4_out[4]
  PIN prt4_out[3] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.4912 LAYER M3 ;
  END prt4_out[3]
  PIN prt4_out[2] 
    ANTENNAPARTIALMETALAREA 0.499 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1956 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.722 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.8208 LAYER M3 ;
  END prt4_out[2]
  PIN prt4_out[1] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.962 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 74.6768 LAYER M6 ;
  END prt4_out[1]
  PIN prt4_out[0] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
  END prt4_out[0]
  PIN prt4_dir[7] 
    ANTENNAPARTIALMETALAREA 0.2915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.546 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.8464 LAYER M3 ;
  END prt4_dir[7]
  PIN prt4_dir[6] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2765 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2606 LAYER M2 ;
  END prt4_dir[6]
  PIN prt4_dir[5] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3222 LAYER M2 ;
  END prt4_dir[5]
  PIN prt4_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.5585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9014 LAYER M2 ;
  END prt4_dir[4]
  PIN prt4_dir[3] 
    ANTENNAPARTIALMETALAREA 0.871 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.898 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.5952 LAYER M3 ;
  END prt4_dir[3]
  PIN prt4_dir[2] 
    ANTENNAPARTIALMETALAREA 0.2965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3046 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.666 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.1744 LAYER M3 ;
  END prt4_dir[2]
  PIN prt4_dir[1] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.722 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.6208 LAYER M6 ;
  END prt4_dir[1]
  PIN prt4_dir[0] 
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 15.942 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 70.1888 LAYER M6 ;
  END prt4_dir[0]
  PIN prt4_ren[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2286 LAYER M2 ;
  END prt4_ren[7]
  PIN prt4_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5825 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.607 LAYER M2 ;
  END prt4_ren[6]
  PIN prt4_ren[5] 
    ANTENNAPARTIALMETALAREA 1.2705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.906 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.8304 LAYER M3 ;
  END prt4_ren[5]
  PIN prt4_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.7425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.711 LAYER M2 ;
  END prt4_ren[4]
  PIN prt4_ren[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.3385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.7334 LAYER M2 ;
  END prt4_ren[3]
  PIN prt4_ren[2] 
    ANTENNAPARTIALMETALAREA 0.6435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8314 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.6848 LAYER M3 ;
  END prt4_ren[2]
  PIN prt4_ren[1] 
    ANTENNAPARTIALMETALAREA 0.8035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 15.942 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 70.1888 LAYER M6 ;
  END prt4_ren[1]
  PIN prt4_ren[0] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 17.122 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 75.3808 LAYER M6 ;
  END prt4_ren[0]
  PIN use_dac_glb_bias 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4375 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.925 LAYER M2 ;
  END use_dac_glb_bias
  PIN en_bias_buf 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 6.563 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.9652 LAYER M2 ;
  END en_bias_buf
  PIN en_bias_gen 
    ANTENNAPARTIALMETALAREA 0.041 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1804 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.558 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6992 LAYER M4 ;
  END en_bias_gen
  PIN BIAS_ADJ[5] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9872 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.918 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.8832 LAYER M6 ;
  END BIAS_ADJ[5]
  PIN BIAS_ADJ[4] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
  END BIAS_ADJ[4]
  PIN BIAS_ADJ[3] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.658 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.7392 LAYER M4 ;
  END BIAS_ADJ[3]
  PIN BIAS_ADJ[2] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.262 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M4 ;
  END BIAS_ADJ[2]
  PIN BIAS_ADJ[1] 
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3 ;
  END BIAS_ADJ[1]
  PIN BIAS_ADJ[0] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.4305 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3382 LAYER M3 ;
  END BIAS_ADJ[0]
  PIN BIAS_DBP[13] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.35 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.472 LAYER M3 ;
  END BIAS_DBP[13]
  PIN BIAS_DBP[12] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3 ;
  END BIAS_DBP[12]
  PIN BIAS_DBP[11] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1648 LAYER M3 ;
  END BIAS_DBP[11]
  PIN BIAS_DBP[10] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1562 LAYER M2 ;
  END BIAS_DBP[10]
  PIN BIAS_DBP[9] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1008 LAYER M3 ;
  END BIAS_DBP[9]
  PIN BIAS_DBP[8] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.562 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9168 LAYER M3 ;
  END BIAS_DBP[8]
  PIN BIAS_DBP[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.916 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1184 LAYER M2 ;
  END BIAS_DBP[7]
  PIN BIAS_DBP[6] 
    ANTENNAPARTIALMETALAREA 0.0625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.558 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8992 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.978 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.9472 LAYER M4 ;
  END BIAS_DBP[6]
  PIN BIAS_DBP[5] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
  END BIAS_DBP[5]
  PIN BIAS_DBP[4] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
  END BIAS_DBP[4]
  PIN BIAS_DBP[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.885 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.982 LAYER M2 ;
  END BIAS_DBP[3]
  PIN BIAS_DBP[2] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.402 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M4 ;
  END BIAS_DBP[2]
  PIN BIAS_DBP[1] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.142 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M3 ;
  END BIAS_DBP[1]
  PIN BIAS_DBP[0] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.3475 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.573 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.818 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6432 LAYER M4 ;
  END BIAS_DBP[0]
  PIN BIAS_DBN[13] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 9.064 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 39.9696 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 157.168 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 692.863 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA4 ;
  END BIAS_DBN[13]
  PIN BIAS_DBN[12] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 7.2835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.1794 LAYER M2 ;
  END BIAS_DBN[12]
  PIN BIAS_DBN[11] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.324 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5136 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 6.818 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 30.0432 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.306 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 79.438 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 276.857 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA5 ;
  END BIAS_DBN[11]
  PIN BIAS_DBN[10] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.682 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 7.298 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 32.1552 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 1.068 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7872 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M7 ; 
    ANTENNAMAXAREACAR 63.9214 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 285.117 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.5873 LAYER VIA7 ;
  END BIAS_DBN[10]
  PIN BIAS_DBN[9] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.842 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7488 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.158 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.3392 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.262 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.7968 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 273.064 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1205.8 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA6 ;
  END BIAS_DBN[9]
  PIN BIAS_DBN[8] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.618 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7632 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.626 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 11.5984 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.716 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.0384 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 203.582 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 899.388 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_DBN[8]
  PIN BIAS_DBN[7] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
  END BIAS_DBN[7]
  PIN BIAS_DBN[6] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9152 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.882 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1248 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.398 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 45.7952 LAYER M6 ;
  END BIAS_DBN[6]
  PIN BIAS_DBN[5] 
    ANTENNAPARTIALMETALAREA 7.904 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.8656 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.298 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7552 LAYER M3 ;
  END BIAS_DBN[5]
  PIN BIAS_DBN[4] 
    ANTENNAPARTIALMETALAREA 0.0185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.328 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.478 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 24.1472 LAYER M4 ;
  END BIAS_DBN[4]
  PIN BIAS_DBN[3] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.9408 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.682 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4448 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 102.881 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 450.492 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA4 ;
  END BIAS_DBN[3]
  PIN BIAS_DBN[2] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1008 LAYER M3 ;
  END BIAS_DBN[2]
  PIN BIAS_DBN[1] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.178 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M3 ;
  END BIAS_DBN[1]
  PIN BIAS_DBN[0] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.678 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4272 LAYER M4 ;
  END BIAS_DBN[0]
  PIN BIAS_DBPC[13] 
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
  END BIAS_DBPC[13]
  PIN BIAS_DBPC[12] 
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
  END BIAS_DBPC[12]
  PIN BIAS_DBPC[11] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.476 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1824 LAYER M2 ;
  END BIAS_DBPC[11]
  PIN BIAS_DBPC[10] 
    ANTENNAPARTIALMETALAREA 0.1685 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7854 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.562 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9168 LAYER M3 ;
  END BIAS_DBPC[10]
  PIN BIAS_DBPC[9] 
    ANTENNAPARTIALMETALAREA 0.032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1408 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.866 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8544 LAYER M3 ;
  END BIAS_DBPC[9]
  PIN BIAS_DBPC[8] 
    ANTENNAPARTIALMETALAREA 0.1595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7458 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.466 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4944 LAYER M3 ;
  END BIAS_DBPC[8]
  PIN BIAS_DBPC[7] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.622 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.9808 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.94 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 52.624 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 301.95 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1333.16 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_DBPC[7]
  PIN BIAS_DBPC[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.8545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2038 LAYER M2 ;
  END BIAS_DBPC[6]
  PIN BIAS_DBPC[5] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.272 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2408 LAYER M3 ;
  END BIAS_DBPC[5]
  PIN BIAS_DBPC[4] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.2665 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2166 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.486 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.7824 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.518 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 41.9232 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M6 ; 
    ANTENNAMAXAREACAR 345.836 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1526.84 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VIA6 ;
  END BIAS_DBPC[4]
  PIN BIAS_DBPC[3] 
    ANTENNAPARTIALMETALAREA 0.019 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0836 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9872 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.618 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.5632 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.146 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.598 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 33.4752 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 401.328 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1770.49 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.23625 LAYER VIA6 ;
  END BIAS_DBPC[3]
  PIN BIAS_DBPC[2] 
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6528 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.258 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.738 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.0912 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 179.022 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 790.055 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_DBPC[2]
  PIN BIAS_DBPC[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.025 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.154 LAYER M2 ;
  END BIAS_DBPC[1]
  PIN BIAS_DBPC[0] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.246 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.842 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.5488 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.88 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 43.56 LAYER M6 ;
  END BIAS_DBPC[0]
  PIN BIAS_DBNC[13] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.358 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.258 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.3792 LAYER M4 ;
  END BIAS_DBNC[13]
  PIN BIAS_DBNC[12] 
    ANTENNAPARTIALMETALAREA 0.0225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.099 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.538 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 37.6112 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 165.211 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 729.911 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA4 ;
  END BIAS_DBNC[12]
  PIN BIAS_DBNC[11] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.242 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5088 LAYER M4 ;
  END BIAS_DBNC[11]
  PIN BIAS_DBNC[10] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.438 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 37.1712 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 182.498 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 806.609 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6 ;
  END BIAS_DBNC[10]
  PIN BIAS_DBNC[9] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 6.136 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.0864 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.702 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1328 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.562 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 20.1168 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 224.068 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 989.741 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA6 ;
  END BIAS_DBNC[9]
  PIN BIAS_DBNC[8] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.346 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.1664 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.738 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 47.2912 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 257.246 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1135.5 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.2987 LAYER VIA6 ;
  END BIAS_DBNC[8]
  PIN BIAS_DBNC[7] 
    ANTENNAPARTIALMETALAREA 0.248 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1352 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1648 LAYER M3 ;
  END BIAS_DBNC[7]
  PIN BIAS_DBNC[6] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.136 LAYER M3 ;
  END BIAS_DBNC[6]
  PIN BIAS_DBNC[5] 
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.198 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.9152 LAYER M4 ;
  END BIAS_DBNC[5]
  PIN BIAS_DBNC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2198 LAYER M2 ;
  END BIAS_DBNC[4]
  PIN BIAS_DBNC[3] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
  END BIAS_DBNC[3]
  PIN BIAS_DBNC[2] 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1248 LAYER M3 ;
  END BIAS_DBNC[2]
  PIN BIAS_DBNC[1] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.526 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7584 LAYER M3 ;
  END BIAS_DBNC[1]
  PIN BIAS_DBNC[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.276 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7024 LAYER M2 ;
  END BIAS_DBNC[0]
  PIN BIAS_TC_POT[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.932 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2328 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.422 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9008 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.92965 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 44.7677 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3 ;
  END BIAS_TC_POT[5]
  PIN BIAS_TC_POT[4] 
    ANTENNAPARTIALMETALAREA 0.063 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2772 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.698 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5152 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.15 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 28.876 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 127.142 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.122 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 100.725 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 444.912 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_TC_POT[4]
  PIN BIAS_TC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.1145 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5038 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 51.5008 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 227.49 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3 ;
  END BIAS_TC_POT[3]
  PIN BIAS_TC_POT[2] 
    ANTENNAPARTIALMETALAREA 0.651 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9084 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M2 ; 
    ANTENNAMAXAREACAR 11.6842 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 51.5633 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.333333 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.178 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M3 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.6508 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 65.35 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.333333 LAYER VIA3 ;
  END BIAS_TC_POT[2]
  PIN BIAS_TC_POT[1] 
    ANTENNAPARTIALMETALAREA 0.3065 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.418 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8832 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.482 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1648 LAYER M4 ;
  END BIAS_TC_POT[1]
  PIN BIAS_TC_POT[0] 
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.982 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.7648 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.8734 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 189.72 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3 ;
  END BIAS_TC_POT[0]
  PIN BIAS_LC_POT[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5498 LAYER M2 ;
  END BIAS_LC_POT[5]
  PIN BIAS_LC_POT[4] 
    ANTENNAPARTIALMETALAREA 0.127 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5588 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.225 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.434 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.086 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8224 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ; 
    ANTENNAMAXAREACAR 58.5451 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 257.874 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.63934 LAYER VIA4 ;
  END BIAS_LC_POT[4]
  PIN BIAS_LC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.091 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.442 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.838 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7312 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M5 ; 
    ANTENNAMAXAREACAR 39.05 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 174.937 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA5 ;
  END BIAS_LC_POT[3]
  PIN BIAS_LC_POT[2] 
    ANTENNAPARTIALMETALAREA 0.191 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8404 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.902 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 69.65 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 309.577 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3 ;
  END BIAS_LC_POT[2]
  PIN BIAS_LC_POT[1] 
    ANTENNAPARTIALMETALAREA 0.4535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9954 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.8604 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 132.142 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.647249 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.642 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2688 LAYER M4 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 56.43 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 249.761 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.647249 LAYER VIA4 ;
  END BIAS_LC_POT[1]
  PIN BIAS_LC_POT[0] 
    ANTENNAPARTIALMETALAREA 1.066 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6904 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.344 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.4016 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.9329 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 166.947 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_LC_POT[0]
  PIN BIAS_TIA_G_POT[16] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.261 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1484 LAYER M2 ;
  END BIAS_TIA_G_POT[16]
  PIN BIAS_TIA_G_POT[15] 
    ANTENNAPARTIALMETALAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0164 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.878 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9072 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.122 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.5808 LAYER M5 ;
  END BIAS_TIA_G_POT[15]
  PIN BIAS_TIA_G_POT[14] 
    ANTENNAPARTIALMETALAREA 0.306 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.902 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.2128 LAYER M3 ;
  END BIAS_TIA_G_POT[14]
  PIN BIAS_TIA_G_POT[13] 
    ANTENNAPARTIALMETALAREA 0.3125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.375 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.398 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.3952 LAYER M3 ;
  END BIAS_TIA_G_POT[13]
  PIN BIAS_TIA_G_POT[12] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 4.962 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.8768 LAYER M5 ;
  END BIAS_TIA_G_POT[12]
  PIN BIAS_TIA_G_POT[11] 
    ANTENNAPARTIALMETALAREA 0.3545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5598 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.142 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.886 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1424 LAYER M5 ;
  END BIAS_TIA_G_POT[11]
  PIN BIAS_TIA_G_POT[10] 
    ANTENNAPARTIALMETALAREA 0.389 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7116 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.022 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.7408 LAYER M3 ;
  END BIAS_TIA_G_POT[10]
  PIN BIAS_TIA_G_POT[9] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.0705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7102 LAYER M2 ;
  END BIAS_TIA_G_POT[9]
  PIN BIAS_TIA_G_POT[8] 
    ANTENNAPARTIALMETALAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0164 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.7 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 25.168 LAYER M5 ;
  END BIAS_TIA_G_POT[8]
  PIN BIAS_TIA_G_POT[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.8125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.975 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2704 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.238 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 31.8912 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 16.502 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 72.6528 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.476 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5824 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 2.668 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 11.8272 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M7 ; 
    ANTENNAMAXAREACAR 212.107 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 933.543 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.66667 LAYER VIA7 ;
  END BIAS_TIA_G_POT[7]
  PIN BIAS_TIA_G_POT[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.189 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2756 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.484 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.858 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8192 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 29.918 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 131.683 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.186 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M6 ; 
    ANTENNAMAXAREACAR 97.3048 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 431.874 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.267 LAYER VIA6 ;
  END BIAS_TIA_G_POT[6]
  PIN BIAS_TIA_G_POT[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4134 LAYER M2 ;
  END BIAS_TIA_G_POT[5]
  PIN BIAS_TIA_G_POT[4] 
    ANTENNAPARTIALMETALAREA 0.378 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6632 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.582 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6048 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ; 
    ANTENNAMAXAREACAR 43.5827 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 195.005 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.0929 LAYER VIA4 ;
  END BIAS_TIA_G_POT[4]
  PIN BIAS_TIA_G_POT[3] 
    ANTENNAPARTIALMETALAREA 1.3745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0478 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2 ; 
    ANTENNAMAXAREACAR 20.4563 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 89.8153 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.158 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7392 LAYER M3 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.7363 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 100.482 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3 ;
  END BIAS_TIA_G_POT[3]
  PIN BIAS_TIA_G_POT[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.251 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1924 LAYER M2 ;
  END BIAS_TIA_G_POT[2]
  PIN BIAS_TIA_G_POT[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.8165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6366 LAYER M2 ;
  END BIAS_TIA_G_POT[1]
  PIN BIAS_TIA_G_POT[0] 
    ANTENNAPARTIALMETALAREA 0.257 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1308 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.186 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.862 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8368 LAYER M4 ;
  END BIAS_TIA_G_POT[0]
  PIN BIAS_REV_POT[13] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0816 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.818 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6432 LAYER M4 ;
  END BIAS_REV_POT[13]
  PIN BIAS_REV_POT[12] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.538 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8112 LAYER M4 ;
  END BIAS_REV_POT[12]
  PIN BIAS_REV_POT[11] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
  END BIAS_REV_POT[11]
  PIN BIAS_REV_POT[10] 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9632 LAYER M4 ;
  END BIAS_REV_POT[10]
  PIN BIAS_REV_POT[9] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.558 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6552 LAYER M2 ;
  END BIAS_REV_POT[9]
  PIN BIAS_REV_POT[8] 
    ANTENNAPARTIALMETALAREA 0.0725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.319 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
  END BIAS_REV_POT[8]
  PIN BIAS_REV_POT[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.084 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3696 LAYER M2 ;
  END BIAS_REV_POT[7]
  PIN BIAS_REV_POT[6] 
    ANTENNAPARTIALMETALAREA 0.0215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0946 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.062 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7168 LAYER M3 ;
  END BIAS_REV_POT[6]
  PIN BIAS_REV_POT[5] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
  END BIAS_REV_POT[5]
  PIN BIAS_REV_POT[4] 
    ANTENNAPARTIALMETALAREA 0.0705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3102 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.982 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3648 LAYER M3 ;
  END BIAS_REV_POT[4]
  PIN BIAS_REV_POT[3] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.146 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M3 ;
  END BIAS_REV_POT[3]
  PIN BIAS_REV_POT[2] 
    ANTENNAPARTIALMETALAREA 0.1425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.627 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.646 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8864 LAYER M3 ;
  END BIAS_REV_POT[2]
  PIN BIAS_REV_POT[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.063 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3212 LAYER M2 ;
  END BIAS_REV_POT[1]
  PIN BIAS_REV_POT[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4158 LAYER M2 ;
  END BIAS_REV_POT[0]
  PIN BIAS_TC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.9595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2218 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.042 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.6097 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 199.57 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_TC_DSADC[5]
  PIN BIAS_TC_DSADC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.349 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9796 LAYER M2 ;
  END BIAS_TC_DSADC[4]
  PIN BIAS_TC_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.5695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5058 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.562 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.446 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_TC_DSADC[3]
  PIN BIAS_TC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 1.015 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.466 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.854 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8016 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.4163 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 80.8485 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_TC_DSADC[2]
  PIN BIAS_TC_DSADC[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.8955 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9842 LAYER M2 ;
  END BIAS_TC_DSADC[1]
  PIN BIAS_TC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.086 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3784 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.418 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2832 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 45.2056 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 198.947 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA4 ;
  END BIAS_TC_DSADC[0]
  PIN BIAS_LC_DSADC[5] 
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.2135 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9834 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.97 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.712 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 120.434 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 529.405 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA4 ;
  END BIAS_LC_DSADC[5]
  PIN BIAS_LC_DSADC[4] 
    ANTENNAPARTIALMETALAREA 1.357 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9708 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.854 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.418 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8832 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 62.0477 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 272.712 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA4 ;
  END BIAS_LC_DSADC[4]
  PIN BIAS_LC_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.377 LAYER M2 ;
  END BIAS_LC_DSADC[3]
  PIN BIAS_LC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 1.226 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3944 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3568 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.4786 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 139.262 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3 ;
  END BIAS_LC_DSADC[2]
  PIN BIAS_LC_DSADC[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.0955 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8642 LAYER M2 ;
  END BIAS_LC_DSADC[1]
  PIN BIAS_LC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.131 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5764 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.902 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0128 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.518 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3232 LAYER M4 ;
  END BIAS_LC_DSADC[0]
  PIN BIAS_RIN_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.191 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8404 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.246 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.778 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4672 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M5 ; 
    ANTENNAMAXAREACAR 125.466 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 555.262 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.589 LAYER VIA5 ;
  END BIAS_RIN_DSADC[5]
  PIN BIAS_RIN_DSADC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.147 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0468 LAYER M2 ;
  END BIAS_RIN_DSADC[4]
  PIN BIAS_RIN_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.4215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8546 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.898 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.9806 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 75.7087 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.809061 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.262 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5968 LAYER M4 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 37.4013 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 166.272 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.809061 LAYER VIA4 ;
  END BIAS_RIN_DSADC[3]
  PIN BIAS_RIN_DSADC[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.874 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8896 LAYER M2 ;
  END BIAS_RIN_DSADC[2]
  PIN BIAS_RIN_DSADC[1] 
    ANTENNAPARTIALMETALAREA 1.2265 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3966 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.864 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2896 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 74.5922 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 330.848 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3 ;
  END BIAS_RIN_DSADC[1]
  PIN BIAS_RIN_DSADC[0] 
    ANTENNAPARTIALMETALAREA 1.953 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5932 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.224 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.8736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 68.4693 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 302.971 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3 ;
  END BIAS_RIN_DSADC[0]
  PIN BIAS_RFB_DSADC[5] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6045 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7038 LAYER M2 ;
  END BIAS_RFB_DSADC[5]
  PIN BIAS_RFB_DSADC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.256 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6584 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.686 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4624 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.422 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9008 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 10.93 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 48.18 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.104 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5016 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 5.1 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 22.528 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 176.876 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 776.417 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA7 ;
  END BIAS_RFB_DSADC[4]
  PIN BIAS_RFB_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.742 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3088 LAYER M2 ;
  END BIAS_RFB_DSADC[3]
  PIN BIAS_RFB_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.131 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5764 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.542 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8288 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 LAYER M4 ; 
    ANTENNAMAXAREACAR 74.245 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 327.362 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.854701 LAYER VIA4 ;
  END BIAS_RFB_DSADC[2]
  PIN BIAS_RFB_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.1345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5918 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.822 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6608 LAYER M4 ;
  END BIAS_RFB_DSADC[1]
  PIN BIAS_RFB_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.278 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.938 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1712 LAYER M3 ;
  END BIAS_RFB_DSADC[0]
  PIN BIAS_DSADC_VCM[13] 
    ANTENNAPARTIALMETALAREA 4.315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.03 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.226 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M3 ;
  END BIAS_DSADC_VCM[13]
  PIN BIAS_DSADC_VCM[12] 
    ANTENNAPARTIALMETALAREA 0.1715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7546 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.572 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6048 LAYER M3 ;
  END BIAS_DSADC_VCM[12]
  PIN BIAS_DSADC_VCM[11] 
    ANTENNAPARTIALMETALAREA 0.069 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3 ;
  END BIAS_DSADC_VCM[11]
  PIN BIAS_DSADC_VCM[10] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0684 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.838 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7312 LAYER M4 ;
  END BIAS_DSADC_VCM[10]
  PIN BIAS_DSADC_VCM[9] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.468 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1472 LAYER M3 ;
  END BIAS_DSADC_VCM[9]
  PIN BIAS_DSADC_VCM[8] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3014 LAYER M2 ;
  END BIAS_DSADC_VCM[8]
  PIN BIAS_DSADC_VCM[7] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.698 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1152 LAYER M4 ;
  END BIAS_DSADC_VCM[7]
  PIN BIAS_DSADC_VCM[6] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.692 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
  END BIAS_DSADC_VCM[6]
  PIN BIAS_DSADC_VCM[5] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.298 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3552 LAYER M4 ;
  END BIAS_DSADC_VCM[5]
  PIN BIAS_DSADC_VCM[4] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.692 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3 ;
  END BIAS_DSADC_VCM[4]
  PIN BIAS_DSADC_VCM[3] 
    ANTENNAPARTIALMETALAREA 0.169 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7436 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.746 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3264 LAYER M3 ;
  END BIAS_DSADC_VCM[3]
  PIN BIAS_DSADC_VCM[2] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.882 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9248 LAYER M3 ;
  END BIAS_DSADC_VCM[2]
  PIN BIAS_DSADC_VCM[1] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8048 LAYER M3 ;
  END BIAS_DSADC_VCM[1]
  PIN BIAS_DSADC_VCM[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0275 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.165 LAYER M2 ;
  END BIAS_DSADC_VCM[0]
  PIN dsadc_conv_done 
    ANTENNAPARTIALMETALAREA 0.422 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8568 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.398 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7952 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 11.862 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 52.2368 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M5 ; 
    ANTENNAMAXAREACAR 585.895 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2584.6 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.58303 LAYER VIA5 ;
  END dsadc_conv_done
  PIN dsadc_en 
    ANTENNAPARTIALMETALAREA 0.072 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3168 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.43 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 24.024 LAYER M5 ;
  END dsadc_en
  PIN dsadc_clk 
    ANTENNAPARTIALMETALAREA 0.196 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2156 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 32.962 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.4342 LAYER M3 ;
  END dsadc_clk
  PIN dsadc_switch[2] 
    ANTENNAPARTIALMETALAREA 0.4695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0658 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6928 LAYER M3 ;
  END dsadc_switch[2]
  PIN dsadc_switch[1] 
    ANTENNAPARTIALMETALAREA 0.167 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7348 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.763 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4012 LAYER M3 ;
  END dsadc_switch[1]
  PIN dsadc_switch[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.251 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1044 LAYER M2 ;
  END dsadc_switch[0]
  PIN dac_en_pot 
    ANTENNAPARTIALMETALAREA 0.1265 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5566 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.722 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.582 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6048 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.378 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 14.9072 LAYER M5 ;
  END dac_en_pot
  PIN adc_ext_in 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.337 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5268 LAYER M2 ;
  END adc_ext_in
  PIN atp_en 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5905 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6422 LAYER M2 ;
  END atp_en
  PIN atp_sel 
    ANTENNAPARTIALMETALAREA 0.135 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.594 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.206 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.1504 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.982 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.1648 LAYER M5 ;
  END atp_sel
  PIN adc_sel 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8722 LAYER M2 ;
  END adc_sel
  PIN saradc_clk 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 72.784 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.5904 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.64 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.28 LAYER M4 ;
  END saradc_clk
  PIN saradc_rdy 
    ANTENNAPARTIALMETALAREA 1.3025 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.731 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.978 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.5472 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.086 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4224 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 8.698 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 38.3152 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 2.762 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 12.1968 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0269 LAYER M7 ; 
    ANTENNAMAXAREACAR 195.442 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 854 LAYER M7 ;
    ANTENNAMAXCUTCAR 4.46097 LAYER VIA7 ;
  END saradc_rdy
  PIN saradc_rst 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1242 LAYER M2 ;
  END saradc_rst
  PIN saradc_data[9] 
    ANTENNAPARTIALMETALAREA 0.3315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4586 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.298 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3552 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.112 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9808 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 12.598 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 55.4752 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.246 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6 ; 
    ANTENNAMAXAREACAR 158.027 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 698.988 LAYER M6 ;
    ANTENNAMAXCUTCAR 4.08163 LAYER VIA6 ;
  END saradc_data[9]
  PIN saradc_data[8] 
    ANTENNAPARTIALMETALAREA 0.351 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0935 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4554 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.442 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.678 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4272 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.664 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0096 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6 ; 
    ANTENNAMAXAREACAR 75.4959 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 338.498 LAYER M6 ;
    ANTENNAMAXCUTCAR 4.08163 LAYER VIA6 ;
  END saradc_data[8]
  PIN saradc_data[7] 
    ANTENNAPARTIALMETALAREA 1.2325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.467 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 16.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 72.1248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M3 ; 
    ANTENNAMAXAREACAR 713.21 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3138.14 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.63265 LAYER VIA3 ;
  END saradc_data[7]
  PIN saradc_data[6] 
    ANTENNAPARTIALMETALAREA 0.207 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9108 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.208 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.8032 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M4 ; 
    ANTENNAMAXAREACAR 133.455 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 591.396 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.44898 LAYER VIA4 ;
  END saradc_data[6]
  PIN saradc_data[5] 
    ANTENNAPARTIALMETALAREA 0.351 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.5735 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5674 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.446 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0064 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 15.978 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 70.3472 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.722 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2208 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6 ; 
    ANTENNAMAXAREACAR 47.7306 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 203.29 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.67347 LAYER VIA6 ;
  END saradc_data[5]
  PIN saradc_data[4] 
    ANTENNAPARTIALMETALAREA 0.5715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5146 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.706 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1504 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 13.344 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 58.8016 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 583.822 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2572.75 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.85714 LAYER VIA5 ;
  END saradc_data[4]
  PIN saradc_data[3] 
    ANTENNAPARTIALMETALAREA 0.451 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9844 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.2135 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3834 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.938 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1712 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 5.768 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 25.4672 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M7 ; 
    ANTENNAMAXAREACAR 430.68 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 1903.43 LAYER M7 ;
    ANTENNAMAXCUTCAR 4.89796 LAYER VIA7 ;
  END saradc_data[3]
  PIN saradc_data[2] 
    ANTENNAPARTIALMETALAREA 0.5715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5146 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.518 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3232 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.406 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8304 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M4 ; 
    ANTENNAMAXAREACAR 401.827 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1757.14 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.72911 LAYER VIA4 ;
  END saradc_data[2]
  PIN saradc_data[1] 
    ANTENNAPARTIALMETALAREA 0.7665 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3726 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 15.042 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.2288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.378 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7072 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.666 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9744 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 63.3061 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 284.106 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.85714 LAYER VIA5 ;
  END saradc_data[1]
  PIN saradc_data[0] 
    ANTENNAPARTIALMETALAREA 0.9435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1514 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 16.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.8608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.482 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1648 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M4 ; 
    ANTENNAMAXAREACAR 37.7551 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 169.886 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.04082 LAYER VIA4 ;
  END saradc_data[0]
END MCU

END LIBRARY
