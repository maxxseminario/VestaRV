##
## LEF for PtnCells ;
## created by Innovus v20.12-s088_1 on Mon Nov 17 15:45:30 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO MCU
  CLASS BLOCK ;
  SIZE 1186.000000 BY 686.000000 ;
  FOREIGN MCU 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN resetn_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.442 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 25.842 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 113.749 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6  ;
    ANTENNAMAXAREACAR 974.013 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 4292.32 LAYER M6  ;
    ANTENNAMAXCUTCAR 3.32103 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 131.365000 0.000000 131.465000 0.520000 ;
    END
  END resetn_in
  PIN resetn_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.325 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.474 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 111.130000 0.000000 111.230000 0.520000 ;
    END
  END resetn_out
  PIN resetn_dir
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.6365 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8446 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 121.725000 0.000000 121.825000 0.520000 ;
    END
  END resetn_dir
  PIN resetn_ren
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.5895 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6378 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 125.685000 0.000000 125.785000 0.520000 ;
    END
  END resetn_ren
  PIN prt1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.4155 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.9162 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2  ;
    ANTENNAMAXAREACAR 570.452 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 2511.78 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.369004 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 45.565000 1186.000000 45.665000 ;
    END
  END prt1_in[7]
  PIN prt1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.6125 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 99.495 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 10.962 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.2768 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3  ;
    ANTENNAMAXAREACAR 112.492 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 485.767 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.08401 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 133.565000 1186.000000 133.665000 ;
    END
  END prt1_in[6]
  PIN prt1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0905 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.0422 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 11.706 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.5504 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1305 LAYER M3  ;
    ANTENNAMAXAREACAR 98.311 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 432.269 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAMAXCUTCAR 0.782188 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M4  ;
    ANTENNAGATEAREA 0.2577 LAYER M4  ;
    ANTENNAMAXAREACAR 99.1725 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 436.23 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.782188 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 221.565000 1186.000000 221.665000 ;
    END
  END prt1_in[5]
  PIN prt1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8725 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.439 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 11.59 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.04 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1305 LAYER M3  ;
    ANTENNAMAXAREACAR 97.1232 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 427.042 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAMAXCUTCAR 0.782188 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.178 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M4  ;
    ANTENNAGATEAREA 0.1305 LAYER M4  ;
    ANTENNAMAXAREACAR 98.4872 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 433.381 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAMAXCUTCAR 0.935444 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 6.006 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 26.4704 LAYER M5  ;
    ANTENNAGATEAREA 0.2577 LAYER M5  ;
    ANTENNAMAXAREACAR 121.793 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 536.099 LAYER M5  ;
    ANTENNAMAXCUTCAR 0.935444 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 309.565000 1186.000000 309.665000 ;
    END
  END prt1_in[4]
  PIN prt1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.176 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1936 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4982 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 4.242 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8422 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 LAYER M4  ;
    ANTENNAMAXAREACAR 19.556 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 25.0566 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAMAXCUTCAR 0.314465 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.52 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER M5  ;
    ANTENNAGATEAREA 0.318 LAYER M5  ;
    ANTENNAMAXAREACAR 30.6252 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 45.1069 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.25786 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 397.565000 1186.000000 397.665000 ;
    END
  END prt1_in[3]
  PIN prt1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1135 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3434 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 12.418 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.7712 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1931 LAYER M3  ;
    ANTENNAMAXAREACAR 122.456 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 540.411 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 485.565000 1186.000000 485.665000 ;
    END
  END prt1_in[2]
  PIN prt1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1575 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.937 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 9.782 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.0848 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3  ;
    ANTENNAMAXAREACAR 112.431 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 494.435 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 573.565000 1186.000000 573.665000 ;
    END
  END prt1_in[1]
  PIN prt1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.0995 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 97.2378 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 4.418 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4832 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3  ;
    ANTENNAMAXAREACAR 52.3228 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 229.855 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 661.565000 1186.000000 661.665000 ;
    END
  END prt1_in[0]
  PIN prt1_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 25.330000 1186.000000 25.430000 ;
    END
  END prt1_out[7]
  PIN prt1_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 12.499 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.0836 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 113.330000 1186.000000 113.430000 ;
    END
  END prt1_out[6]
  PIN prt1_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 201.330000 1186.000000 201.430000 ;
    END
  END prt1_out[5]
  PIN prt1_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 289.330000 1186.000000 289.430000 ;
    END
  END prt1_out[4]
  PIN prt1_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.796 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9024 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 8.186 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.0624 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 377.330000 1186.000000 377.430000 ;
    END
  END prt1_out[3]
  PIN prt1_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.092 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 8.804 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.8256 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 465.330000 1186.000000 465.430000 ;
    END
  END prt1_out[2]
  PIN prt1_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 14.535 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.042 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 553.330000 1186.000000 553.430000 ;
    END
  END prt1_out[1]
  PIN prt1_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 11.575 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.018 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 641.330000 1186.000000 641.430000 ;
    END
  END prt1_out[0]
  PIN prt1_dir[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0115 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2506 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 8.782 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.6848 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 35.925000 1186.000000 36.025000 ;
    END
  END prt1_dir[7]
  PIN prt1_dir[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2165 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9526 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.266 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2144 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 123.925000 1186.000000 124.025000 ;
    END
  END prt1_dir[6]
  PIN prt1_dir[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 211.925000 1186.000000 212.025000 ;
    END
  END prt1_dir[5]
  PIN prt1_dir[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8214 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 9.098 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.0752 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 299.925000 1186.000000 300.025000 ;
    END
  END prt1_dir[4]
  PIN prt1_dir[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 7.064 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.1696 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 387.925000 1186.000000 388.025000 ;
    END
  END prt1_dir[3]
  PIN prt1_dir[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0855 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4202 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 475.925000 1186.000000 476.025000 ;
    END
  END prt1_dir[2]
  PIN prt1_dir[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 563.925000 1186.000000 564.025000 ;
    END
  END prt1_dir[1]
  PIN prt1_dir[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 12.2345 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.9198 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 651.925000 1186.000000 652.025000 ;
    END
  END prt1_dir[0]
  PIN prt1_ren[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0855 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4202 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 39.885000 1186.000000 39.985000 ;
    END
  END prt1_ren[7]
  PIN prt1_ren[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1805 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1942 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.466 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4944 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 127.885000 1186.000000 127.985000 ;
    END
  END prt1_ren[6]
  PIN prt1_ren[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 215.885000 1186.000000 215.985000 ;
    END
  END prt1_ren[5]
  PIN prt1_ren[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2985 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5574 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 9.362 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.2368 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 303.885000 1186.000000 303.985000 ;
    END
  END prt1_ren[4]
  PIN prt1_ren[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2475 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.089 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 3.566 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.7344 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 391.885000 1186.000000 391.985000 ;
    END
  END prt1_ren[3]
  PIN prt1_ren[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5295 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7738 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.702 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5328 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 479.885000 1186.000000 479.985000 ;
    END
  END prt1_ren[2]
  PIN prt1_ren[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 567.885000 1186.000000 567.985000 ;
    END
  END prt1_ren[1]
  PIN prt1_ren[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 12.3905 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.6062 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 655.885000 1186.000000 655.985000 ;
    END
  END prt1_ren[0]
  PIN prt2_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7785 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5134 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0595 LAYER M2  ;
    ANTENNAMAXAREACAR 18.0714 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 78.4706 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.336134 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 302.965000 0.000000 303.065000 0.520000 ;
    END
  END prt2_in[7]
  PIN prt2_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4122 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2  ;
    ANTENNAMAXAREACAR 27.7954 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 121.522 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 388.765000 0.000000 388.865000 0.520000 ;
    END
  END prt2_in[6]
  PIN prt2_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7125 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.135 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 LAYER M2  ;
    ANTENNAMAXAREACAR 7.72407 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 32.9611 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.185185 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 474.565000 0.000000 474.665000 0.520000 ;
    END
  END prt2_in[5]
  PIN prt2_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 4.362 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2368 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3  ;
    ANTENNAMAXAREACAR 146.784 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 630.772 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 560.365000 0.000000 560.465000 0.520000 ;
    END
  END prt2_in[4]
  PIN prt2_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.234 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5334 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M2  ;
    ANTENNAMAXAREACAR 6.88784 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 9.43291 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.104822 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 646.165000 0.000000 646.265000 0.520000 ;
    END
  END prt2_in[3]
  PIN prt2_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6785 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9854 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0893 LAYER M2  ;
    ANTENNAMAXAREACAR 11.5812 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 48.6697 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.223964 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 731.965000 0.000000 732.065000 0.520000 ;
    END
  END prt2_in[2]
  PIN prt2_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7155 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1482 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0893 LAYER M2  ;
    ANTENNAMAXAREACAR 11.3908 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 48.0739 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.223964 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 817.765000 0.000000 817.865000 0.520000 ;
    END
  END prt2_in[1]
  PIN prt2_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 30.982 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.365 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0381 LAYER M3  ;
    ANTENNAMAXAREACAR 850.332 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 3731.77 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.04987 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 903.565000 0.000000 903.665000 0.520000 ;
    END
  END prt2_in[0]
  PIN prt2_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.471 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0724 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 9.862 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.4368 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 282.730000 0.000000 282.830000 0.520000 ;
    END
  END prt2_out[7]
  PIN prt2_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.681 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 368.530000 0.000000 368.630000 0.520000 ;
    END
  END prt2_out[6]
  PIN prt2_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.577 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6708 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 454.330000 0.000000 454.430000 0.520000 ;
    END
  END prt2_out[5]
  PIN prt2_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.679 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9876 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 10.038 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.2112 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 540.130000 0.000000 540.230000 0.520000 ;
    END
  END prt2_out[4]
  PIN prt2_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 625.930000 0.000000 626.030000 0.520000 ;
    END
  END prt2_out[3]
  PIN prt2_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.152 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 13.586 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.8224 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 711.730000 0.000000 711.830000 0.520000 ;
    END
  END prt2_out[2]
  PIN prt2_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.279 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2276 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 797.530000 0.000000 797.630000 0.520000 ;
    END
  END prt2_out[1]
  PIN prt2_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.512 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 883.330000 0.000000 883.430000 0.520000 ;
    END
  END prt2_out[0]
  PIN prt2_dir[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.711 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1284 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 8.602 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.8928 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 293.325000 0.000000 293.425000 0.520000 ;
    END
  END prt2_dir[7]
  PIN prt2_dir[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.5835 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6554 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 379.125000 0.000000 379.225000 0.520000 ;
    END
  END prt2_dir[6]
  PIN prt2_dir[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.6815 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0426 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 464.925000 0.000000 465.025000 0.520000 ;
    END
  END prt2_dir[5]
  PIN prt2_dir[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.2715 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1946 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 550.725000 0.000000 550.825000 0.520000 ;
    END
  END prt2_dir[4]
  PIN prt2_dir[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.2715 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1946 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 636.525000 0.000000 636.625000 0.520000 ;
    END
  END prt2_dir[3]
  PIN prt2_dir[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.531 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3364 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.362 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.2368 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 722.325000 0.000000 722.425000 0.520000 ;
    END
  END prt2_dir[2]
  PIN prt2_dir[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.6595 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9018 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 808.125000 0.000000 808.225000 0.520000 ;
    END
  END prt2_dir[1]
  PIN prt2_dir[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.2785 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2254 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 893.925000 0.000000 894.025000 0.520000 ;
    END
  END prt2_dir[0]
  PIN prt2_ren[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6435 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8314 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 8.878 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.1072 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 297.285000 0.000000 297.385000 0.520000 ;
    END
  END prt2_ren[7]
  PIN prt2_ren[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.7235 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2714 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 383.085000 0.000000 383.185000 0.520000 ;
    END
  END prt2_ren[6]
  PIN prt2_ren[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7345 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2318 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.758 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7792 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 468.885000 0.000000 468.985000 0.520000 ;
    END
  END prt2_ren[5]
  PIN prt2_ren[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.5625 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.519 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 554.685000 0.000000 554.785000 0.520000 ;
    END
  END prt2_ren[4]
  PIN prt2_ren[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8875 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.905 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 3.146 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8864 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 640.485000 0.000000 640.585000 0.520000 ;
    END
  END prt2_ren[3]
  PIN prt2_ren[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.667 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9348 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.2095 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7658 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 726.285000 0.000000 726.385000 0.520000 ;
    END
  END prt2_ren[2]
  PIN prt2_ren[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.2855 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3002 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 812.085000 0.000000 812.185000 0.520000 ;
    END
  END prt2_ren[1]
  PIN prt2_ren[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.6855 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0602 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 897.885000 0.000000 897.985000 0.520000 ;
    END
  END prt2_ren[0]
  PIN prt3_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.7995 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.8058 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2  ;
    ANTENNAMAXAREACAR 698.801 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 3074.69 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.738007 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 641.335000 0.520000 641.435000 ;
    END
  END prt3_in[7]
  PIN prt3_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.9905 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.4022 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 16.178 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.2272 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 610.052 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 2670.41 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 553.335000 0.520000 553.435000 ;
    END
  END prt3_in[6]
  PIN prt3_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9325 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.903 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 15.938 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.1712 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 2.258 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9792 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4  ;
    ANTENNAMAXAREACAR 39.3685 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 175.57 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 465.335000 0.520000 465.435000 ;
    END
  END prt3_in[5]
  PIN prt3_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6325 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.783 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 13.382 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.9248 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.278 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.622 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9808 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M5  ;
    ANTENNAMAXAREACAR 47.4781 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 209.971 LAYER M5  ;
    ANTENNAMAXCUTCAR 0.876988 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 377.335000 0.520000 377.435000 ;
    END
  END prt3_in[4]
  PIN prt3_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7355 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8362 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 18.226 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.2384 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1707 LAYER M3  ;
    ANTENNAMAXAREACAR 119.268 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 524.402 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 289.335000 0.520000 289.435000 ;
    END
  END prt3_in[3]
  PIN prt3_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5755 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5322 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 16.952 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.7648 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 644.59 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 2824.86 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 201.335000 0.520000 201.435000 ;
    END
  END prt3_in[2]
  PIN prt3_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.5355 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.9562 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 4.722 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8208 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 285.009 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1255.83 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 113.335000 0.520000 113.435000 ;
    END
  END prt3_in[1]
  PIN prt3_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9105 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4502 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 9.438 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.5712 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3  ;
    ANTENNAMAXAREACAR 294.622 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1280.64 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 25.335000 0.520000 25.435000 ;
    END
  END prt3_in[0]
  PIN prt3_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 14.743 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.9572 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 661.570000 0.520000 661.670000 ;
    END
  END prt3_out[7]
  PIN prt3_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 6.423 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.3492 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 573.570000 0.520000 573.670000 ;
    END
  END prt3_out[6]
  PIN prt3_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.036 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5584 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.766 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8144 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 485.570000 0.520000 485.670000 ;
    END
  END prt3_out[5]
  PIN prt3_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.379 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1556 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 397.570000 0.520000 397.670000 ;
    END
  END prt3_out[4]
  PIN prt3_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.792 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8848 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.806 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9904 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 309.570000 0.520000 309.670000 ;
    END
  END prt3_out[3]
  PIN prt3_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.175 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.458 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 221.570000 0.520000 221.670000 ;
    END
  END prt3_out[2]
  PIN prt3_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 12.855 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.65 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 133.570000 0.520000 133.670000 ;
    END
  END prt3_out[1]
  PIN prt3_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.901 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2084 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 45.570000 0.520000 45.670000 ;
    END
  END prt3_out[0]
  PIN prt3_dir[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 14.2415 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.7066 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 650.975000 0.520000 651.075000 ;
    END
  END prt3_dir[7]
  PIN prt3_dir[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 5.0055 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1562 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 562.975000 0.520000 563.075000 ;
    END
  END prt3_dir[6]
  PIN prt3_dir[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.186 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 474.975000 0.520000 475.075000 ;
    END
  END prt3_dir[5]
  PIN prt3_dir[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4165 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8326 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.842 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.3488 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 386.975000 0.520000 387.075000 ;
    END
  END prt3_dir[4]
  PIN prt3_dir[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1515 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6666 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.646 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.4864 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 298.975000 0.520000 299.075000 ;
    END
  END prt3_dir[3]
  PIN prt3_dir[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 13.7345 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.5198 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 210.975000 0.520000 211.075000 ;
    END
  END prt3_dir[2]
  PIN prt3_dir[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0495 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.8618 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.646 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8864 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 122.975000 0.520000 123.075000 ;
    END
  END prt3_dir[1]
  PIN prt3_dir[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.1345 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8798 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 34.975000 0.520000 35.075000 ;
    END
  END prt3_dir[0]
  PIN prt3_ren[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 13.3255 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.7642 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 647.015000 0.520000 647.115000 ;
    END
  END prt3_ren[7]
  PIN prt3_ren[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 5.1075 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.561 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 559.015000 0.520000 559.115000 ;
    END
  END prt3_ren[6]
  PIN prt3_ren[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1462 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 471.015000 0.520000 471.115000 ;
    END
  END prt3_ren[5]
  PIN prt3_ren[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9062 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.77 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.032 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0582 LAYER M3  ;
    ANTENNAMAXAREACAR 258.459 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1136.85 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.687285 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 383.015000 0.520000 383.115000 ;
    END
  END prt3_ren[4]
  PIN prt3_ren[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 6.568 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.9872 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 295.015000 0.520000 295.115000 ;
    END
  END prt3_ren[3]
  PIN prt3_ren[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 9.6885 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.7614 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 207.015000 0.520000 207.115000 ;
    END
  END prt3_ren[2]
  PIN prt3_ren[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 14.3125 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.107 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 119.015000 0.520000 119.115000 ;
    END
  END prt3_ren[1]
  PIN prt3_ren[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5805 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5542 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.118 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 31.015000 0.520000 31.115000 ;
    END
  END prt3_ren[0]
  PIN prt4_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6042 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 26.828 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.131 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3  ;
    ANTENNAMAXAREACAR 389.192 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1708.37 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 646.165000 685.480000 646.265000 686.000000 ;
    END
  END prt4_in[7]
  PIN prt4_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1642 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 19.838 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.4192 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3  ;
    ANTENNAMAXAREACAR 198.371 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 873.831 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.08401 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 560.365000 685.480000 560.465000 686.000000 ;
    END
  END prt4_in[6]
  PIN prt4_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6785 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3854 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 9.504 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.9056 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3  ;
    ANTENNAMAXAREACAR 251.47 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1102.34 LAYER M3  ;
    ANTENNAMAXCUTCAR 2.16802 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 474.565000 685.480000 474.665000 686.000000 ;
    END
  END prt4_in[5]
  PIN prt4_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9755 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6922 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 4.858 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.4192 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1204 LAYER M4  ;
    ANTENNAMAXAREACAR 63.5979 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 279.093 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.25012 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 388.765000 685.480000 388.865000 686.000000 ;
    END
  END prt4_in[4]
  PIN prt4_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4505 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.4262 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.246 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5264 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1456 LAYER M3  ;
    ANTENNAMAXAREACAR 15.2257 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 66.8666 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.08401 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 302.965000 685.480000 303.065000 686.000000 ;
    END
  END prt4_in[3]
  PIN prt4_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 11.998 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.8352 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 6.818 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0432 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4  ;
    ANTENNAMAXAREACAR 96.3583 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 423.219 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.81869 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 217.165000 685.480000 217.265000 686.000000 ;
    END
  END prt4_in[2]
  PIN prt4_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.731 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 20.818 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.6432 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 6.556 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.9344 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0636 LAYER M4  ;
    ANTENNAMAXAREACAR 126.222 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 557.921 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAMAXCUTCAR 1.41509 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.506 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2704 LAYER M5  ;
    ANTENNAGATEAREA 0.1305 LAYER M5  ;
    ANTENNAMAXAREACAR 130.099 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 575.319 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.41509 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 131.365000 685.480000 131.465000 686.000000 ;
    END
  END prt4_in[1]
  PIN prt4_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2725 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 27.886 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.742 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 1080.52 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 4736.44 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 45.565000 685.480000 45.665000 686.000000 ;
    END
  END prt4_in[0]
  PIN prt4_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.292 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8806 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 82.8 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.256 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 625.930000 685.480000 626.030000 686.000000 ;
    END
  END prt4_out[7]
  PIN prt4_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.332 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4246 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 9.6 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.736 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 540.130000 685.480000 540.230000 686.000000 ;
    END
  END prt4_out[6]
  PIN prt4_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.43 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.473 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 19.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 22 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 454.330000 685.480000 454.430000 686.000000 ;
    END
  END prt4_out[5]
  PIN prt4_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 7.922 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8902 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 368.530000 685.480000 368.630000 686.000000 ;
    END
  END prt4_out[4]
  PIN prt4_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.968 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 5.998 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.4352 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 282.730000 685.480000 282.830000 686.000000 ;
    END
  END prt4_out[3]
  PIN prt4_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4564 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.278 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.8672 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 196.930000 685.480000 197.030000 686.000000 ;
    END
  END prt4_out[2]
  PIN prt4_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.922 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 74.5008 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 111.130000 685.480000 111.230000 686.000000 ;
    END
  END prt4_out[1]
  PIN prt4_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 25.330000 685.480000 25.430000 686.000000 ;
    END
  END prt4_out[0]
  PIN prt4_dir[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2915 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 11.506 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.6704 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 636.525000 685.480000 636.625000 686.000000 ;
    END
  END prt4_dir[7]
  PIN prt4_dir[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 2.3785 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5534 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 550.725000 685.480000 550.825000 686.000000 ;
    END
  END prt4_dir[6]
  PIN prt4_dir[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.968 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 2.5785 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4334 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 464.925000 685.480000 465.025000 686.000000 ;
    END
  END prt4_dir[5]
  PIN prt4_dir[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.968 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.6385 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0974 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 379.125000 685.480000 379.225000 686.000000 ;
    END
  END prt4_dir[4]
  PIN prt4_dir[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.871 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8324 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.968 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 5.242 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.1088 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 293.325000 685.480000 293.425000 686.000000 ;
    END
  END prt4_dir[3]
  PIN prt4_dir[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.511 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2484 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 13.278 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.4672 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 207.525000 685.480000 207.625000 686.000000 ;
    END
  END prt4_dir[2]
  PIN prt4_dir[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 17.122 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 75.3808 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 121.725000 685.480000 121.825000 686.000000 ;
    END
  END prt4_dir[1]
  PIN prt4_dir[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.386 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 72.1424 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 35.925000 685.480000 36.025000 686.000000 ;
    END
  END prt4_dir[0]
  PIN prt4_ren[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5075 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.233 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 13.502 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.4528 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 640.485000 685.480000 640.585000 686.000000 ;
    END
  END prt4_ren[7]
  PIN prt4_ren[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.9475 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.257 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 554.685000 685.480000 554.785000 686.000000 ;
    END
  END prt4_ren[6]
  PIN prt4_ren[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2105 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3262 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 7.066 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.1344 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 468.885000 685.480000 468.985000 686.000000 ;
    END
  END prt4_ren[5]
  PIN prt4_ren[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.7055 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5482 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 383.085000 685.480000 383.185000 686.000000 ;
    END
  END prt4_ren[4]
  PIN prt4_ren[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.1625 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.159 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 297.285000 685.480000 297.385000 686.000000 ;
    END
  END prt4_ren[3]
  PIN prt4_ren[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4435 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9514 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 13.202 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.1328 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 211.485000 685.480000 211.585000 686.000000 ;
    END
  END prt4_ren[2]
  PIN prt4_ren[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8035 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5354 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.342 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 71.9488 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 125.685000 685.480000 125.785000 686.000000 ;
    END
  END prt4_ren[1]
  PIN prt4_ren[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 17.146 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 75.4864 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 39.885000 685.480000 39.985000 686.000000 ;
    END
  END prt4_ren[0]
  PIN use_dac_glb_bias
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 614.515000 389.000000 614.615000 ;
    END
  END use_dac_glb_bias
  PIN en_bias_buf
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.246 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 613.970000 389.000000 614.070000 ;
    END
  END en_bias_buf
  PIN en_bias_gen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.041 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1804 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.566 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5344 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 6.096 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.9104 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 612.880000 389.000000 612.980000 ;
    END
  END en_bias_gen
  PIN BIAS_ADJ[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.358 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 609.610000 389.000000 609.710000 ;
    END
  END BIAS_ADJ[5]
  PIN BIAS_ADJ[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 2.438 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7712 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 610.155000 389.000000 610.255000 ;
    END
  END BIAS_ADJ[4]
  PIN BIAS_ADJ[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.019 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0836 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.178 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 610.700000 389.000000 610.800000 ;
    END
  END BIAS_ADJ[3]
  PIN BIAS_ADJ[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.344 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6016 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 611.245000 389.000000 611.345000 ;
    END
  END BIAS_ADJ[2]
  PIN BIAS_ADJ[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 611.790000 389.000000 611.890000 ;
    END
  END BIAS_ADJ[1]
  PIN BIAS_ADJ[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.278 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 612.335000 389.000000 612.435000 ;
    END
  END BIAS_ADJ[0]
  PIN BIAS_DBP[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.031 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1364 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.446 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0064 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.718 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2032 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 1.426 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3184 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 601.980000 389.000000 602.080000 ;
    END
  END BIAS_DBP[13]
  PIN BIAS_DBP[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 2.7985 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.4014 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 602.525000 389.000000 602.625000 ;
    END
  END BIAS_DBP[12]
  PIN BIAS_DBP[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 603.070000 389.000000 603.170000 ;
    END
  END BIAS_DBP[11]
  PIN BIAS_DBP[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1185 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5654 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.442 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3888 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2688 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 603.615000 389.000000 603.715000 ;
    END
  END BIAS_DBP[10]
  PIN BIAS_DBP[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 6.278 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6672 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 604.160000 389.000000 604.260000 ;
    END
  END BIAS_DBP[9]
  PIN BIAS_DBP[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.542 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8288 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 604.705000 389.000000 604.805000 ;
    END
  END BIAS_DBP[8]
  PIN BIAS_DBP[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 605.250000 389.000000 605.350000 ;
    END
  END BIAS_DBP[7]
  PIN BIAS_DBP[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0675 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.341 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 605.795000 389.000000 605.895000 ;
    END
  END BIAS_DBP[6]
  PIN BIAS_DBP[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.064 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3256 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 606.340000 389.000000 606.440000 ;
    END
  END BIAS_DBP[5]
  PIN BIAS_DBP[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.4255 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9162 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.178 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0544 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 4.158 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 18.3392 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 606.885000 389.000000 606.985000 ;
    END
  END BIAS_DBP[4]
  PIN BIAS_DBP[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.988 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4352 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 607.430000 389.000000 607.530000 ;
    END
  END BIAS_DBP[3]
  PIN BIAS_DBP[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.122 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9808 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 607.975000 389.000000 608.075000 ;
    END
  END BIAS_DBP[2]
  PIN BIAS_DBP[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.782 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 608.520000 389.000000 608.620000 ;
    END
  END BIAS_DBP[1]
  PIN BIAS_DBP[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.566 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9344 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 2.098 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2752 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 609.065000 389.000000 609.165000 ;
    END
  END BIAS_DBP[0]
  PIN BIAS_DBN[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.613 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7412 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 579.090000 389.000000 579.190000 ;
    END
  END BIAS_DBN[13]
  PIN BIAS_DBN[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.626 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1984 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 4.258 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7792 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 3.918 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2832 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 579.635000 389.000000 579.735000 ;
    END
  END BIAS_DBN[12]
  PIN BIAS_DBN[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 580.180000 389.000000 580.280000 ;
    END
  END BIAS_DBN[11]
  PIN BIAS_DBN[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.3935 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7754 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 5.998 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.4352 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 580.725000 389.000000 580.825000 ;
    END
  END BIAS_DBN[10]
  PIN BIAS_DBN[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.22 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.422 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9008 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.186 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4624 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 8.978 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 39.5472 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 581.270000 389.000000 581.370000 ;
    END
  END BIAS_DBN[9]
  PIN BIAS_DBN[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.702 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1328 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 581.815000 389.000000 581.915000 ;
    END
  END BIAS_DBN[8]
  PIN BIAS_DBN[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 582.360000 389.000000 582.460000 ;
    END
  END BIAS_DBN[7]
  PIN BIAS_DBN[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 4.658 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.5392 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 6.302 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.7728 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 3.098 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6752 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6  ;
    ANTENNAMAXAREACAR 162.882 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 719.276 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 582.905000 389.000000 583.005000 ;
    END
  END BIAS_DBN[6]
  PIN BIAS_DBN[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.458 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0592 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.138 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0512 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 583.450000 389.000000 583.550000 ;
    END
  END BIAS_DBN[5]
  PIN BIAS_DBN[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 5.964 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.3296 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 583.995000 389.000000 584.095000 ;
    END
  END BIAS_DBN[4]
  PIN BIAS_DBN[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.158 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1392 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 584.540000 389.000000 584.640000 ;
    END
  END BIAS_DBN[3]
  PIN BIAS_DBN[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.6275 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.249 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 585.085000 389.000000 585.185000 ;
    END
  END BIAS_DBN[2]
  PIN BIAS_DBN[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 8.418 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.0832 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 585.630000 389.000000 585.730000 ;
    END
  END BIAS_DBN[1]
  PIN BIAS_DBN[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.978 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3472 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 586.175000 389.000000 586.275000 ;
    END
  END BIAS_DBN[0]
  PIN BIAS_DBPC[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.858 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8192 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 594.350000 389.000000 594.450000 ;
    END
  END BIAS_DBPC[13]
  PIN BIAS_DBPC[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.2625 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.243 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 594.895000 389.000000 594.995000 ;
    END
  END BIAS_DBPC[12]
  PIN BIAS_DBPC[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.442 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 5.018 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1232 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 595.440000 389.000000 595.540000 ;
    END
  END BIAS_DBPC[11]
  PIN BIAS_DBPC[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.476 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3824 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 595.985000 389.000000 596.085000 ;
    END
  END BIAS_DBPC[10]
  PIN BIAS_DBPC[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 596.530000 389.000000 596.630000 ;
    END
  END BIAS_DBPC[9]
  PIN BIAS_DBPC[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 597.075000 389.000000 597.175000 ;
    END
  END BIAS_DBPC[8]
  PIN BIAS_DBPC[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.008 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5232 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 597.620000 389.000000 597.720000 ;
    END
  END BIAS_DBPC[7]
  PIN BIAS_DBPC[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.338 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 3.898 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1952 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 598.165000 389.000000 598.265000 ;
    END
  END BIAS_DBPC[6]
  PIN BIAS_DBPC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.302 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7728 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 598.710000 389.000000 598.810000 ;
    END
  END BIAS_DBPC[5]
  PIN BIAS_DBPC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.7105 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4142 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 599.255000 389.000000 599.355000 ;
    END
  END BIAS_DBPC[4]
  PIN BIAS_DBPC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.019 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0836 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 599.800000 389.000000 599.900000 ;
    END
  END BIAS_DBPC[3]
  PIN BIAS_DBPC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6528 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 600.345000 389.000000 600.445000 ;
    END
  END BIAS_DBPC[2]
  PIN BIAS_DBPC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 2.422 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7008 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 600.890000 389.000000 600.990000 ;
    END
  END BIAS_DBPC[1]
  PIN BIAS_DBPC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.278 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6672 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 601.435000 389.000000 601.535000 ;
    END
  END BIAS_DBPC[0]
  PIN BIAS_DBNC[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.173 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8052 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.862 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8368 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 586.720000 389.000000 586.820000 ;
    END
  END BIAS_DBNC[13]
  PIN BIAS_DBNC[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.426 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3184 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 587.265000 389.000000 587.365000 ;
    END
  END BIAS_DBNC[12]
  PIN BIAS_DBNC[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.706 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5504 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 587.810000 389.000000 587.910000 ;
    END
  END BIAS_DBNC[11]
  PIN BIAS_DBNC[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.744 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7616 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 588.355000 389.000000 588.455000 ;
    END
  END BIAS_DBNC[10]
  PIN BIAS_DBNC[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.019 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0836 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.878 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3072 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 588.900000 389.000000 589.000000 ;
    END
  END BIAS_DBNC[9]
  PIN BIAS_DBNC[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.618 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7632 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 589.445000 389.000000 589.545000 ;
    END
  END BIAS_DBNC[8]
  PIN BIAS_DBNC[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.03 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.132 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 589.990000 389.000000 590.090000 ;
    END
  END BIAS_DBNC[7]
  PIN BIAS_DBNC[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0615 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3146 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 590.535000 389.000000 590.635000 ;
    END
  END BIAS_DBNC[6]
  PIN BIAS_DBNC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 1.038 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6112 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 1.226 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4384 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 7.418 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6832 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 591.080000 389.000000 591.180000 ;
    END
  END BIAS_DBNC[5]
  PIN BIAS_DBNC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 591.625000 389.000000 591.725000 ;
    END
  END BIAS_DBNC[4]
  PIN BIAS_DBNC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6528 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 592.170000 389.000000 592.270000 ;
    END
  END BIAS_DBNC[3]
  PIN BIAS_DBNC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1105 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5302 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.918 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0832 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 592.715000 389.000000 592.815000 ;
    END
  END BIAS_DBNC[2]
  PIN BIAS_DBNC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.104 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9456 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 593.260000 389.000000 593.360000 ;
    END
  END BIAS_DBNC[1]
  PIN BIAS_DBNC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0245 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1518 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 593.805000 389.000000 593.905000 ;
    END
  END BIAS_DBNC[0]
  PIN BIAS_TC_POT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5305 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3782 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2  ;
    ANTENNAMAXAREACAR 8.27742 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 36.8629 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3  ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 10.0379 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 45.2439 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.922 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1008 LAYER M4  ;
    ANTENNAGATEAREA 0.0693 LAYER M4  ;
    ANTENNAMAXAREACAR 23.3424 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 104.418 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1052.065000 445.480000 1052.165000 446.000000 ;
    END
  END BIAS_TC_POT[5]
  PIN BIAS_TC_POT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.535 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.442 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1052.610000 445.480000 1052.710000 446.000000 ;
    END
  END BIAS_TC_POT[4]
  PIN BIAS_TC_POT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2135 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9394 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.586 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6224 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.618 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7632 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1053.155000 445.480000 1053.255000 446.000000 ;
    END
  END BIAS_TC_POT[3]
  PIN BIAS_TC_POT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3288 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.498 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2352 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1053.700000 445.480000 1053.800000 446.000000 ;
    END
  END BIAS_TC_POT[2]
  PIN BIAS_TC_POT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.2665 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2166 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 2.062 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1168 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1054.245000 445.480000 1054.345000 446.000000 ;
    END
  END BIAS_TC_POT[1]
  PIN BIAS_TC_POT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.207 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9108 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1054.790000 445.480000 1054.890000 446.000000 ;
    END
  END BIAS_TC_POT[0]
  PIN BIAS_LC_POT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1325 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.583 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.69 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.48 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 28.7482 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 126.309 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1055.335000 445.480000 1055.435000 446.000000 ;
    END
  END BIAS_LC_POT[5]
  PIN BIAS_LC_POT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.091 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.139 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6556 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 2.32 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.296 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M4  ;
    ANTENNAMAXAREACAR 85.1298 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 376.552 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.63934 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1055.880000 445.480000 1055.980000 446.000000 ;
    END
  END BIAS_LC_POT[4]
  PIN BIAS_LC_POT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.928 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.402 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2128 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 24.7583 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 108.713 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1056.425000 445.480000 1056.525000 446.000000 ;
    END
  END BIAS_LC_POT[3]
  PIN BIAS_LC_POT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.767 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3748 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M2  ;
    ANTENNAMAXAREACAR 18.357 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 78.2922 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAMAXCUTCAR 0.823045 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.858 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8192 LAYER M3  ;
    ANTENNAGATEAREA 0.0486 LAYER M3  ;
    ANTENNAMAXAREACAR 36.0113 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 156.877 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.823045 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1056.970000 445.480000 1057.070000 446.000000 ;
    END
  END BIAS_LC_POT[2]
  PIN BIAS_LC_POT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6805 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9942 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.318 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4432 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1057.515000 445.480000 1057.615000 446.000000 ;
    END
  END BIAS_LC_POT[1]
  PIN BIAS_LC_POT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6984 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1058.060000 445.480000 1058.160000 446.000000 ;
    END
  END BIAS_LC_POT[0]
  PIN BIAS_TIA_G_POT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.298 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3112 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1059.150000 445.480000 1059.250000 446.000000 ;
    END
  END BIAS_TIA_G_POT[16]
  PIN BIAS_TIA_G_POT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9965 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3846 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 2.886 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7424 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 6.678 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 29.4272 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1043.345000 445.480000 1043.445000 446.000000 ;
    END
  END BIAS_TIA_G_POT[15]
  PIN BIAS_TIA_G_POT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.087 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3828 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.726 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2384 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.562 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5168 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 3.946 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4064 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1043.890000 445.480000 1043.990000 446.000000 ;
    END
  END BIAS_TIA_G_POT[14]
  PIN BIAS_TIA_G_POT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2455 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0802 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.802 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 3.878 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1072 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1044.435000 445.480000 1044.535000 446.000000 ;
    END
  END BIAS_TIA_G_POT[13]
  PIN BIAS_TIA_G_POT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.214 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3416 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 6.542 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.8288 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1044.980000 445.480000 1045.080000 446.000000 ;
    END
  END BIAS_TIA_G_POT[12]
  PIN BIAS_TIA_G_POT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.171 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7524 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.418 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8832 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.062 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 17.9168 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 0.402 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 1045.525000 445.480000 1045.625000 446.000000 ;
    END
  END BIAS_TIA_G_POT[11]
  PIN BIAS_TIA_G_POT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.109 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8796 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 6.678 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.4272 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1046.070000 445.480000 1046.170000 446.000000 ;
    END
  END BIAS_TIA_G_POT[10]
  PIN BIAS_TIA_G_POT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3475 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.529 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.782 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1046.615000 445.480000 1046.715000 446.000000 ;
    END
  END BIAS_TIA_G_POT[9]
  PIN BIAS_TIA_G_POT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.301 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3684 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 3.202 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.1328 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1047.160000 445.480000 1047.260000 446.000000 ;
    END
  END BIAS_TIA_G_POT[8]
  PIN BIAS_TIA_G_POT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0695 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3058 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.566 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5344 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.838 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7312 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1047.705000 445.480000 1047.805000 446.000000 ;
    END
  END BIAS_TIA_G_POT[7]
  PIN BIAS_TIA_G_POT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.347 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5268 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.466 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0944 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1048.250000 445.480000 1048.350000 446.000000 ;
    END
  END BIAS_TIA_G_POT[6]
  PIN BIAS_TIA_G_POT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6974 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.446 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0064 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1048.795000 445.480000 1048.895000 446.000000 ;
    END
  END BIAS_TIA_G_POT[5]
  PIN BIAS_TIA_G_POT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.253 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1132 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.526 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1049.340000 445.480000 1049.440000 446.000000 ;
    END
  END BIAS_TIA_G_POT[4]
  PIN BIAS_TIA_G_POT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.087 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3828 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.766 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4144 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4  ;
    ANTENNAMAXAREACAR 17.7363 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 79.7518 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1049.885000 445.480000 1049.985000 446.000000 ;
    END
  END BIAS_TIA_G_POT[3]
  PIN BIAS_TIA_G_POT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.615 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.75 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2  ;
    ANTENNAMAXAREACAR 9.49675 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 42.228 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAMAXCUTCAR 0.2886 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 10.2471 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 46.1645 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.742 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3088 LAYER M4  ;
    ANTENNAGATEAREA 0.0693 LAYER M4  ;
    ANTENNAMAXAREACAR 20.9542 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 93.9105 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1050.430000 445.480000 1050.530000 446.000000 ;
    END
  END BIAS_TIA_G_POT[2]
  PIN BIAS_TIA_G_POT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0765 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3366 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.146 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 2.318 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2432 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1050.975000 445.480000 1051.075000 446.000000 ;
    END
  END BIAS_TIA_G_POT[1]
  PIN BIAS_TIA_G_POT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.278 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7112 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2  ;
    ANTENNAMAXAREACAR 19.0639 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 84.9582 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.1443 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 1051.520000 445.480000 1051.620000 446.000000 ;
    END
  END BIAS_TIA_G_POT[0]
  PIN BIAS_REV_POT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.318 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6432 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 607.010000 1139.520000 607.110000 ;
    END
  END BIAS_REV_POT[13]
  PIN BIAS_REV_POT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.868 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9072 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 607.555000 1139.520000 607.655000 ;
    END
  END BIAS_REV_POT[12]
  PIN BIAS_REV_POT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.818 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6432 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 608.100000 1139.520000 608.200000 ;
    END
  END BIAS_REV_POT[11]
  PIN BIAS_REV_POT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7465 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2846 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.606 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7104 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.938 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5712 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 608.645000 1139.520000 608.745000 ;
    END
  END BIAS_REV_POT[10]
  PIN BIAS_REV_POT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.398 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4392 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 609.190000 1139.520000 609.290000 ;
    END
  END BIAS_REV_POT[9]
  PIN BIAS_REV_POT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.138 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0512 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 609.735000 1139.520000 609.835000 ;
    END
  END BIAS_REV_POT[8]
  PIN BIAS_REV_POT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.484 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.722 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2208 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 610.280000 1139.520000 610.380000 ;
    END
  END BIAS_REV_POT[7]
  PIN BIAS_REV_POT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0215 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0946 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.678 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0272 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 610.825000 1139.520000 610.925000 ;
    END
  END BIAS_REV_POT[6]
  PIN BIAS_REV_POT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.141 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6644 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 611.370000 1139.520000 611.470000 ;
    END
  END BIAS_REV_POT[5]
  PIN BIAS_REV_POT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0705 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3102 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.662 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9568 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 611.915000 1139.520000 612.015000 ;
    END
  END BIAS_REV_POT[4]
  PIN BIAS_REV_POT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.528 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3672 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 612.460000 1139.520000 612.560000 ;
    END
  END BIAS_REV_POT[3]
  PIN BIAS_REV_POT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0245 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1518 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 613.005000 1139.520000 613.105000 ;
    END
  END BIAS_REV_POT[2]
  PIN BIAS_REV_POT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.718 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2032 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 613.550000 1139.520000 613.650000 ;
    END
  END BIAS_REV_POT[1]
  PIN BIAS_REV_POT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0845 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4158 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 614.095000 1139.520000 614.195000 ;
    END
  END BIAS_REV_POT[0]
  PIN BIAS_TC_DSADC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0174 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.738 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2912 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1019.335000 445.480000 1019.435000 446.000000 ;
    END
  END BIAS_TC_DSADC[5]
  PIN BIAS_TC_DSADC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.65 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.904 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.478 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5472 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3  ;
    ANTENNAMAXAREACAR 26.45 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 117.297 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.333333 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1019.880000 445.480000 1019.980000 446.000000 ;
    END
  END BIAS_TC_DSADC[4]
  PIN BIAS_TC_DSADC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0735 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7234 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.838 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1312 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 33.539 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 147.388 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1020.425000 445.480000 1020.525000 446.000000 ;
    END
  END BIAS_TC_DSADC[3]
  PIN BIAS_TC_DSADC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.671 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9524 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.342 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9488 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 24.715 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 108.257 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1020.970000 445.480000 1021.070000 446.000000 ;
    END
  END BIAS_TC_DSADC[2]
  PIN BIAS_TC_DSADC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6105 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6862 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.306 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7904 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1021.515000 445.480000 1021.615000 446.000000 ;
    END
  END BIAS_TC_DSADC[1]
  PIN BIAS_TC_DSADC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.045 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.642 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.182 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2448 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 24.8737 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 109.221 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1022.060000 445.480000 1022.160000 446.000000 ;
    END
  END BIAS_TC_DSADC[0]
  PIN BIAS_LC_DSADC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.1165 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0006 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.616 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1984 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3  ;
    ANTENNAMAXAREACAR 60.0332 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 264.524 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1022.605000 445.480000 1022.705000 446.000000 ;
    END
  END BIAS_LC_DSADC[5]
  PIN BIAS_LC_DSADC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 2.029 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0596 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.502 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3  ;
    ANTENNAMAXAREACAR 55.6448 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 241.042 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1023.150000 445.480000 1023.250000 446.000000 ;
    END
  END BIAS_LC_DSADC[4]
  PIN BIAS_LC_DSADC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.0215 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5386 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.822 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0608 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3  ;
    ANTENNAMAXAREACAR 68.5121 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 300.175 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1023.695000 445.480000 1023.795000 446.000000 ;
    END
  END BIAS_LC_DSADC[3]
  PIN BIAS_LC_DSADC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.49 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1024.240000 445.480000 1024.340000 446.000000 ;
    END
  END BIAS_LC_DSADC[2]
  PIN BIAS_LC_DSADC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.1155 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9522 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1024.785000 445.480000 1024.885000 446.000000 ;
    END
  END BIAS_LC_DSADC[1]
  PIN BIAS_LC_DSADC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.132 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9808 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.566 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9344 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 30.9488 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 134.231 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1025.330000 445.480000 1025.430000 446.000000 ;
    END
  END BIAS_LC_DSADC[0]
  PIN BIAS_RIN_DSADC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8162 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.542 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4288 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 1.618 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1632 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M5  ;
    ANTENNAMAXAREACAR 102.165 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 453.592 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.26537 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1016.065000 445.480000 1016.165000 446.000000 ;
    END
  END BIAS_RIN_DSADC[5]
  PIN BIAS_RIN_DSADC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.775 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.41 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.058 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6992 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3  ;
    ANTENNAMAXAREACAR 54.4628 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 240.854 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1016.610000 445.480000 1016.710000 446.000000 ;
    END
  END BIAS_RIN_DSADC[4]
  PIN BIAS_RIN_DSADC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.402 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M2  ;
    ANTENNAMAXAREACAR 48.3463 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 213.942 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.323625 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 1017.155000 445.480000 1017.255000 446.000000 ;
    END
  END BIAS_RIN_DSADC[3]
  PIN BIAS_RIN_DSADC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.118 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9632 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1017.700000 445.480000 1017.800000 446.000000 ;
    END
  END BIAS_RIN_DSADC[2]
  PIN BIAS_RIN_DSADC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8305 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6542 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.684 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4976 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3  ;
    ANTENNAMAXAREACAR 63.4595 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 281.864 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1018.245000 445.480000 1018.345000 446.000000 ;
    END
  END BIAS_RIN_DSADC[1]
  PIN BIAS_RIN_DSADC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.613 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1852 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1018.790000 445.480000 1018.890000 446.000000 ;
    END
  END BIAS_RIN_DSADC[0]
  PIN BIAS_RFB_DSADC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5346 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.962 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6768 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 LAYER M3  ;
    ANTENNAMAXAREACAR 51.7748 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 227.908 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1012.795000 445.480000 1012.895000 446.000000 ;
    END
  END BIAS_RFB_DSADC[5]
  PIN BIAS_RFB_DSADC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.153 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6732 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.442 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.502 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 21.28 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 93.72 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 1.082 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8048 LAYER M6  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6  ;
    ANTENNADIFFAREA 1.696 LAYER M7  ;
    ANTENNAPARTIALMETALAREA 3.588 LAYER M7  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8752 LAYER M7  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M7  ;
    ANTENNAMAXAREACAR 288.189 LAYER M7  ;
    ANTENNAMAXSIDEAREACAR 1260.12 LAYER M7  ;
    ANTENNAMAXCUTCAR 3.8835 LAYER VIA7  ;
    PORT
      LAYER M2 ;
        RECT 1013.340000 445.480000 1013.440000 446.000000 ;
    END
  END BIAS_RFB_DSADC[4]
  PIN BIAS_RFB_DSADC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.4415 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9866 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.762 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3968 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 LAYER M4  ;
    ANTENNAMAXAREACAR 41.6223 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 184.461 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1013.885000 445.480000 1013.985000 446.000000 ;
    END
  END BIAS_RFB_DSADC[3]
  PIN BIAS_RFB_DSADC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.085 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.374 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.958 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2592 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.246 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 1.598 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0752 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M5  ;
    ANTENNAMAXAREACAR 277.204 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 1225.4 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.589 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1014.430000 445.480000 1014.530000 446.000000 ;
    END
  END BIAS_RFB_DSADC[2]
  PIN BIAS_RFB_DSADC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3755 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6522 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.802 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5728 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4  ;
    ANTENNAMAXAREACAR 103.852 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 457.327 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1014.975000 445.480000 1015.075000 446.000000 ;
    END
  END BIAS_RFB_DSADC[1]
  PIN BIAS_RFB_DSADC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.137 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6028 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.766 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4144 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.898 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9952 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 0.226 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6  ;
    ANTENNAMAXAREACAR 441.294 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1949.05 LAYER M6  ;
    ANTENNAMAXCUTCAR 3.23625 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 1015.520000 445.480000 1015.620000 446.000000 ;
    END
  END BIAS_RFB_DSADC[0]
  PIN BIAS_DSADC_VCM[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 5.715 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.19 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 599.380000 1139.520000 599.480000 ;
    END
  END BIAS_DSADC_VCM[13]
  PIN BIAS_DSADC_VCM[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.942 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1888 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 599.925000 1139.520000 600.025000 ;
    END
  END BIAS_DSADC_VCM[12]
  PIN BIAS_DSADC_VCM[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.529 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1276 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.426 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9184 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.778 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8672 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 600.470000 1139.520000 600.570000 ;
    END
  END BIAS_DSADC_VCM[11]
  PIN BIAS_DSADC_VCM[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 601.015000 1139.520000 601.115000 ;
    END
  END BIAS_DSADC_VCM[10]
  PIN BIAS_DSADC_VCM[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.411 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4964 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 601.560000 1139.520000 601.660000 ;
    END
  END BIAS_DSADC_VCM[9]
  PIN BIAS_DSADC_VCM[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.158 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1392 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 602.105000 1139.520000 602.205000 ;
    END
  END BIAS_DSADC_VCM[8]
  PIN BIAS_DSADC_VCM[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.158 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7392 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.662 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9568 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 602.650000 1139.520000 602.750000 ;
    END
  END BIAS_DSADC_VCM[7]
  PIN BIAS_DSADC_VCM[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0625 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 603.195000 1139.520000 603.295000 ;
    END
  END BIAS_DSADC_VCM[6]
  PIN BIAS_DSADC_VCM[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.758 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3792 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 603.740000 1139.520000 603.840000 ;
    END
  END BIAS_DSADC_VCM[5]
  PIN BIAS_DSADC_VCM[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.458 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 604.285000 1139.520000 604.385000 ;
    END
  END BIAS_DSADC_VCM[4]
  PIN BIAS_DSADC_VCM[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.008 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 6.802 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 29.9728 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5  ;
    ANTENNAMAXAREACAR 102.543 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 452.277 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 604.830000 1139.520000 604.930000 ;
    END
  END BIAS_DSADC_VCM[3]
  PIN BIAS_DSADC_VCM[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0655 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3322 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 605.375000 1139.520000 605.475000 ;
    END
  END BIAS_DSADC_VCM[2]
  PIN BIAS_DSADC_VCM[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 605.920000 1139.520000 606.020000 ;
    END
  END BIAS_DSADC_VCM[1]
  PIN BIAS_DSADC_VCM[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.546 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4464 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 606.465000 1139.520000 606.565000 ;
    END
  END BIAS_DSADC_VCM[0]
  PIN dsadc_conv_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.042 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1848 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.278 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 1.402 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2128 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 12.446 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 54.8944 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0381 LAYER M5  ;
    ANTENNAMAXAREACAR 384.411 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 1684.27 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.09974 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 998.030000 445.480000 998.130000 446.000000 ;
    END
  END dsadc_conv_done
  PIN dsadc_en
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.288 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3112 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1042.800000 445.480000 1042.900000 446.000000 ;
    END
  END dsadc_en
  PIN dsadc_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2156 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 61.202 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.4982 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1027.510000 445.480000 1027.610000 446.000000 ;
    END
  END dsadc_clk
  PIN dsadc_switch[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.2695 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1858 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1025.875000 445.480000 1025.975000 446.000000 ;
    END
  END dsadc_switch[2]
  PIN dsadc_switch[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.244 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0736 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.938 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5712 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1026.420000 445.480000 1026.520000 446.000000 ;
    END
  END dsadc_switch[1]
  PIN dsadc_switch[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6225 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.739 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.862 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8368 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1026.965000 445.480000 1027.065000 446.000000 ;
    END
  END dsadc_switch[0]
  PIN dac_en_pot
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8065 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 6.026 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.5584 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1042.255000 445.480000 1042.355000 446.000000 ;
    END
  END dac_en_pot
  PIN adc_ext_in
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1012.250000 445.480000 1012.350000 446.000000 ;
    END
  END adc_ext_in
  PIN atp_en
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4445 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9558 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 7.002 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.8528 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1010.615000 445.480000 1010.715000 446.000000 ;
    END
  END atp_en
  PIN atp_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.385 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.738 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1011.160000 445.480000 1011.260000 446.000000 ;
    END
  END atp_sel
  PIN adc_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.4115 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8546 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1011.705000 445.480000 1011.805000 446.000000 ;
    END
  END adc_sel
  PIN saradc_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 9.662 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8042 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 874.605000 445.480000 874.705000 446.000000 ;
    END
  END saradc_clk
  PIN saradc_rdy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.131 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5764 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.1 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.484 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.618 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7632 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M5  ;
    ANTENNAMAXAREACAR 278.703 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 1227.84 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.30548 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 874.205000 445.480000 874.305000 446.000000 ;
    END
  END saradc_rdy
  PIN saradc_rst
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.5155 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2682 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 873.805000 445.480000 873.905000 446.000000 ;
    END
  END saradc_rst
  PIN saradc_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.087 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3828 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.8215 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6586 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 1.404 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2656 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.778 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 21.0672 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 0.606 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7104 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6  ;
    ANTENNAMAXAREACAR 195.333 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 865.486 LAYER M6  ;
    ANTENNAMAXCUTCAR 4.08163 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 873.405000 445.480000 873.505000 446.000000 ;
    END
  END saradc_data[9]
  PIN saradc_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1515 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6666 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 6.844 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.2016 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 6.678 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 29.4272 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M6  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6  ;
    ANTENNAPARTIALMETALAREA 0.946 LAYER M7  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2064 LAYER M7  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M7  ;
    ANTENNAMAXAREACAR 174.435 LAYER M7  ;
    ANTENNAMAXSIDEAREACAR 759.135 LAYER M7  ;
    ANTENNAMAXCUTCAR 4.89796 LAYER VIA7  ;
    PORT
      LAYER M2 ;
        RECT 873.005000 445.480000 873.105000 446.000000 ;
    END
  END saradc_data[8]
  PIN saradc_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3515 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5466 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.642 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8688 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.946 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2064 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 16.424 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 72.3536 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5  ;
    ANTENNAMAXAREACAR 723.796 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 3192.06 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.85714 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 872.605000 445.480000 872.705000 446.000000 ;
    END
  END saradc_data[7]
  PIN saradc_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1915 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8426 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.782 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 15.778 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 69.4672 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 1.418 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2832 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6  ;
    ANTENNAMAXAREACAR 78.0265 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 349.306 LAYER M6  ;
    ANTENNAMAXCUTCAR 4.08163 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 872.205000 445.480000 872.305000 446.000000 ;
    END
  END saradc_data[6]
  PIN saradc_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2315 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0186 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 2.026 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9584 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.222 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6208 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M5  ;
    ANTENNAMAXAREACAR 140.579 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 617.929 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.01511 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 871.805000 445.480000 871.905000 446.000000 ;
    END
  END saradc_data[5]
  PIN saradc_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7425 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.267 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.978 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3472 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 12.378 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 54.5072 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5  ;
    ANTENNAMAXAREACAR 683.186 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 2995.25 LAYER M5  ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 871.405000 445.480000 871.505000 446.000000 ;
    END
  END saradc_data[4]
  PIN saradc_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5845 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6158 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 3.558 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.6992 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.146 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 9.196 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 40.5504 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5  ;
    ANTENNAMAXAREACAR 399.659 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 1761.26 LAYER M5  ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 871.005000 445.480000 871.105000 446.000000 ;
    END
  END saradc_data[3]
  PIN saradc_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M2  ;
    ANTENNAMAXAREACAR 9.62972 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6625 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.251889 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 870.605000 445.480000 870.705000 446.000000 ;
    END
  END saradc_data[2]
  PIN saradc_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9025 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.971 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 5.762 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.3968 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 7.818 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 34.4432 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 0.622 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7808 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6  ;
    ANTENNAMAXAREACAR 206.859 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 901.796 LAYER M6  ;
    ANTENNAMAXCUTCAR 4.08163 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 870.205000 445.480000 870.305000 446.000000 ;
    END
  END saradc_data[1]
  PIN saradc_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3595 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5818 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 9.742 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.9088 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3  ;
    ANTENNAMAXAREACAR 266.826 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1167.91 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 869.805000 445.480000 869.905000 446.000000 ;
    END
  END saradc_data[0]
  PIN a0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[31]
  PIN a0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[30]
  PIN a0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[29]
  PIN a0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[28]
  PIN a0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[27]
  PIN a0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[26]
  PIN a0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[25]
  PIN a0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[24]
  PIN a0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[23]
  PIN a0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[22]
  PIN a0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[21]
  PIN a0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[20]
  PIN a0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[19]
  PIN a0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[18]
  PIN a0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[17]
  PIN a0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[16]
  PIN a0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[15]
  PIN a0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[14]
  PIN a0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[13]
  PIN a0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[12]
  PIN a0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[11]
  PIN a0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[10]
  PIN a0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[9]
  PIN a0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[8]
  PIN a0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[7]
  PIN a0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[6]
  PIN a0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[5]
  PIN a0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[4]
  PIN a0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[3]
  PIN a0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[2]
  PIN a0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[1]
  PIN a0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[0]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M7 ;
        RECT 51.000000 0.000000 56.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 51.000000 681.000000 56.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 101.000000 0.000000 106.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 101.000000 681.000000 106.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 151.000000 0.000000 156.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 151.000000 681.000000 156.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 201.000000 0.000000 206.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 201.000000 681.000000 206.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 251.000000 0.000000 256.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 251.000000 681.000000 256.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 301.000000 0.000000 306.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 301.000000 681.000000 306.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 351.000000 0.000000 356.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 351.000000 681.000000 356.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 401.000000 0.000000 406.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 401.000000 501.000000 406.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 401.000000 656.000000 406.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 401.000000 681.000000 406.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 451.000000 0.000000 456.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 451.000000 501.000000 456.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 451.000000 656.000000 456.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 451.000000 681.000000 456.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 501.000000 0.000000 506.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 501.000000 501.000000 506.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 501.000000 656.000000 506.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 501.000000 681.000000 506.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 551.000000 0.000000 556.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 551.000000 501.000000 556.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 551.000000 656.000000 556.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 551.000000 681.000000 556.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 601.000000 0.000000 606.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 601.000000 501.000000 606.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 601.000000 656.000000 606.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 601.000000 681.000000 606.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 651.000000 0.000000 656.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 651.000000 501.000000 656.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 651.000000 656.000000 656.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 651.000000 681.000000 656.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 701.000000 0.000000 706.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 701.000000 501.000000 706.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 751.000000 0.000000 756.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 751.000000 441.000000 756.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 801.000000 0.000000 806.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 801.000000 441.000000 806.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 851.000000 0.000000 856.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 851.000000 441.000000 856.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 901.000000 0.000000 906.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 901.000000 441.000000 906.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 951.000000 0.000000 956.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 951.000000 441.000000 956.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1001.000000 0.000000 1006.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1001.000000 441.000000 1006.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1051.000000 0.000000 1056.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1051.000000 441.000000 1056.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1101.000000 0.000000 1106.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1101.000000 441.000000 1106.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1151.000000 0.000000 1156.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1151.000000 681.000000 1156.000000 686.000000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER M2 ;
        RECT 4.000000 5.850000 14.000000 6.150000 ;
        RECT 51.000000 5.850000 56.000000 6.150000 ;
        RECT 51.000000 1.850000 56.000000 2.150000 ;
        RECT 101.000000 1.850000 106.000000 2.150000 ;
        RECT 101.000000 5.850000 106.000000 6.150000 ;
        RECT 151.000000 1.850000 156.000000 2.150000 ;
        RECT 151.000000 5.850000 156.000000 6.150000 ;
        RECT 201.000000 1.850000 206.000000 2.150000 ;
        RECT 201.000000 5.850000 206.000000 6.150000 ;
        RECT 251.000000 1.850000 256.000000 2.150000 ;
        RECT 251.000000 5.850000 256.000000 6.150000 ;
        RECT 301.000000 1.850000 306.000000 2.150000 ;
        RECT 301.000000 5.850000 306.000000 6.150000 ;
        RECT 351.000000 1.850000 356.000000 2.150000 ;
        RECT 351.000000 5.850000 356.000000 6.150000 ;
        RECT 401.000000 1.850000 406.000000 2.150000 ;
        RECT 401.000000 5.850000 406.000000 6.150000 ;
        RECT 451.000000 1.850000 456.000000 2.150000 ;
        RECT 451.000000 5.850000 456.000000 6.150000 ;
        RECT 501.000000 1.850000 506.000000 2.150000 ;
        RECT 501.000000 5.850000 506.000000 6.150000 ;
        RECT 551.000000 1.850000 556.000000 2.150000 ;
        RECT 551.000000 5.850000 556.000000 6.150000 ;
        RECT 4.000000 265.850000 14.000000 266.150000 ;
        RECT 4.000000 261.850000 14.000000 262.150000 ;
        RECT 51.000000 265.850000 56.000000 266.150000 ;
        RECT 51.000000 261.850000 56.000000 262.150000 ;
        RECT 101.000000 265.850000 106.000000 266.150000 ;
        RECT 101.000000 261.850000 106.000000 262.150000 ;
        RECT 51.000000 305.850000 56.000000 306.150000 ;
        RECT 4.000000 305.850000 14.000000 306.150000 ;
        RECT 4.000000 285.850000 14.000000 286.150000 ;
        RECT 4.000000 281.850000 14.000000 282.150000 ;
        RECT 4.000000 269.850000 14.000000 270.150000 ;
        RECT 4.000000 273.850000 14.000000 274.150000 ;
        RECT 4.000000 277.850000 14.000000 278.150000 ;
        RECT 4.000000 289.850000 14.000000 290.150000 ;
        RECT 4.000000 293.850000 14.000000 294.150000 ;
        RECT 4.000000 297.850000 14.000000 298.150000 ;
        RECT 4.000000 301.850000 14.000000 302.150000 ;
        RECT 51.000000 269.850000 56.000000 270.150000 ;
        RECT 51.000000 273.850000 56.000000 274.150000 ;
        RECT 51.000000 277.850000 56.000000 278.150000 ;
        RECT 51.000000 281.850000 56.000000 282.150000 ;
        RECT 51.000000 285.850000 56.000000 286.150000 ;
        RECT 51.000000 301.850000 56.000000 302.150000 ;
        RECT 51.000000 297.850000 56.000000 298.150000 ;
        RECT 51.000000 293.850000 56.000000 294.150000 ;
        RECT 51.000000 289.850000 56.000000 290.150000 ;
        RECT 4.000000 321.850000 14.000000 322.150000 ;
        RECT 4.000000 317.850000 14.000000 318.150000 ;
        RECT 4.000000 309.850000 14.000000 310.150000 ;
        RECT 4.000000 313.850000 14.000000 314.150000 ;
        RECT 4.000000 325.850000 14.000000 326.150000 ;
        RECT 4.000000 329.850000 14.000000 330.150000 ;
        RECT 4.000000 333.850000 14.000000 334.150000 ;
        RECT 4.000000 337.850000 14.000000 338.150000 ;
        RECT 4.000000 341.850000 14.000000 342.150000 ;
        RECT 51.000000 313.850000 56.000000 314.150000 ;
        RECT 51.000000 309.850000 56.000000 310.150000 ;
        RECT 51.000000 317.850000 56.000000 318.150000 ;
        RECT 51.000000 321.850000 56.000000 322.150000 ;
        RECT 51.000000 341.850000 56.000000 342.150000 ;
        RECT 51.000000 337.850000 56.000000 338.150000 ;
        RECT 51.000000 333.850000 56.000000 334.150000 ;
        RECT 51.000000 329.850000 56.000000 330.150000 ;
        RECT 51.000000 325.850000 56.000000 326.150000 ;
        RECT 101.000000 305.850000 106.000000 306.150000 ;
        RECT 101.000000 285.850000 106.000000 286.150000 ;
        RECT 101.000000 269.850000 106.000000 270.150000 ;
        RECT 101.000000 273.850000 106.000000 274.150000 ;
        RECT 101.000000 277.850000 106.000000 278.150000 ;
        RECT 101.000000 281.850000 106.000000 282.150000 ;
        RECT 101.000000 301.850000 106.000000 302.150000 ;
        RECT 101.000000 297.850000 106.000000 298.150000 ;
        RECT 101.000000 293.850000 106.000000 294.150000 ;
        RECT 101.000000 289.850000 106.000000 290.150000 ;
        RECT 101.000000 321.850000 106.000000 322.150000 ;
        RECT 101.000000 317.850000 106.000000 318.150000 ;
        RECT 101.000000 313.850000 106.000000 314.150000 ;
        RECT 101.000000 309.850000 106.000000 310.150000 ;
        RECT 101.000000 325.850000 106.000000 326.150000 ;
        RECT 101.000000 329.850000 106.000000 330.150000 ;
        RECT 101.000000 333.850000 106.000000 334.150000 ;
        RECT 101.000000 337.850000 106.000000 338.150000 ;
        RECT 101.000000 341.850000 106.000000 342.150000 ;
        RECT 151.000000 261.850000 156.000000 262.150000 ;
        RECT 151.000000 265.850000 156.000000 266.150000 ;
        RECT 201.000000 265.850000 206.000000 266.150000 ;
        RECT 201.000000 261.850000 206.000000 262.150000 ;
        RECT 251.000000 265.850000 256.000000 266.150000 ;
        RECT 251.000000 261.850000 256.000000 262.150000 ;
        RECT 201.000000 305.850000 206.000000 306.150000 ;
        RECT 151.000000 305.850000 156.000000 306.150000 ;
        RECT 151.000000 277.850000 156.000000 278.150000 ;
        RECT 151.000000 273.850000 156.000000 274.150000 ;
        RECT 151.000000 269.850000 156.000000 270.150000 ;
        RECT 151.000000 281.850000 156.000000 282.150000 ;
        RECT 151.000000 285.850000 156.000000 286.150000 ;
        RECT 151.000000 289.850000 156.000000 290.150000 ;
        RECT 151.000000 293.850000 156.000000 294.150000 ;
        RECT 151.000000 301.850000 156.000000 302.150000 ;
        RECT 151.000000 297.850000 156.000000 298.150000 ;
        RECT 201.000000 269.850000 206.000000 270.150000 ;
        RECT 201.000000 273.850000 206.000000 274.150000 ;
        RECT 201.000000 277.850000 206.000000 278.150000 ;
        RECT 201.000000 281.850000 206.000000 282.150000 ;
        RECT 201.000000 285.850000 206.000000 286.150000 ;
        RECT 201.000000 301.850000 206.000000 302.150000 ;
        RECT 201.000000 297.850000 206.000000 298.150000 ;
        RECT 201.000000 293.850000 206.000000 294.150000 ;
        RECT 201.000000 289.850000 206.000000 290.150000 ;
        RECT 151.000000 313.850000 156.000000 314.150000 ;
        RECT 151.000000 309.850000 156.000000 310.150000 ;
        RECT 151.000000 321.850000 156.000000 322.150000 ;
        RECT 151.000000 317.850000 156.000000 318.150000 ;
        RECT 151.000000 329.850000 156.000000 330.150000 ;
        RECT 151.000000 325.850000 156.000000 326.150000 ;
        RECT 151.000000 333.850000 156.000000 334.150000 ;
        RECT 151.000000 337.850000 156.000000 338.150000 ;
        RECT 151.000000 341.850000 156.000000 342.150000 ;
        RECT 201.000000 313.850000 206.000000 314.150000 ;
        RECT 201.000000 309.850000 206.000000 310.150000 ;
        RECT 201.000000 317.850000 206.000000 318.150000 ;
        RECT 201.000000 321.850000 206.000000 322.150000 ;
        RECT 201.000000 341.850000 206.000000 342.150000 ;
        RECT 201.000000 337.850000 206.000000 338.150000 ;
        RECT 201.000000 333.850000 206.000000 334.150000 ;
        RECT 201.000000 329.850000 206.000000 330.150000 ;
        RECT 201.000000 325.850000 206.000000 326.150000 ;
        RECT 251.000000 305.850000 256.000000 306.150000 ;
        RECT 251.000000 285.850000 256.000000 286.150000 ;
        RECT 251.000000 269.850000 256.000000 270.150000 ;
        RECT 251.000000 273.850000 256.000000 274.150000 ;
        RECT 251.000000 277.850000 256.000000 278.150000 ;
        RECT 251.000000 281.850000 256.000000 282.150000 ;
        RECT 251.000000 293.850000 256.000000 294.150000 ;
        RECT 251.000000 289.850000 256.000000 290.150000 ;
        RECT 251.000000 297.850000 256.000000 298.150000 ;
        RECT 251.000000 301.850000 256.000000 302.150000 ;
        RECT 251.000000 309.850000 256.000000 310.150000 ;
        RECT 251.000000 313.850000 256.000000 314.150000 ;
        RECT 251.000000 321.850000 256.000000 322.150000 ;
        RECT 251.000000 317.850000 256.000000 318.150000 ;
        RECT 251.000000 325.850000 256.000000 326.150000 ;
        RECT 251.000000 329.850000 256.000000 330.150000 ;
        RECT 251.000000 333.850000 256.000000 334.150000 ;
        RECT 251.000000 337.850000 256.000000 338.150000 ;
        RECT 251.000000 341.850000 256.000000 342.150000 ;
        RECT 301.000000 265.850000 306.000000 266.150000 ;
        RECT 301.000000 261.850000 306.000000 262.150000 ;
        RECT 351.000000 265.850000 356.000000 266.150000 ;
        RECT 351.000000 261.850000 356.000000 262.150000 ;
        RECT 401.000000 261.850000 406.000000 262.150000 ;
        RECT 401.000000 265.850000 406.000000 266.150000 ;
        RECT 301.000000 305.850000 306.000000 306.150000 ;
        RECT 351.000000 305.850000 356.000000 306.150000 ;
        RECT 301.000000 277.850000 306.000000 278.150000 ;
        RECT 301.000000 269.850000 306.000000 270.150000 ;
        RECT 301.000000 273.850000 306.000000 274.150000 ;
        RECT 301.000000 281.850000 306.000000 282.150000 ;
        RECT 301.000000 285.850000 306.000000 286.150000 ;
        RECT 301.000000 293.850000 306.000000 294.150000 ;
        RECT 301.000000 289.850000 306.000000 290.150000 ;
        RECT 301.000000 301.850000 306.000000 302.150000 ;
        RECT 301.000000 297.850000 306.000000 298.150000 ;
        RECT 351.000000 269.850000 356.000000 270.150000 ;
        RECT 351.000000 273.850000 356.000000 274.150000 ;
        RECT 351.000000 277.850000 356.000000 278.150000 ;
        RECT 351.000000 281.850000 356.000000 282.150000 ;
        RECT 351.000000 285.850000 356.000000 286.150000 ;
        RECT 351.000000 289.850000 356.000000 290.150000 ;
        RECT 351.000000 293.850000 356.000000 294.150000 ;
        RECT 351.000000 297.850000 356.000000 298.150000 ;
        RECT 351.000000 301.850000 356.000000 302.150000 ;
        RECT 301.000000 313.850000 306.000000 314.150000 ;
        RECT 301.000000 309.850000 306.000000 310.150000 ;
        RECT 301.000000 317.850000 306.000000 318.150000 ;
        RECT 301.000000 321.850000 306.000000 322.150000 ;
        RECT 301.000000 329.850000 306.000000 330.150000 ;
        RECT 301.000000 325.850000 306.000000 326.150000 ;
        RECT 301.000000 341.850000 306.000000 342.150000 ;
        RECT 301.000000 337.850000 306.000000 338.150000 ;
        RECT 301.000000 333.850000 306.000000 334.150000 ;
        RECT 351.000000 313.850000 356.000000 314.150000 ;
        RECT 351.000000 309.850000 356.000000 310.150000 ;
        RECT 351.000000 317.850000 356.000000 318.150000 ;
        RECT 351.000000 321.850000 356.000000 322.150000 ;
        RECT 351.000000 341.850000 356.000000 342.150000 ;
        RECT 351.000000 337.850000 356.000000 338.150000 ;
        RECT 351.000000 333.850000 356.000000 334.150000 ;
        RECT 351.000000 329.850000 356.000000 330.150000 ;
        RECT 351.000000 325.850000 356.000000 326.150000 ;
        RECT 401.000000 305.850000 406.000000 306.150000 ;
        RECT 401.000000 285.850000 406.000000 286.150000 ;
        RECT 401.000000 273.850000 406.000000 274.150000 ;
        RECT 401.000000 269.850000 406.000000 270.150000 ;
        RECT 401.000000 277.850000 406.000000 278.150000 ;
        RECT 401.000000 281.850000 406.000000 282.150000 ;
        RECT 401.000000 293.850000 406.000000 294.150000 ;
        RECT 401.000000 289.850000 406.000000 290.150000 ;
        RECT 401.000000 297.850000 406.000000 298.150000 ;
        RECT 401.000000 301.850000 406.000000 302.150000 ;
        RECT 401.000000 309.850000 406.000000 310.150000 ;
        RECT 401.000000 313.850000 406.000000 314.150000 ;
        RECT 401.000000 317.850000 406.000000 318.150000 ;
        RECT 401.000000 321.850000 406.000000 322.150000 ;
        RECT 401.000000 329.850000 406.000000 330.150000 ;
        RECT 401.000000 325.850000 406.000000 326.150000 ;
        RECT 401.000000 333.850000 406.000000 334.150000 ;
        RECT 401.000000 337.850000 406.000000 338.150000 ;
        RECT 401.000000 341.850000 406.000000 342.150000 ;
        RECT 451.000000 265.850000 456.000000 266.150000 ;
        RECT 451.000000 261.850000 456.000000 262.150000 ;
        RECT 501.000000 261.850000 506.000000 262.150000 ;
        RECT 501.000000 265.850000 506.000000 266.150000 ;
        RECT 551.000000 265.850000 556.000000 266.150000 ;
        RECT 551.000000 261.850000 556.000000 262.150000 ;
        RECT 501.000000 305.850000 506.000000 306.150000 ;
        RECT 451.000000 277.850000 456.000000 278.150000 ;
        RECT 451.000000 273.850000 456.000000 274.150000 ;
        RECT 451.000000 269.850000 456.000000 270.150000 ;
        RECT 451.000000 285.850000 456.000000 286.150000 ;
        RECT 451.000000 281.850000 456.000000 282.150000 ;
        RECT 451.000000 293.850000 456.000000 294.150000 ;
        RECT 451.000000 289.850000 456.000000 290.150000 ;
        RECT 451.000000 297.850000 456.000000 298.150000 ;
        RECT 501.000000 277.850000 506.000000 278.150000 ;
        RECT 501.000000 269.850000 506.000000 270.150000 ;
        RECT 501.000000 273.850000 506.000000 274.150000 ;
        RECT 501.000000 281.850000 506.000000 282.150000 ;
        RECT 501.000000 285.850000 506.000000 286.150000 ;
        RECT 501.000000 289.850000 506.000000 290.150000 ;
        RECT 501.000000 293.850000 506.000000 294.150000 ;
        RECT 501.000000 301.850000 506.000000 302.150000 ;
        RECT 501.000000 297.850000 506.000000 298.150000 ;
        RECT 451.000000 321.850000 456.000000 322.150000 ;
        RECT 451.000000 333.850000 456.000000 334.150000 ;
        RECT 451.000000 329.850000 456.000000 330.150000 ;
        RECT 451.000000 325.850000 456.000000 326.150000 ;
        RECT 451.000000 337.850000 456.000000 338.150000 ;
        RECT 451.000000 341.850000 456.000000 342.150000 ;
        RECT 501.000000 313.850000 506.000000 314.150000 ;
        RECT 501.000000 309.850000 506.000000 310.150000 ;
        RECT 501.000000 317.850000 506.000000 318.150000 ;
        RECT 501.000000 321.850000 506.000000 322.150000 ;
        RECT 501.000000 329.850000 506.000000 330.150000 ;
        RECT 501.000000 325.850000 506.000000 326.150000 ;
        RECT 501.000000 333.850000 506.000000 334.150000 ;
        RECT 501.000000 337.850000 506.000000 338.150000 ;
        RECT 501.000000 341.850000 506.000000 342.150000 ;
        RECT 551.000000 305.850000 556.000000 306.150000 ;
        RECT 551.000000 277.850000 556.000000 278.150000 ;
        RECT 551.000000 269.850000 556.000000 270.150000 ;
        RECT 551.000000 273.850000 556.000000 274.150000 ;
        RECT 551.000000 285.850000 556.000000 286.150000 ;
        RECT 551.000000 281.850000 556.000000 282.150000 ;
        RECT 551.000000 301.850000 556.000000 302.150000 ;
        RECT 551.000000 297.850000 556.000000 298.150000 ;
        RECT 551.000000 293.850000 556.000000 294.150000 ;
        RECT 551.000000 289.850000 556.000000 290.150000 ;
        RECT 551.000000 309.850000 556.000000 310.150000 ;
        RECT 551.000000 313.850000 556.000000 314.150000 ;
        RECT 551.000000 317.850000 556.000000 318.150000 ;
        RECT 551.000000 321.850000 556.000000 322.150000 ;
        RECT 551.000000 325.850000 556.000000 326.150000 ;
        RECT 551.000000 329.850000 556.000000 330.150000 ;
        RECT 551.000000 333.850000 556.000000 334.150000 ;
        RECT 551.000000 337.850000 556.000000 338.150000 ;
        RECT 551.000000 341.850000 556.000000 342.150000 ;
        RECT 601.000000 1.850000 606.000000 2.150000 ;
        RECT 601.000000 5.850000 606.000000 6.150000 ;
        RECT 651.000000 1.850000 656.000000 2.150000 ;
        RECT 651.000000 5.850000 656.000000 6.150000 ;
        RECT 701.000000 1.850000 706.000000 2.150000 ;
        RECT 701.000000 5.850000 706.000000 6.150000 ;
        RECT 751.000000 1.850000 756.000000 2.150000 ;
        RECT 751.000000 5.850000 756.000000 6.150000 ;
        RECT 801.000000 1.850000 806.000000 2.150000 ;
        RECT 801.000000 5.850000 806.000000 6.150000 ;
        RECT 851.000000 1.850000 856.000000 2.150000 ;
        RECT 851.000000 5.850000 856.000000 6.150000 ;
        RECT 901.000000 1.850000 906.000000 2.150000 ;
        RECT 901.000000 5.850000 906.000000 6.150000 ;
        RECT 951.000000 1.850000 956.000000 2.150000 ;
        RECT 951.000000 5.850000 956.000000 6.150000 ;
        RECT 1001.000000 1.850000 1006.000000 2.150000 ;
        RECT 1001.000000 5.850000 1006.000000 6.150000 ;
        RECT 1051.000000 1.850000 1056.000000 2.150000 ;
        RECT 1051.000000 5.850000 1056.000000 6.150000 ;
        RECT 1101.000000 1.850000 1106.000000 2.150000 ;
        RECT 1101.000000 5.850000 1106.000000 6.150000 ;
        RECT 1151.000000 5.850000 1156.000000 6.150000 ;
        RECT 1172.000000 5.850000 1182.000000 6.150000 ;
        RECT 1151.000000 1.850000 1156.000000 2.150000 ;
        RECT 1172.000000 17.850000 1182.000000 18.150000 ;
        RECT 1172.000000 13.850000 1182.000000 14.150000 ;
        RECT 1172.000000 9.850000 1182.000000 10.150000 ;
        RECT 1172.000000 21.850000 1182.000000 22.150000 ;
        RECT 1172.000000 25.850000 1182.000000 26.150000 ;
        RECT 1172.000000 33.850000 1182.000000 34.150000 ;
        RECT 1172.000000 29.850000 1182.000000 30.150000 ;
        RECT 1172.000000 41.850000 1182.000000 42.150000 ;
        RECT 1172.000000 37.850000 1182.000000 38.150000 ;
        RECT 1172.000000 45.850000 1182.000000 46.150000 ;
        RECT 601.000000 265.850000 606.000000 266.150000 ;
        RECT 601.000000 261.850000 606.000000 262.150000 ;
        RECT 651.000000 261.850000 656.000000 262.150000 ;
        RECT 651.000000 265.850000 656.000000 266.150000 ;
        RECT 701.000000 265.850000 706.000000 266.150000 ;
        RECT 701.000000 261.850000 706.000000 262.150000 ;
        RECT 601.000000 305.850000 606.000000 306.150000 ;
        RECT 651.000000 305.850000 656.000000 306.150000 ;
        RECT 601.000000 277.850000 606.000000 278.150000 ;
        RECT 601.000000 269.850000 606.000000 270.150000 ;
        RECT 601.000000 273.850000 606.000000 274.150000 ;
        RECT 601.000000 281.850000 606.000000 282.150000 ;
        RECT 601.000000 285.850000 606.000000 286.150000 ;
        RECT 601.000000 289.850000 606.000000 290.150000 ;
        RECT 601.000000 293.850000 606.000000 294.150000 ;
        RECT 601.000000 297.850000 606.000000 298.150000 ;
        RECT 601.000000 301.850000 606.000000 302.150000 ;
        RECT 651.000000 277.850000 656.000000 278.150000 ;
        RECT 651.000000 273.850000 656.000000 274.150000 ;
        RECT 651.000000 269.850000 656.000000 270.150000 ;
        RECT 651.000000 281.850000 656.000000 282.150000 ;
        RECT 651.000000 285.850000 656.000000 286.150000 ;
        RECT 651.000000 289.850000 656.000000 290.150000 ;
        RECT 651.000000 293.850000 656.000000 294.150000 ;
        RECT 651.000000 301.850000 656.000000 302.150000 ;
        RECT 651.000000 297.850000 656.000000 298.150000 ;
        RECT 601.000000 321.850000 606.000000 322.150000 ;
        RECT 601.000000 317.850000 606.000000 318.150000 ;
        RECT 601.000000 309.850000 606.000000 310.150000 ;
        RECT 601.000000 313.850000 606.000000 314.150000 ;
        RECT 601.000000 325.850000 606.000000 326.150000 ;
        RECT 601.000000 329.850000 606.000000 330.150000 ;
        RECT 601.000000 333.850000 606.000000 334.150000 ;
        RECT 601.000000 337.850000 606.000000 338.150000 ;
        RECT 601.000000 341.850000 606.000000 342.150000 ;
        RECT 651.000000 313.850000 656.000000 314.150000 ;
        RECT 651.000000 309.850000 656.000000 310.150000 ;
        RECT 651.000000 321.850000 656.000000 322.150000 ;
        RECT 651.000000 317.850000 656.000000 318.150000 ;
        RECT 651.000000 329.850000 656.000000 330.150000 ;
        RECT 651.000000 325.850000 656.000000 326.150000 ;
        RECT 651.000000 333.850000 656.000000 334.150000 ;
        RECT 651.000000 337.850000 656.000000 338.150000 ;
        RECT 651.000000 341.850000 656.000000 342.150000 ;
        RECT 701.000000 305.850000 706.000000 306.150000 ;
        RECT 701.000000 281.850000 706.000000 282.150000 ;
        RECT 701.000000 277.850000 706.000000 278.150000 ;
        RECT 701.000000 273.850000 706.000000 274.150000 ;
        RECT 701.000000 269.850000 706.000000 270.150000 ;
        RECT 701.000000 285.850000 706.000000 286.150000 ;
        RECT 701.000000 301.850000 706.000000 302.150000 ;
        RECT 701.000000 297.850000 706.000000 298.150000 ;
        RECT 701.000000 293.850000 706.000000 294.150000 ;
        RECT 701.000000 289.850000 706.000000 290.150000 ;
        RECT 701.000000 309.850000 706.000000 310.150000 ;
        RECT 701.000000 313.850000 706.000000 314.150000 ;
        RECT 701.000000 317.850000 706.000000 318.150000 ;
        RECT 701.000000 321.850000 706.000000 322.150000 ;
        RECT 701.000000 325.850000 706.000000 326.150000 ;
        RECT 701.000000 329.850000 706.000000 330.150000 ;
        RECT 701.000000 333.850000 706.000000 334.150000 ;
        RECT 701.000000 337.850000 706.000000 338.150000 ;
        RECT 701.000000 341.850000 706.000000 342.150000 ;
        RECT 751.000000 261.850000 756.000000 262.150000 ;
        RECT 751.000000 265.850000 756.000000 266.150000 ;
        RECT 801.000000 261.850000 806.000000 262.150000 ;
        RECT 801.000000 265.850000 806.000000 266.150000 ;
        RECT 851.000000 265.850000 856.000000 266.150000 ;
        RECT 851.000000 261.850000 856.000000 262.150000 ;
        RECT 801.000000 305.850000 806.000000 306.150000 ;
        RECT 751.000000 305.850000 756.000000 306.150000 ;
        RECT 751.000000 285.850000 756.000000 286.150000 ;
        RECT 751.000000 281.850000 756.000000 282.150000 ;
        RECT 751.000000 269.850000 756.000000 270.150000 ;
        RECT 751.000000 273.850000 756.000000 274.150000 ;
        RECT 751.000000 277.850000 756.000000 278.150000 ;
        RECT 751.000000 289.850000 756.000000 290.150000 ;
        RECT 751.000000 293.850000 756.000000 294.150000 ;
        RECT 751.000000 297.850000 756.000000 298.150000 ;
        RECT 751.000000 301.850000 756.000000 302.150000 ;
        RECT 801.000000 277.850000 806.000000 278.150000 ;
        RECT 801.000000 269.850000 806.000000 270.150000 ;
        RECT 801.000000 273.850000 806.000000 274.150000 ;
        RECT 801.000000 281.850000 806.000000 282.150000 ;
        RECT 801.000000 285.850000 806.000000 286.150000 ;
        RECT 801.000000 289.850000 806.000000 290.150000 ;
        RECT 801.000000 293.850000 806.000000 294.150000 ;
        RECT 801.000000 301.850000 806.000000 302.150000 ;
        RECT 801.000000 297.850000 806.000000 298.150000 ;
        RECT 751.000000 321.850000 756.000000 322.150000 ;
        RECT 751.000000 317.850000 756.000000 318.150000 ;
        RECT 751.000000 309.850000 756.000000 310.150000 ;
        RECT 751.000000 313.850000 756.000000 314.150000 ;
        RECT 751.000000 325.850000 756.000000 326.150000 ;
        RECT 751.000000 329.850000 756.000000 330.150000 ;
        RECT 751.000000 333.850000 756.000000 334.150000 ;
        RECT 751.000000 337.850000 756.000000 338.150000 ;
        RECT 751.000000 341.850000 756.000000 342.150000 ;
        RECT 801.000000 313.850000 806.000000 314.150000 ;
        RECT 801.000000 309.850000 806.000000 310.150000 ;
        RECT 801.000000 321.850000 806.000000 322.150000 ;
        RECT 801.000000 317.850000 806.000000 318.150000 ;
        RECT 801.000000 329.850000 806.000000 330.150000 ;
        RECT 801.000000 325.850000 806.000000 326.150000 ;
        RECT 801.000000 333.850000 806.000000 334.150000 ;
        RECT 801.000000 337.850000 806.000000 338.150000 ;
        RECT 801.000000 341.850000 806.000000 342.150000 ;
        RECT 851.000000 305.850000 856.000000 306.150000 ;
        RECT 851.000000 281.850000 856.000000 282.150000 ;
        RECT 851.000000 277.850000 856.000000 278.150000 ;
        RECT 851.000000 273.850000 856.000000 274.150000 ;
        RECT 851.000000 269.850000 856.000000 270.150000 ;
        RECT 851.000000 285.850000 856.000000 286.150000 ;
        RECT 851.000000 301.850000 856.000000 302.150000 ;
        RECT 851.000000 297.850000 856.000000 298.150000 ;
        RECT 851.000000 293.850000 856.000000 294.150000 ;
        RECT 851.000000 289.850000 856.000000 290.150000 ;
        RECT 851.000000 309.850000 856.000000 310.150000 ;
        RECT 851.000000 313.850000 856.000000 314.150000 ;
        RECT 851.000000 317.850000 856.000000 318.150000 ;
        RECT 851.000000 321.850000 856.000000 322.150000 ;
        RECT 851.000000 325.850000 856.000000 326.150000 ;
        RECT 851.000000 329.850000 856.000000 330.150000 ;
        RECT 851.000000 333.850000 856.000000 334.150000 ;
        RECT 851.000000 337.850000 856.000000 338.150000 ;
        RECT 851.000000 341.850000 856.000000 342.150000 ;
        RECT 1172.000000 61.850000 1182.000000 62.150000 ;
        RECT 1172.000000 57.850000 1182.000000 58.150000 ;
        RECT 1172.000000 53.850000 1182.000000 54.150000 ;
        RECT 1172.000000 49.850000 1182.000000 50.150000 ;
        RECT 1172.000000 73.850000 1182.000000 74.150000 ;
        RECT 1172.000000 69.850000 1182.000000 70.150000 ;
        RECT 1172.000000 65.850000 1182.000000 66.150000 ;
        RECT 1172.000000 77.850000 1182.000000 78.150000 ;
        RECT 1172.000000 81.850000 1182.000000 82.150000 ;
        RECT 1172.000000 101.850000 1182.000000 102.150000 ;
        RECT 1172.000000 89.850000 1182.000000 90.150000 ;
        RECT 1172.000000 85.850000 1182.000000 86.150000 ;
        RECT 1172.000000 93.850000 1182.000000 94.150000 ;
        RECT 1172.000000 97.850000 1182.000000 98.150000 ;
        RECT 1172.000000 117.850000 1182.000000 118.150000 ;
        RECT 1172.000000 113.850000 1182.000000 114.150000 ;
        RECT 1172.000000 105.850000 1182.000000 106.150000 ;
        RECT 1172.000000 109.850000 1182.000000 110.150000 ;
        RECT 1151.000000 133.850000 1156.000000 134.150000 ;
        RECT 1172.000000 129.850000 1182.000000 130.150000 ;
        RECT 1172.000000 125.850000 1182.000000 126.150000 ;
        RECT 1172.000000 121.850000 1182.000000 122.150000 ;
        RECT 1172.000000 133.850000 1182.000000 134.150000 ;
        RECT 1172.000000 137.850000 1182.000000 138.150000 ;
        RECT 1172.000000 141.850000 1182.000000 142.150000 ;
        RECT 1172.000000 145.850000 1182.000000 146.150000 ;
        RECT 1172.000000 149.850000 1182.000000 150.150000 ;
        RECT 1172.000000 153.850000 1182.000000 154.150000 ;
        RECT 1172.000000 165.850000 1182.000000 166.150000 ;
        RECT 1172.000000 161.850000 1182.000000 162.150000 ;
        RECT 1172.000000 157.850000 1182.000000 158.150000 ;
        RECT 1172.000000 169.850000 1182.000000 170.150000 ;
        RECT 1172.000000 173.850000 1182.000000 174.150000 ;
        RECT 1172.000000 177.850000 1182.000000 178.150000 ;
        RECT 1172.000000 181.850000 1182.000000 182.150000 ;
        RECT 1172.000000 185.850000 1182.000000 186.150000 ;
        RECT 1172.000000 189.850000 1182.000000 190.150000 ;
        RECT 1172.000000 193.850000 1182.000000 194.150000 ;
        RECT 901.000000 261.850000 906.000000 262.150000 ;
        RECT 901.000000 265.850000 906.000000 266.150000 ;
        RECT 951.000000 265.850000 956.000000 266.150000 ;
        RECT 951.000000 261.850000 956.000000 262.150000 ;
        RECT 1001.000000 261.850000 1006.000000 262.150000 ;
        RECT 1001.000000 265.850000 1006.000000 266.150000 ;
        RECT 951.000000 305.850000 956.000000 306.150000 ;
        RECT 901.000000 305.850000 906.000000 306.150000 ;
        RECT 901.000000 285.850000 906.000000 286.150000 ;
        RECT 901.000000 281.850000 906.000000 282.150000 ;
        RECT 901.000000 269.850000 906.000000 270.150000 ;
        RECT 901.000000 273.850000 906.000000 274.150000 ;
        RECT 901.000000 277.850000 906.000000 278.150000 ;
        RECT 901.000000 289.850000 906.000000 290.150000 ;
        RECT 901.000000 293.850000 906.000000 294.150000 ;
        RECT 901.000000 297.850000 906.000000 298.150000 ;
        RECT 901.000000 301.850000 906.000000 302.150000 ;
        RECT 951.000000 269.850000 956.000000 270.150000 ;
        RECT 951.000000 273.850000 956.000000 274.150000 ;
        RECT 951.000000 277.850000 956.000000 278.150000 ;
        RECT 951.000000 281.850000 956.000000 282.150000 ;
        RECT 951.000000 285.850000 956.000000 286.150000 ;
        RECT 951.000000 301.850000 956.000000 302.150000 ;
        RECT 951.000000 297.850000 956.000000 298.150000 ;
        RECT 951.000000 293.850000 956.000000 294.150000 ;
        RECT 951.000000 289.850000 956.000000 290.150000 ;
        RECT 901.000000 321.850000 906.000000 322.150000 ;
        RECT 901.000000 309.850000 906.000000 310.150000 ;
        RECT 901.000000 313.850000 906.000000 314.150000 ;
        RECT 901.000000 317.850000 906.000000 318.150000 ;
        RECT 901.000000 325.850000 906.000000 326.150000 ;
        RECT 901.000000 329.850000 906.000000 330.150000 ;
        RECT 901.000000 333.850000 906.000000 334.150000 ;
        RECT 901.000000 337.850000 906.000000 338.150000 ;
        RECT 901.000000 341.850000 906.000000 342.150000 ;
        RECT 951.000000 313.850000 956.000000 314.150000 ;
        RECT 951.000000 309.850000 956.000000 310.150000 ;
        RECT 951.000000 317.850000 956.000000 318.150000 ;
        RECT 951.000000 321.850000 956.000000 322.150000 ;
        RECT 951.000000 325.850000 956.000000 326.150000 ;
        RECT 951.000000 329.850000 956.000000 330.150000 ;
        RECT 951.000000 333.850000 956.000000 334.150000 ;
        RECT 951.000000 337.850000 956.000000 338.150000 ;
        RECT 951.000000 341.850000 956.000000 342.150000 ;
        RECT 1001.000000 305.850000 1006.000000 306.150000 ;
        RECT 1001.000000 277.850000 1006.000000 278.150000 ;
        RECT 1001.000000 269.850000 1006.000000 270.150000 ;
        RECT 1001.000000 273.850000 1006.000000 274.150000 ;
        RECT 1001.000000 285.850000 1006.000000 286.150000 ;
        RECT 1001.000000 281.850000 1006.000000 282.150000 ;
        RECT 1001.000000 289.850000 1006.000000 290.150000 ;
        RECT 1001.000000 293.850000 1006.000000 294.150000 ;
        RECT 1001.000000 301.850000 1006.000000 302.150000 ;
        RECT 1001.000000 297.850000 1006.000000 298.150000 ;
        RECT 1001.000000 313.850000 1006.000000 314.150000 ;
        RECT 1001.000000 309.850000 1006.000000 310.150000 ;
        RECT 1001.000000 317.850000 1006.000000 318.150000 ;
        RECT 1001.000000 321.850000 1006.000000 322.150000 ;
        RECT 1001.000000 329.850000 1006.000000 330.150000 ;
        RECT 1001.000000 325.850000 1006.000000 326.150000 ;
        RECT 1001.000000 333.850000 1006.000000 334.150000 ;
        RECT 1001.000000 337.850000 1006.000000 338.150000 ;
        RECT 1001.000000 341.850000 1006.000000 342.150000 ;
        RECT 1051.000000 261.850000 1056.000000 262.150000 ;
        RECT 1051.000000 265.850000 1056.000000 266.150000 ;
        RECT 1101.000000 265.850000 1106.000000 266.150000 ;
        RECT 1101.000000 261.850000 1106.000000 262.150000 ;
        RECT 1172.000000 197.850000 1182.000000 198.150000 ;
        RECT 1172.000000 201.850000 1182.000000 202.150000 ;
        RECT 1172.000000 205.850000 1182.000000 206.150000 ;
        RECT 1172.000000 209.850000 1182.000000 210.150000 ;
        RECT 1172.000000 221.850000 1182.000000 222.150000 ;
        RECT 1172.000000 217.850000 1182.000000 218.150000 ;
        RECT 1172.000000 213.850000 1182.000000 214.150000 ;
        RECT 1172.000000 225.850000 1182.000000 226.150000 ;
        RECT 1172.000000 229.850000 1182.000000 230.150000 ;
        RECT 1172.000000 233.850000 1182.000000 234.150000 ;
        RECT 1172.000000 237.850000 1182.000000 238.150000 ;
        RECT 1172.000000 241.850000 1182.000000 242.150000 ;
        RECT 1172.000000 245.850000 1182.000000 246.150000 ;
        RECT 1172.000000 249.850000 1182.000000 250.150000 ;
        RECT 1151.000000 257.850000 1156.000000 258.150000 ;
        RECT 1151.000000 265.850000 1156.000000 266.150000 ;
        RECT 1151.000000 261.850000 1156.000000 262.150000 ;
        RECT 1172.000000 265.850000 1182.000000 266.150000 ;
        RECT 1172.000000 253.850000 1182.000000 254.150000 ;
        RECT 1172.000000 257.850000 1182.000000 258.150000 ;
        RECT 1172.000000 261.850000 1182.000000 262.150000 ;
        RECT 1101.000000 305.850000 1106.000000 306.150000 ;
        RECT 1051.000000 305.850000 1056.000000 306.150000 ;
        RECT 1051.000000 285.850000 1056.000000 286.150000 ;
        RECT 1051.000000 281.850000 1056.000000 282.150000 ;
        RECT 1051.000000 273.850000 1056.000000 274.150000 ;
        RECT 1051.000000 269.850000 1056.000000 270.150000 ;
        RECT 1051.000000 277.850000 1056.000000 278.150000 ;
        RECT 1051.000000 289.850000 1056.000000 290.150000 ;
        RECT 1051.000000 293.850000 1056.000000 294.150000 ;
        RECT 1051.000000 297.850000 1056.000000 298.150000 ;
        RECT 1051.000000 301.850000 1056.000000 302.150000 ;
        RECT 1101.000000 269.850000 1106.000000 270.150000 ;
        RECT 1101.000000 273.850000 1106.000000 274.150000 ;
        RECT 1101.000000 277.850000 1106.000000 278.150000 ;
        RECT 1101.000000 281.850000 1106.000000 282.150000 ;
        RECT 1101.000000 285.850000 1106.000000 286.150000 ;
        RECT 1101.000000 301.850000 1106.000000 302.150000 ;
        RECT 1101.000000 297.850000 1106.000000 298.150000 ;
        RECT 1101.000000 293.850000 1106.000000 294.150000 ;
        RECT 1101.000000 289.850000 1106.000000 290.150000 ;
        RECT 1051.000000 321.850000 1056.000000 322.150000 ;
        RECT 1051.000000 309.850000 1056.000000 310.150000 ;
        RECT 1051.000000 313.850000 1056.000000 314.150000 ;
        RECT 1051.000000 317.850000 1056.000000 318.150000 ;
        RECT 1051.000000 325.850000 1056.000000 326.150000 ;
        RECT 1051.000000 329.850000 1056.000000 330.150000 ;
        RECT 1051.000000 333.850000 1056.000000 334.150000 ;
        RECT 1051.000000 337.850000 1056.000000 338.150000 ;
        RECT 1051.000000 341.850000 1056.000000 342.150000 ;
        RECT 1101.000000 313.850000 1106.000000 314.150000 ;
        RECT 1101.000000 309.850000 1106.000000 310.150000 ;
        RECT 1101.000000 317.850000 1106.000000 318.150000 ;
        RECT 1101.000000 321.850000 1106.000000 322.150000 ;
        RECT 1101.000000 325.850000 1106.000000 326.150000 ;
        RECT 1101.000000 329.850000 1106.000000 330.150000 ;
        RECT 1101.000000 333.850000 1106.000000 334.150000 ;
        RECT 1101.000000 337.850000 1106.000000 338.150000 ;
        RECT 1101.000000 341.850000 1106.000000 342.150000 ;
        RECT 1151.000000 305.850000 1156.000000 306.150000 ;
        RECT 1172.000000 305.850000 1182.000000 306.150000 ;
        RECT 1151.000000 277.850000 1156.000000 278.150000 ;
        RECT 1151.000000 269.850000 1156.000000 270.150000 ;
        RECT 1151.000000 273.850000 1156.000000 274.150000 ;
        RECT 1151.000000 281.850000 1156.000000 282.150000 ;
        RECT 1151.000000 285.850000 1156.000000 286.150000 ;
        RECT 1172.000000 277.850000 1182.000000 278.150000 ;
        RECT 1172.000000 269.850000 1182.000000 270.150000 ;
        RECT 1172.000000 273.850000 1182.000000 274.150000 ;
        RECT 1172.000000 281.850000 1182.000000 282.150000 ;
        RECT 1172.000000 285.850000 1182.000000 286.150000 ;
        RECT 1151.000000 301.850000 1156.000000 302.150000 ;
        RECT 1151.000000 297.850000 1156.000000 298.150000 ;
        RECT 1151.000000 289.850000 1156.000000 290.150000 ;
        RECT 1151.000000 293.850000 1156.000000 294.150000 ;
        RECT 1172.000000 301.850000 1182.000000 302.150000 ;
        RECT 1172.000000 289.850000 1182.000000 290.150000 ;
        RECT 1172.000000 293.850000 1182.000000 294.150000 ;
        RECT 1172.000000 297.850000 1182.000000 298.150000 ;
        RECT 1151.000000 321.850000 1156.000000 322.150000 ;
        RECT 1151.000000 317.850000 1156.000000 318.150000 ;
        RECT 1151.000000 309.850000 1156.000000 310.150000 ;
        RECT 1151.000000 313.850000 1156.000000 314.150000 ;
        RECT 1172.000000 321.850000 1182.000000 322.150000 ;
        RECT 1172.000000 309.850000 1182.000000 310.150000 ;
        RECT 1172.000000 313.850000 1182.000000 314.150000 ;
        RECT 1172.000000 317.850000 1182.000000 318.150000 ;
        RECT 1151.000000 329.850000 1156.000000 330.150000 ;
        RECT 1151.000000 325.850000 1156.000000 326.150000 ;
        RECT 1151.000000 333.850000 1156.000000 334.150000 ;
        RECT 1151.000000 337.850000 1156.000000 338.150000 ;
        RECT 1151.000000 341.850000 1156.000000 342.150000 ;
        RECT 1172.000000 329.850000 1182.000000 330.150000 ;
        RECT 1172.000000 325.850000 1182.000000 326.150000 ;
        RECT 1172.000000 333.850000 1182.000000 334.150000 ;
        RECT 1172.000000 337.850000 1182.000000 338.150000 ;
        RECT 1172.000000 341.850000 1182.000000 342.150000 ;
        RECT 4.000000 357.850000 14.000000 358.150000 ;
        RECT 4.000000 353.850000 14.000000 354.150000 ;
        RECT 4.000000 345.850000 14.000000 346.150000 ;
        RECT 4.000000 349.850000 14.000000 350.150000 ;
        RECT 4.000000 369.850000 14.000000 370.150000 ;
        RECT 4.000000 365.850000 14.000000 366.150000 ;
        RECT 4.000000 361.850000 14.000000 362.150000 ;
        RECT 4.000000 377.850000 14.000000 378.150000 ;
        RECT 4.000000 373.850000 14.000000 374.150000 ;
        RECT 51.000000 345.850000 56.000000 346.150000 ;
        RECT 51.000000 369.850000 56.000000 370.150000 ;
        RECT 51.000000 365.850000 56.000000 366.150000 ;
        RECT 51.000000 361.850000 56.000000 362.150000 ;
        RECT 51.000000 373.850000 56.000000 374.150000 ;
        RECT 51.000000 377.850000 56.000000 378.150000 ;
        RECT 4.000000 393.850000 14.000000 394.150000 ;
        RECT 4.000000 389.850000 14.000000 390.150000 ;
        RECT 4.000000 381.850000 14.000000 382.150000 ;
        RECT 4.000000 385.850000 14.000000 386.150000 ;
        RECT 4.000000 397.850000 14.000000 398.150000 ;
        RECT 4.000000 401.850000 14.000000 402.150000 ;
        RECT 4.000000 405.850000 14.000000 406.150000 ;
        RECT 4.000000 409.850000 14.000000 410.150000 ;
        RECT 4.000000 413.850000 14.000000 414.150000 ;
        RECT 51.000000 397.850000 56.000000 398.150000 ;
        RECT 51.000000 385.850000 56.000000 386.150000 ;
        RECT 51.000000 381.850000 56.000000 382.150000 ;
        RECT 51.000000 389.850000 56.000000 390.150000 ;
        RECT 51.000000 393.850000 56.000000 394.150000 ;
        RECT 51.000000 413.850000 56.000000 414.150000 ;
        RECT 51.000000 409.850000 56.000000 410.150000 ;
        RECT 51.000000 405.850000 56.000000 406.150000 ;
        RECT 51.000000 401.850000 56.000000 402.150000 ;
        RECT 101.000000 345.850000 106.000000 346.150000 ;
        RECT 101.000000 349.850000 106.000000 350.150000 ;
        RECT 101.000000 353.850000 106.000000 354.150000 ;
        RECT 101.000000 357.850000 106.000000 358.150000 ;
        RECT 101.000000 361.850000 106.000000 362.150000 ;
        RECT 101.000000 365.850000 106.000000 366.150000 ;
        RECT 101.000000 369.850000 106.000000 370.150000 ;
        RECT 101.000000 373.850000 106.000000 374.150000 ;
        RECT 101.000000 377.850000 106.000000 378.150000 ;
        RECT 101.000000 397.850000 106.000000 398.150000 ;
        RECT 101.000000 381.850000 106.000000 382.150000 ;
        RECT 101.000000 385.850000 106.000000 386.150000 ;
        RECT 101.000000 389.850000 106.000000 390.150000 ;
        RECT 101.000000 393.850000 106.000000 394.150000 ;
        RECT 101.000000 413.850000 106.000000 414.150000 ;
        RECT 101.000000 409.850000 106.000000 410.150000 ;
        RECT 101.000000 405.850000 106.000000 406.150000 ;
        RECT 101.000000 401.850000 106.000000 402.150000 ;
        RECT 4.000000 433.850000 14.000000 434.150000 ;
        RECT 4.000000 429.850000 14.000000 430.150000 ;
        RECT 4.000000 421.850000 14.000000 422.150000 ;
        RECT 4.000000 417.850000 14.000000 418.150000 ;
        RECT 4.000000 425.850000 14.000000 426.150000 ;
        RECT 4.000000 437.850000 14.000000 438.150000 ;
        RECT 4.000000 441.850000 14.000000 442.150000 ;
        RECT 4.000000 445.850000 14.000000 446.150000 ;
        RECT 4.000000 449.850000 14.000000 450.150000 ;
        RECT 4.000000 453.850000 14.000000 454.150000 ;
        RECT 51.000000 417.850000 56.000000 418.150000 ;
        RECT 51.000000 421.850000 56.000000 422.150000 ;
        RECT 51.000000 425.850000 56.000000 426.150000 ;
        RECT 51.000000 429.850000 56.000000 430.150000 ;
        RECT 51.000000 433.850000 56.000000 434.150000 ;
        RECT 51.000000 453.850000 56.000000 454.150000 ;
        RECT 51.000000 449.850000 56.000000 450.150000 ;
        RECT 51.000000 445.850000 56.000000 446.150000 ;
        RECT 51.000000 441.850000 56.000000 442.150000 ;
        RECT 51.000000 437.850000 56.000000 438.150000 ;
        RECT 4.000000 469.850000 14.000000 470.150000 ;
        RECT 4.000000 465.850000 14.000000 466.150000 ;
        RECT 4.000000 457.850000 14.000000 458.150000 ;
        RECT 4.000000 461.850000 14.000000 462.150000 ;
        RECT 4.000000 473.850000 14.000000 474.150000 ;
        RECT 4.000000 477.850000 14.000000 478.150000 ;
        RECT 4.000000 481.850000 14.000000 482.150000 ;
        RECT 4.000000 485.850000 14.000000 486.150000 ;
        RECT 4.000000 489.850000 14.000000 490.150000 ;
        RECT 51.000000 461.850000 56.000000 462.150000 ;
        RECT 51.000000 457.850000 56.000000 458.150000 ;
        RECT 51.000000 465.850000 56.000000 466.150000 ;
        RECT 51.000000 469.850000 56.000000 470.150000 ;
        RECT 51.000000 489.850000 56.000000 490.150000 ;
        RECT 51.000000 485.850000 56.000000 486.150000 ;
        RECT 51.000000 481.850000 56.000000 482.150000 ;
        RECT 51.000000 477.850000 56.000000 478.150000 ;
        RECT 51.000000 473.850000 56.000000 474.150000 ;
        RECT 101.000000 433.850000 106.000000 434.150000 ;
        RECT 101.000000 417.850000 106.000000 418.150000 ;
        RECT 101.000000 421.850000 106.000000 422.150000 ;
        RECT 101.000000 425.850000 106.000000 426.150000 ;
        RECT 101.000000 429.850000 106.000000 430.150000 ;
        RECT 101.000000 437.850000 106.000000 438.150000 ;
        RECT 101.000000 441.850000 106.000000 442.150000 ;
        RECT 101.000000 445.850000 106.000000 446.150000 ;
        RECT 101.000000 449.850000 106.000000 450.150000 ;
        RECT 101.000000 453.850000 106.000000 454.150000 ;
        RECT 101.000000 469.850000 106.000000 470.150000 ;
        RECT 101.000000 465.850000 106.000000 466.150000 ;
        RECT 101.000000 461.850000 106.000000 462.150000 ;
        RECT 101.000000 457.850000 106.000000 458.150000 ;
        RECT 101.000000 473.850000 106.000000 474.150000 ;
        RECT 101.000000 477.850000 106.000000 478.150000 ;
        RECT 101.000000 481.850000 106.000000 482.150000 ;
        RECT 101.000000 485.850000 106.000000 486.150000 ;
        RECT 101.000000 489.850000 106.000000 490.150000 ;
        RECT 151.000000 349.850000 156.000000 350.150000 ;
        RECT 151.000000 345.850000 156.000000 346.150000 ;
        RECT 151.000000 353.850000 156.000000 354.150000 ;
        RECT 151.000000 357.850000 156.000000 358.150000 ;
        RECT 151.000000 361.850000 156.000000 362.150000 ;
        RECT 151.000000 365.850000 156.000000 366.150000 ;
        RECT 151.000000 369.850000 156.000000 370.150000 ;
        RECT 151.000000 377.850000 156.000000 378.150000 ;
        RECT 151.000000 373.850000 156.000000 374.150000 ;
        RECT 201.000000 349.850000 206.000000 350.150000 ;
        RECT 201.000000 345.850000 206.000000 346.150000 ;
        RECT 201.000000 353.850000 206.000000 354.150000 ;
        RECT 201.000000 357.850000 206.000000 358.150000 ;
        RECT 201.000000 361.850000 206.000000 362.150000 ;
        RECT 201.000000 365.850000 206.000000 366.150000 ;
        RECT 201.000000 369.850000 206.000000 370.150000 ;
        RECT 201.000000 373.850000 206.000000 374.150000 ;
        RECT 201.000000 377.850000 206.000000 378.150000 ;
        RECT 151.000000 385.850000 156.000000 386.150000 ;
        RECT 151.000000 381.850000 156.000000 382.150000 ;
        RECT 151.000000 393.850000 156.000000 394.150000 ;
        RECT 151.000000 389.850000 156.000000 390.150000 ;
        RECT 151.000000 397.850000 156.000000 398.150000 ;
        RECT 151.000000 401.850000 156.000000 402.150000 ;
        RECT 201.000000 381.850000 206.000000 382.150000 ;
        RECT 201.000000 385.850000 206.000000 386.150000 ;
        RECT 201.000000 397.850000 206.000000 398.150000 ;
        RECT 201.000000 393.850000 206.000000 394.150000 ;
        RECT 201.000000 389.850000 206.000000 390.150000 ;
        RECT 201.000000 413.850000 206.000000 414.150000 ;
        RECT 201.000000 409.850000 206.000000 410.150000 ;
        RECT 201.000000 405.850000 206.000000 406.150000 ;
        RECT 201.000000 401.850000 206.000000 402.150000 ;
        RECT 251.000000 345.850000 256.000000 346.150000 ;
        RECT 251.000000 349.850000 256.000000 350.150000 ;
        RECT 251.000000 353.850000 256.000000 354.150000 ;
        RECT 251.000000 357.850000 256.000000 358.150000 ;
        RECT 251.000000 369.850000 256.000000 370.150000 ;
        RECT 251.000000 365.850000 256.000000 366.150000 ;
        RECT 251.000000 361.850000 256.000000 362.150000 ;
        RECT 251.000000 373.850000 256.000000 374.150000 ;
        RECT 251.000000 377.850000 256.000000 378.150000 ;
        RECT 251.000000 381.850000 256.000000 382.150000 ;
        RECT 251.000000 385.850000 256.000000 386.150000 ;
        RECT 251.000000 397.850000 256.000000 398.150000 ;
        RECT 251.000000 393.850000 256.000000 394.150000 ;
        RECT 251.000000 389.850000 256.000000 390.150000 ;
        RECT 251.000000 401.850000 256.000000 402.150000 ;
        RECT 151.000000 453.850000 156.000000 454.150000 ;
        RECT 201.000000 429.850000 206.000000 430.150000 ;
        RECT 201.000000 425.850000 206.000000 426.150000 ;
        RECT 201.000000 421.850000 206.000000 422.150000 ;
        RECT 201.000000 417.850000 206.000000 418.150000 ;
        RECT 201.000000 433.850000 206.000000 434.150000 ;
        RECT 201.000000 453.850000 206.000000 454.150000 ;
        RECT 201.000000 449.850000 206.000000 450.150000 ;
        RECT 201.000000 445.850000 206.000000 446.150000 ;
        RECT 201.000000 441.850000 206.000000 442.150000 ;
        RECT 201.000000 437.850000 206.000000 438.150000 ;
        RECT 151.000000 461.850000 156.000000 462.150000 ;
        RECT 151.000000 457.850000 156.000000 458.150000 ;
        RECT 151.000000 469.850000 156.000000 470.150000 ;
        RECT 151.000000 465.850000 156.000000 466.150000 ;
        RECT 151.000000 481.850000 156.000000 482.150000 ;
        RECT 151.000000 477.850000 156.000000 478.150000 ;
        RECT 151.000000 473.850000 156.000000 474.150000 ;
        RECT 151.000000 489.850000 156.000000 490.150000 ;
        RECT 151.000000 485.850000 156.000000 486.150000 ;
        RECT 201.000000 461.850000 206.000000 462.150000 ;
        RECT 201.000000 457.850000 206.000000 458.150000 ;
        RECT 201.000000 465.850000 206.000000 466.150000 ;
        RECT 201.000000 469.850000 206.000000 470.150000 ;
        RECT 201.000000 489.850000 206.000000 490.150000 ;
        RECT 201.000000 485.850000 206.000000 486.150000 ;
        RECT 201.000000 481.850000 206.000000 482.150000 ;
        RECT 201.000000 477.850000 206.000000 478.150000 ;
        RECT 201.000000 473.850000 206.000000 474.150000 ;
        RECT 251.000000 453.850000 256.000000 454.150000 ;
        RECT 251.000000 457.850000 256.000000 458.150000 ;
        RECT 251.000000 461.850000 256.000000 462.150000 ;
        RECT 251.000000 465.850000 256.000000 466.150000 ;
        RECT 251.000000 469.850000 256.000000 470.150000 ;
        RECT 251.000000 481.850000 256.000000 482.150000 ;
        RECT 251.000000 473.850000 256.000000 474.150000 ;
        RECT 251.000000 477.850000 256.000000 478.150000 ;
        RECT 251.000000 485.850000 256.000000 486.150000 ;
        RECT 251.000000 489.850000 256.000000 490.150000 ;
        RECT 4.000000 505.850000 14.000000 506.150000 ;
        RECT 4.000000 501.850000 14.000000 502.150000 ;
        RECT 4.000000 497.850000 14.000000 498.150000 ;
        RECT 4.000000 493.850000 14.000000 494.150000 ;
        RECT 4.000000 513.850000 14.000000 514.150000 ;
        RECT 4.000000 509.850000 14.000000 510.150000 ;
        RECT 51.000000 493.850000 56.000000 494.150000 ;
        RECT 51.000000 497.850000 56.000000 498.150000 ;
        RECT 51.000000 501.850000 56.000000 502.150000 ;
        RECT 51.000000 505.850000 56.000000 506.150000 ;
        RECT 51.000000 513.850000 56.000000 514.150000 ;
        RECT 51.000000 509.850000 56.000000 510.150000 ;
        RECT 101.000000 505.850000 106.000000 506.150000 ;
        RECT 101.000000 501.850000 106.000000 502.150000 ;
        RECT 101.000000 497.850000 106.000000 498.150000 ;
        RECT 101.000000 493.850000 106.000000 494.150000 ;
        RECT 101.000000 513.850000 106.000000 514.150000 ;
        RECT 101.000000 509.850000 106.000000 510.150000 ;
        RECT 151.000000 493.850000 156.000000 494.150000 ;
        RECT 151.000000 497.850000 156.000000 498.150000 ;
        RECT 151.000000 501.850000 156.000000 502.150000 ;
        RECT 151.000000 505.850000 156.000000 506.150000 ;
        RECT 151.000000 513.850000 156.000000 514.150000 ;
        RECT 151.000000 509.850000 156.000000 510.150000 ;
        RECT 201.000000 497.850000 206.000000 498.150000 ;
        RECT 201.000000 493.850000 206.000000 494.150000 ;
        RECT 201.000000 501.850000 206.000000 502.150000 ;
        RECT 201.000000 505.850000 206.000000 506.150000 ;
        RECT 201.000000 513.850000 206.000000 514.150000 ;
        RECT 201.000000 509.850000 206.000000 510.150000 ;
        RECT 251.000000 493.850000 256.000000 494.150000 ;
        RECT 251.000000 497.850000 256.000000 498.150000 ;
        RECT 251.000000 505.850000 256.000000 506.150000 ;
        RECT 251.000000 501.850000 256.000000 502.150000 ;
        RECT 251.000000 513.850000 256.000000 514.150000 ;
        RECT 251.000000 509.850000 256.000000 510.150000 ;
        RECT 301.000000 345.850000 306.000000 346.150000 ;
        RECT 301.000000 349.850000 306.000000 350.150000 ;
        RECT 301.000000 353.850000 306.000000 354.150000 ;
        RECT 301.000000 357.850000 306.000000 358.150000 ;
        RECT 301.000000 369.850000 306.000000 370.150000 ;
        RECT 301.000000 365.850000 306.000000 366.150000 ;
        RECT 301.000000 361.850000 306.000000 362.150000 ;
        RECT 301.000000 377.850000 306.000000 378.150000 ;
        RECT 301.000000 373.850000 306.000000 374.150000 ;
        RECT 351.000000 349.850000 356.000000 350.150000 ;
        RECT 351.000000 345.850000 356.000000 346.150000 ;
        RECT 351.000000 353.850000 356.000000 354.150000 ;
        RECT 351.000000 357.850000 356.000000 358.150000 ;
        RECT 351.000000 361.850000 356.000000 362.150000 ;
        RECT 351.000000 365.850000 356.000000 366.150000 ;
        RECT 351.000000 369.850000 356.000000 370.150000 ;
        RECT 351.000000 373.850000 356.000000 374.150000 ;
        RECT 351.000000 377.850000 356.000000 378.150000 ;
        RECT 301.000000 385.850000 306.000000 386.150000 ;
        RECT 301.000000 381.850000 306.000000 382.150000 ;
        RECT 301.000000 397.850000 306.000000 398.150000 ;
        RECT 301.000000 389.850000 306.000000 390.150000 ;
        RECT 301.000000 393.850000 306.000000 394.150000 ;
        RECT 301.000000 405.850000 306.000000 406.150000 ;
        RECT 301.000000 401.850000 306.000000 402.150000 ;
        RECT 301.000000 409.850000 306.000000 410.150000 ;
        RECT 301.000000 413.850000 306.000000 414.150000 ;
        RECT 351.000000 381.850000 356.000000 382.150000 ;
        RECT 351.000000 385.850000 356.000000 386.150000 ;
        RECT 351.000000 393.850000 356.000000 394.150000 ;
        RECT 351.000000 389.850000 356.000000 390.150000 ;
        RECT 351.000000 397.850000 356.000000 398.150000 ;
        RECT 351.000000 413.850000 356.000000 414.150000 ;
        RECT 351.000000 409.850000 356.000000 410.150000 ;
        RECT 351.000000 405.850000 356.000000 406.150000 ;
        RECT 351.000000 401.850000 356.000000 402.150000 ;
        RECT 401.000000 345.850000 406.000000 346.150000 ;
        RECT 401.000000 349.850000 406.000000 350.150000 ;
        RECT 401.000000 353.850000 406.000000 354.150000 ;
        RECT 401.000000 357.850000 406.000000 358.150000 ;
        RECT 401.000000 365.850000 406.000000 366.150000 ;
        RECT 401.000000 361.850000 406.000000 362.150000 ;
        RECT 401.000000 369.850000 406.000000 370.150000 ;
        RECT 401.000000 373.850000 406.000000 374.150000 ;
        RECT 401.000000 377.850000 406.000000 378.150000 ;
        RECT 401.000000 381.850000 406.000000 382.150000 ;
        RECT 401.000000 385.850000 406.000000 386.150000 ;
        RECT 401.000000 393.850000 406.000000 394.150000 ;
        RECT 401.000000 389.850000 406.000000 390.150000 ;
        RECT 401.000000 397.850000 406.000000 398.150000 ;
        RECT 401.000000 401.850000 406.000000 402.150000 ;
        RECT 401.000000 405.850000 406.000000 406.150000 ;
        RECT 401.000000 409.850000 406.000000 410.150000 ;
        RECT 401.000000 413.850000 406.000000 414.150000 ;
        RECT 301.000000 425.850000 306.000000 426.150000 ;
        RECT 301.000000 417.850000 306.000000 418.150000 ;
        RECT 301.000000 421.850000 306.000000 422.150000 ;
        RECT 301.000000 429.850000 306.000000 430.150000 ;
        RECT 301.000000 433.850000 306.000000 434.150000 ;
        RECT 301.000000 441.850000 306.000000 442.150000 ;
        RECT 301.000000 437.850000 306.000000 438.150000 ;
        RECT 301.000000 453.850000 306.000000 454.150000 ;
        RECT 301.000000 449.850000 306.000000 450.150000 ;
        RECT 301.000000 445.850000 306.000000 446.150000 ;
        RECT 351.000000 425.850000 356.000000 426.150000 ;
        RECT 351.000000 421.850000 356.000000 422.150000 ;
        RECT 351.000000 417.850000 356.000000 418.150000 ;
        RECT 351.000000 433.850000 356.000000 434.150000 ;
        RECT 351.000000 429.850000 356.000000 430.150000 ;
        RECT 351.000000 453.850000 356.000000 454.150000 ;
        RECT 351.000000 449.850000 356.000000 450.150000 ;
        RECT 351.000000 445.850000 356.000000 446.150000 ;
        RECT 351.000000 441.850000 356.000000 442.150000 ;
        RECT 351.000000 437.850000 356.000000 438.150000 ;
        RECT 301.000000 457.850000 306.000000 458.150000 ;
        RECT 301.000000 461.850000 306.000000 462.150000 ;
        RECT 301.000000 465.850000 306.000000 466.150000 ;
        RECT 301.000000 469.850000 306.000000 470.150000 ;
        RECT 301.000000 481.850000 306.000000 482.150000 ;
        RECT 301.000000 477.850000 306.000000 478.150000 ;
        RECT 301.000000 473.850000 306.000000 474.150000 ;
        RECT 301.000000 489.850000 306.000000 490.150000 ;
        RECT 301.000000 485.850000 306.000000 486.150000 ;
        RECT 351.000000 461.850000 356.000000 462.150000 ;
        RECT 351.000000 457.850000 356.000000 458.150000 ;
        RECT 351.000000 465.850000 356.000000 466.150000 ;
        RECT 351.000000 469.850000 356.000000 470.150000 ;
        RECT 351.000000 481.850000 356.000000 482.150000 ;
        RECT 351.000000 473.850000 356.000000 474.150000 ;
        RECT 351.000000 477.850000 356.000000 478.150000 ;
        RECT 351.000000 485.850000 356.000000 486.150000 ;
        RECT 351.000000 489.850000 356.000000 490.150000 ;
        RECT 401.000000 417.850000 406.000000 418.150000 ;
        RECT 401.000000 421.850000 406.000000 422.150000 ;
        RECT 401.000000 425.850000 406.000000 426.150000 ;
        RECT 401.000000 433.850000 406.000000 434.150000 ;
        RECT 401.000000 429.850000 406.000000 430.150000 ;
        RECT 401.000000 441.850000 406.000000 442.150000 ;
        RECT 401.000000 437.850000 406.000000 438.150000 ;
        RECT 401.000000 445.850000 406.000000 446.150000 ;
        RECT 401.000000 453.850000 406.000000 454.150000 ;
        RECT 401.000000 449.850000 406.000000 450.150000 ;
        RECT 401.000000 457.850000 406.000000 458.150000 ;
        RECT 401.000000 461.850000 406.000000 462.150000 ;
        RECT 401.000000 465.850000 406.000000 466.150000 ;
        RECT 401.000000 469.850000 406.000000 470.150000 ;
        RECT 401.000000 481.850000 406.000000 482.150000 ;
        RECT 401.000000 473.850000 406.000000 474.150000 ;
        RECT 401.000000 477.850000 406.000000 478.150000 ;
        RECT 401.000000 485.850000 406.000000 486.150000 ;
        RECT 401.000000 489.850000 406.000000 490.150000 ;
        RECT 451.000000 345.850000 456.000000 346.150000 ;
        RECT 451.000000 369.850000 456.000000 370.150000 ;
        RECT 451.000000 373.850000 456.000000 374.150000 ;
        RECT 451.000000 377.850000 456.000000 378.150000 ;
        RECT 501.000000 345.850000 506.000000 346.150000 ;
        RECT 501.000000 349.850000 506.000000 350.150000 ;
        RECT 501.000000 353.850000 506.000000 354.150000 ;
        RECT 501.000000 357.850000 506.000000 358.150000 ;
        RECT 501.000000 365.850000 506.000000 366.150000 ;
        RECT 501.000000 361.850000 506.000000 362.150000 ;
        RECT 501.000000 369.850000 506.000000 370.150000 ;
        RECT 501.000000 377.850000 506.000000 378.150000 ;
        RECT 501.000000 373.850000 506.000000 374.150000 ;
        RECT 451.000000 381.850000 456.000000 382.150000 ;
        RECT 451.000000 385.850000 456.000000 386.150000 ;
        RECT 451.000000 397.850000 456.000000 398.150000 ;
        RECT 451.000000 393.850000 456.000000 394.150000 ;
        RECT 451.000000 389.850000 456.000000 390.150000 ;
        RECT 501.000000 385.850000 506.000000 386.150000 ;
        RECT 501.000000 381.850000 506.000000 382.150000 ;
        RECT 501.000000 393.850000 506.000000 394.150000 ;
        RECT 501.000000 389.850000 506.000000 390.150000 ;
        RECT 501.000000 397.850000 506.000000 398.150000 ;
        RECT 501.000000 401.850000 506.000000 402.150000 ;
        RECT 501.000000 405.850000 506.000000 406.150000 ;
        RECT 501.000000 409.850000 506.000000 410.150000 ;
        RECT 501.000000 413.850000 506.000000 414.150000 ;
        RECT 551.000000 357.850000 556.000000 358.150000 ;
        RECT 551.000000 353.850000 556.000000 354.150000 ;
        RECT 551.000000 349.850000 556.000000 350.150000 ;
        RECT 551.000000 345.850000 556.000000 346.150000 ;
        RECT 551.000000 361.850000 556.000000 362.150000 ;
        RECT 551.000000 365.850000 556.000000 366.150000 ;
        RECT 551.000000 369.850000 556.000000 370.150000 ;
        RECT 551.000000 373.850000 556.000000 374.150000 ;
        RECT 551.000000 377.850000 556.000000 378.150000 ;
        RECT 551.000000 385.850000 556.000000 386.150000 ;
        RECT 551.000000 381.850000 556.000000 382.150000 ;
        RECT 551.000000 397.850000 556.000000 398.150000 ;
        RECT 551.000000 393.850000 556.000000 394.150000 ;
        RECT 551.000000 389.850000 556.000000 390.150000 ;
        RECT 551.000000 413.850000 556.000000 414.150000 ;
        RECT 551.000000 409.850000 556.000000 410.150000 ;
        RECT 551.000000 405.850000 556.000000 406.150000 ;
        RECT 551.000000 401.850000 556.000000 402.150000 ;
        RECT 451.000000 425.850000 456.000000 426.150000 ;
        RECT 451.000000 421.850000 456.000000 422.150000 ;
        RECT 451.000000 429.850000 456.000000 430.150000 ;
        RECT 451.000000 433.850000 456.000000 434.150000 ;
        RECT 451.000000 441.850000 456.000000 442.150000 ;
        RECT 451.000000 437.850000 456.000000 438.150000 ;
        RECT 451.000000 453.850000 456.000000 454.150000 ;
        RECT 451.000000 449.850000 456.000000 450.150000 ;
        RECT 451.000000 445.850000 456.000000 446.150000 ;
        RECT 501.000000 417.850000 506.000000 418.150000 ;
        RECT 501.000000 421.850000 506.000000 422.150000 ;
        RECT 501.000000 425.850000 506.000000 426.150000 ;
        RECT 501.000000 429.850000 506.000000 430.150000 ;
        RECT 501.000000 433.850000 506.000000 434.150000 ;
        RECT 501.000000 437.850000 506.000000 438.150000 ;
        RECT 501.000000 441.850000 506.000000 442.150000 ;
        RECT 501.000000 445.850000 506.000000 446.150000 ;
        RECT 501.000000 449.850000 506.000000 450.150000 ;
        RECT 501.000000 453.850000 506.000000 454.150000 ;
        RECT 451.000000 461.850000 456.000000 462.150000 ;
        RECT 451.000000 457.850000 456.000000 458.150000 ;
        RECT 451.000000 465.850000 456.000000 466.150000 ;
        RECT 451.000000 469.850000 456.000000 470.150000 ;
        RECT 451.000000 481.850000 456.000000 482.150000 ;
        RECT 451.000000 477.850000 456.000000 478.150000 ;
        RECT 451.000000 473.850000 456.000000 474.150000 ;
        RECT 451.000000 489.850000 456.000000 490.150000 ;
        RECT 451.000000 485.850000 456.000000 486.150000 ;
        RECT 501.000000 457.850000 506.000000 458.150000 ;
        RECT 501.000000 461.850000 506.000000 462.150000 ;
        RECT 501.000000 465.850000 506.000000 466.150000 ;
        RECT 501.000000 469.850000 506.000000 470.150000 ;
        RECT 501.000000 481.850000 506.000000 482.150000 ;
        RECT 501.000000 473.850000 506.000000 474.150000 ;
        RECT 501.000000 477.850000 506.000000 478.150000 ;
        RECT 501.000000 485.850000 506.000000 486.150000 ;
        RECT 501.000000 489.850000 506.000000 490.150000 ;
        RECT 551.000000 429.850000 556.000000 430.150000 ;
        RECT 551.000000 425.850000 556.000000 426.150000 ;
        RECT 551.000000 417.850000 556.000000 418.150000 ;
        RECT 551.000000 421.850000 556.000000 422.150000 ;
        RECT 551.000000 433.850000 556.000000 434.150000 ;
        RECT 551.000000 437.850000 556.000000 438.150000 ;
        RECT 551.000000 441.850000 556.000000 442.150000 ;
        RECT 551.000000 445.850000 556.000000 446.150000 ;
        RECT 551.000000 449.850000 556.000000 450.150000 ;
        RECT 551.000000 453.850000 556.000000 454.150000 ;
        RECT 551.000000 457.850000 556.000000 458.150000 ;
        RECT 551.000000 461.850000 556.000000 462.150000 ;
        RECT 551.000000 465.850000 556.000000 466.150000 ;
        RECT 551.000000 469.850000 556.000000 470.150000 ;
        RECT 551.000000 481.850000 556.000000 482.150000 ;
        RECT 551.000000 473.850000 556.000000 474.150000 ;
        RECT 551.000000 477.850000 556.000000 478.150000 ;
        RECT 551.000000 485.850000 556.000000 486.150000 ;
        RECT 551.000000 489.850000 556.000000 490.150000 ;
        RECT 301.000000 497.850000 306.000000 498.150000 ;
        RECT 301.000000 493.850000 306.000000 494.150000 ;
        RECT 301.000000 501.850000 306.000000 502.150000 ;
        RECT 301.000000 505.850000 306.000000 506.150000 ;
        RECT 301.000000 517.850000 306.000000 518.150000 ;
        RECT 301.000000 513.850000 306.000000 514.150000 ;
        RECT 301.000000 509.850000 306.000000 510.150000 ;
        RECT 351.000000 493.850000 356.000000 494.150000 ;
        RECT 351.000000 497.850000 356.000000 498.150000 ;
        RECT 351.000000 505.850000 356.000000 506.150000 ;
        RECT 351.000000 501.850000 356.000000 502.150000 ;
        RECT 351.000000 509.850000 356.000000 510.150000 ;
        RECT 351.000000 513.850000 356.000000 514.150000 ;
        RECT 351.000000 517.850000 356.000000 518.150000 ;
        RECT 351.000000 521.850000 356.000000 522.150000 ;
        RECT 351.000000 525.850000 356.000000 526.150000 ;
        RECT 351.000000 533.850000 356.000000 534.150000 ;
        RECT 351.000000 529.850000 356.000000 530.150000 ;
        RECT 351.000000 537.850000 356.000000 538.150000 ;
        RECT 351.000000 541.850000 356.000000 542.150000 ;
        RECT 351.000000 545.850000 356.000000 546.150000 ;
        RECT 351.000000 561.850000 356.000000 562.150000 ;
        RECT 351.000000 557.850000 356.000000 558.150000 ;
        RECT 351.000000 553.850000 356.000000 554.150000 ;
        RECT 351.000000 549.850000 356.000000 550.150000 ;
        RECT 375.000000 493.850000 385.000000 494.150000 ;
        RECT 375.000000 497.850000 385.000000 498.150000 ;
        RECT 375.000000 501.850000 385.000000 502.150000 ;
        RECT 375.000000 505.850000 385.000000 506.150000 ;
        RECT 401.000000 493.850000 406.000000 494.150000 ;
        RECT 401.000000 497.850000 406.000000 498.150000 ;
        RECT 401.000000 501.850000 406.000000 502.150000 ;
        RECT 375.000000 509.850000 385.000000 510.150000 ;
        RECT 375.000000 513.850000 385.000000 514.150000 ;
        RECT 375.000000 517.850000 385.000000 518.150000 ;
        RECT 375.000000 521.850000 385.000000 522.150000 ;
        RECT 375.000000 525.850000 385.000000 526.150000 ;
        RECT 375.000000 545.850000 385.000000 546.150000 ;
        RECT 375.000000 541.850000 385.000000 542.150000 ;
        RECT 375.000000 537.850000 385.000000 538.150000 ;
        RECT 375.000000 533.850000 385.000000 534.150000 ;
        RECT 375.000000 529.850000 385.000000 530.150000 ;
        RECT 375.000000 561.850000 385.000000 562.150000 ;
        RECT 375.000000 557.850000 385.000000 558.150000 ;
        RECT 375.000000 553.850000 385.000000 554.150000 ;
        RECT 375.000000 549.850000 385.000000 550.150000 ;
        RECT 351.000000 565.850000 356.000000 566.150000 ;
        RECT 351.000000 569.850000 356.000000 570.150000 ;
        RECT 351.000000 573.850000 356.000000 574.150000 ;
        RECT 351.000000 577.850000 356.000000 578.150000 ;
        RECT 351.000000 581.850000 356.000000 582.150000 ;
        RECT 351.000000 601.850000 356.000000 602.150000 ;
        RECT 351.000000 597.850000 356.000000 598.150000 ;
        RECT 351.000000 593.850000 356.000000 594.150000 ;
        RECT 351.000000 589.850000 356.000000 590.150000 ;
        RECT 351.000000 585.850000 356.000000 586.150000 ;
        RECT 351.000000 609.850000 356.000000 610.150000 ;
        RECT 351.000000 605.850000 356.000000 606.150000 ;
        RECT 351.000000 613.850000 356.000000 614.150000 ;
        RECT 351.000000 617.850000 356.000000 618.150000 ;
        RECT 351.000000 621.850000 356.000000 622.150000 ;
        RECT 351.000000 625.850000 356.000000 626.150000 ;
        RECT 351.000000 629.850000 356.000000 630.150000 ;
        RECT 351.000000 633.850000 356.000000 634.150000 ;
        RECT 351.000000 637.850000 356.000000 638.150000 ;
        RECT 375.000000 565.850000 385.000000 566.150000 ;
        RECT 375.000000 569.850000 385.000000 570.150000 ;
        RECT 375.000000 573.850000 385.000000 574.150000 ;
        RECT 375.000000 577.850000 385.000000 578.150000 ;
        RECT 375.000000 581.850000 385.000000 582.150000 ;
        RECT 375.000000 585.850000 385.000000 586.150000 ;
        RECT 375.000000 589.850000 385.000000 590.150000 ;
        RECT 375.000000 593.850000 385.000000 594.150000 ;
        RECT 375.000000 597.850000 385.000000 598.150000 ;
        RECT 375.000000 601.850000 385.000000 602.150000 ;
        RECT 375.000000 617.850000 385.000000 618.150000 ;
        RECT 375.000000 613.850000 385.000000 614.150000 ;
        RECT 375.000000 609.850000 385.000000 610.150000 ;
        RECT 375.000000 605.850000 385.000000 606.150000 ;
        RECT 375.000000 621.850000 385.000000 622.150000 ;
        RECT 375.000000 625.850000 385.000000 626.150000 ;
        RECT 375.000000 629.850000 385.000000 630.150000 ;
        RECT 375.000000 633.850000 385.000000 634.150000 ;
        RECT 375.000000 637.850000 385.000000 638.150000 ;
        RECT 451.000000 493.850000 456.000000 494.150000 ;
        RECT 451.000000 497.850000 456.000000 498.150000 ;
        RECT 451.000000 501.850000 456.000000 502.150000 ;
        RECT 501.000000 497.850000 506.000000 498.150000 ;
        RECT 501.000000 493.850000 506.000000 494.150000 ;
        RECT 501.000000 501.850000 506.000000 502.150000 ;
        RECT 551.000000 493.850000 556.000000 494.150000 ;
        RECT 551.000000 497.850000 556.000000 498.150000 ;
        RECT 551.000000 501.850000 556.000000 502.150000 ;
        RECT 351.000000 657.850000 356.000000 658.150000 ;
        RECT 351.000000 641.850000 356.000000 642.150000 ;
        RECT 351.000000 645.850000 356.000000 646.150000 ;
        RECT 351.000000 649.850000 356.000000 650.150000 ;
        RECT 351.000000 653.850000 356.000000 654.150000 ;
        RECT 351.000000 673.850000 356.000000 674.150000 ;
        RECT 351.000000 669.850000 356.000000 670.150000 ;
        RECT 351.000000 665.850000 356.000000 666.150000 ;
        RECT 351.000000 661.850000 356.000000 662.150000 ;
        RECT 301.000000 681.850000 306.000000 682.150000 ;
        RECT 301.000000 677.850000 306.000000 678.150000 ;
        RECT 351.000000 677.850000 356.000000 678.150000 ;
        RECT 351.000000 681.850000 356.000000 682.150000 ;
        RECT 375.000000 657.850000 385.000000 658.150000 ;
        RECT 401.000000 657.850000 406.000000 658.150000 ;
        RECT 375.000000 641.850000 385.000000 642.150000 ;
        RECT 375.000000 645.850000 385.000000 646.150000 ;
        RECT 375.000000 649.850000 385.000000 650.150000 ;
        RECT 375.000000 653.850000 385.000000 654.150000 ;
        RECT 375.000000 665.850000 385.000000 666.150000 ;
        RECT 375.000000 661.850000 385.000000 662.150000 ;
        RECT 375.000000 669.850000 385.000000 670.150000 ;
        RECT 375.000000 673.850000 385.000000 674.150000 ;
        RECT 401.000000 665.850000 406.000000 666.150000 ;
        RECT 401.000000 661.850000 406.000000 662.150000 ;
        RECT 401.000000 669.850000 406.000000 670.150000 ;
        RECT 401.000000 673.850000 406.000000 674.150000 ;
        RECT 401.000000 677.850000 406.000000 678.150000 ;
        RECT 375.000000 677.850000 385.000000 678.150000 ;
        RECT 401.000000 681.850000 406.000000 682.150000 ;
        RECT 375.000000 681.850000 385.000000 682.150000 ;
        RECT 451.000000 657.850000 456.000000 658.150000 ;
        RECT 451.000000 673.850000 456.000000 674.150000 ;
        RECT 451.000000 669.850000 456.000000 670.150000 ;
        RECT 451.000000 665.850000 456.000000 666.150000 ;
        RECT 451.000000 661.850000 456.000000 662.150000 ;
        RECT 501.000000 657.850000 506.000000 658.150000 ;
        RECT 501.000000 661.850000 506.000000 662.150000 ;
        RECT 501.000000 665.850000 506.000000 666.150000 ;
        RECT 501.000000 673.850000 506.000000 674.150000 ;
        RECT 501.000000 669.850000 506.000000 670.150000 ;
        RECT 451.000000 677.850000 456.000000 678.150000 ;
        RECT 451.000000 681.850000 456.000000 682.150000 ;
        RECT 501.000000 677.850000 506.000000 678.150000 ;
        RECT 501.000000 681.850000 506.000000 682.150000 ;
        RECT 551.000000 673.850000 556.000000 674.150000 ;
        RECT 551.000000 657.850000 556.000000 658.150000 ;
        RECT 551.000000 661.850000 556.000000 662.150000 ;
        RECT 551.000000 665.850000 556.000000 666.150000 ;
        RECT 551.000000 669.850000 556.000000 670.150000 ;
        RECT 551.000000 681.850000 556.000000 682.150000 ;
        RECT 551.000000 677.850000 556.000000 678.150000 ;
        RECT 601.000000 357.850000 606.000000 358.150000 ;
        RECT 601.000000 353.850000 606.000000 354.150000 ;
        RECT 601.000000 345.850000 606.000000 346.150000 ;
        RECT 601.000000 349.850000 606.000000 350.150000 ;
        RECT 601.000000 361.850000 606.000000 362.150000 ;
        RECT 601.000000 365.850000 606.000000 366.150000 ;
        RECT 601.000000 369.850000 606.000000 370.150000 ;
        RECT 601.000000 373.850000 606.000000 374.150000 ;
        RECT 601.000000 377.850000 606.000000 378.150000 ;
        RECT 651.000000 349.850000 656.000000 350.150000 ;
        RECT 651.000000 345.850000 656.000000 346.150000 ;
        RECT 651.000000 353.850000 656.000000 354.150000 ;
        RECT 651.000000 357.850000 656.000000 358.150000 ;
        RECT 651.000000 361.850000 656.000000 362.150000 ;
        RECT 651.000000 365.850000 656.000000 366.150000 ;
        RECT 651.000000 369.850000 656.000000 370.150000 ;
        RECT 651.000000 377.850000 656.000000 378.150000 ;
        RECT 651.000000 373.850000 656.000000 374.150000 ;
        RECT 601.000000 385.850000 606.000000 386.150000 ;
        RECT 601.000000 381.850000 606.000000 382.150000 ;
        RECT 601.000000 397.850000 606.000000 398.150000 ;
        RECT 601.000000 389.850000 606.000000 390.150000 ;
        RECT 601.000000 393.850000 606.000000 394.150000 ;
        RECT 601.000000 405.850000 606.000000 406.150000 ;
        RECT 601.000000 401.850000 606.000000 402.150000 ;
        RECT 601.000000 413.850000 606.000000 414.150000 ;
        RECT 601.000000 409.850000 606.000000 410.150000 ;
        RECT 651.000000 385.850000 656.000000 386.150000 ;
        RECT 651.000000 381.850000 656.000000 382.150000 ;
        RECT 651.000000 393.850000 656.000000 394.150000 ;
        RECT 651.000000 389.850000 656.000000 390.150000 ;
        RECT 651.000000 397.850000 656.000000 398.150000 ;
        RECT 651.000000 405.850000 656.000000 406.150000 ;
        RECT 651.000000 401.850000 656.000000 402.150000 ;
        RECT 651.000000 409.850000 656.000000 410.150000 ;
        RECT 651.000000 413.850000 656.000000 414.150000 ;
        RECT 701.000000 357.850000 706.000000 358.150000 ;
        RECT 701.000000 353.850000 706.000000 354.150000 ;
        RECT 701.000000 349.850000 706.000000 350.150000 ;
        RECT 701.000000 345.850000 706.000000 346.150000 ;
        RECT 701.000000 361.850000 706.000000 362.150000 ;
        RECT 701.000000 365.850000 706.000000 366.150000 ;
        RECT 701.000000 369.850000 706.000000 370.150000 ;
        RECT 701.000000 373.850000 706.000000 374.150000 ;
        RECT 701.000000 377.850000 706.000000 378.150000 ;
        RECT 701.000000 385.850000 706.000000 386.150000 ;
        RECT 701.000000 381.850000 706.000000 382.150000 ;
        RECT 701.000000 397.850000 706.000000 398.150000 ;
        RECT 701.000000 393.850000 706.000000 394.150000 ;
        RECT 701.000000 389.850000 706.000000 390.150000 ;
        RECT 701.000000 413.850000 706.000000 414.150000 ;
        RECT 701.000000 409.850000 706.000000 410.150000 ;
        RECT 701.000000 405.850000 706.000000 406.150000 ;
        RECT 701.000000 401.850000 706.000000 402.150000 ;
        RECT 601.000000 417.850000 606.000000 418.150000 ;
        RECT 601.000000 421.850000 606.000000 422.150000 ;
        RECT 601.000000 425.850000 606.000000 426.150000 ;
        RECT 601.000000 429.850000 606.000000 430.150000 ;
        RECT 601.000000 433.850000 606.000000 434.150000 ;
        RECT 601.000000 441.850000 606.000000 442.150000 ;
        RECT 601.000000 437.850000 606.000000 438.150000 ;
        RECT 601.000000 453.850000 606.000000 454.150000 ;
        RECT 601.000000 449.850000 606.000000 450.150000 ;
        RECT 601.000000 445.850000 606.000000 446.150000 ;
        RECT 651.000000 417.850000 656.000000 418.150000 ;
        RECT 651.000000 425.850000 656.000000 426.150000 ;
        RECT 651.000000 421.850000 656.000000 422.150000 ;
        RECT 651.000000 429.850000 656.000000 430.150000 ;
        RECT 651.000000 433.850000 656.000000 434.150000 ;
        RECT 651.000000 437.850000 656.000000 438.150000 ;
        RECT 651.000000 441.850000 656.000000 442.150000 ;
        RECT 651.000000 445.850000 656.000000 446.150000 ;
        RECT 651.000000 449.850000 656.000000 450.150000 ;
        RECT 651.000000 453.850000 656.000000 454.150000 ;
        RECT 601.000000 469.850000 606.000000 470.150000 ;
        RECT 601.000000 465.850000 606.000000 466.150000 ;
        RECT 601.000000 457.850000 606.000000 458.150000 ;
        RECT 601.000000 461.850000 606.000000 462.150000 ;
        RECT 601.000000 481.850000 606.000000 482.150000 ;
        RECT 601.000000 477.850000 606.000000 478.150000 ;
        RECT 601.000000 473.850000 606.000000 474.150000 ;
        RECT 601.000000 489.850000 606.000000 490.150000 ;
        RECT 601.000000 485.850000 606.000000 486.150000 ;
        RECT 651.000000 461.850000 656.000000 462.150000 ;
        RECT 651.000000 457.850000 656.000000 458.150000 ;
        RECT 651.000000 469.850000 656.000000 470.150000 ;
        RECT 651.000000 465.850000 656.000000 466.150000 ;
        RECT 651.000000 481.850000 656.000000 482.150000 ;
        RECT 651.000000 477.850000 656.000000 478.150000 ;
        RECT 651.000000 473.850000 656.000000 474.150000 ;
        RECT 651.000000 489.850000 656.000000 490.150000 ;
        RECT 651.000000 485.850000 656.000000 486.150000 ;
        RECT 701.000000 425.850000 706.000000 426.150000 ;
        RECT 701.000000 421.850000 706.000000 422.150000 ;
        RECT 701.000000 417.850000 706.000000 418.150000 ;
        RECT 701.000000 429.850000 706.000000 430.150000 ;
        RECT 701.000000 433.850000 706.000000 434.150000 ;
        RECT 701.000000 437.850000 706.000000 438.150000 ;
        RECT 701.000000 441.850000 706.000000 442.150000 ;
        RECT 701.000000 445.850000 706.000000 446.150000 ;
        RECT 701.000000 449.850000 706.000000 450.150000 ;
        RECT 701.000000 453.850000 706.000000 454.150000 ;
        RECT 725.000000 433.850000 735.000000 434.150000 ;
        RECT 725.000000 437.850000 735.000000 438.150000 ;
        RECT 725.000000 441.850000 735.000000 442.150000 ;
        RECT 725.000000 453.850000 735.000000 454.150000 ;
        RECT 725.000000 449.850000 735.000000 450.150000 ;
        RECT 725.000000 445.850000 735.000000 446.150000 ;
        RECT 701.000000 457.850000 706.000000 458.150000 ;
        RECT 701.000000 461.850000 706.000000 462.150000 ;
        RECT 701.000000 465.850000 706.000000 466.150000 ;
        RECT 701.000000 469.850000 706.000000 470.150000 ;
        RECT 701.000000 481.850000 706.000000 482.150000 ;
        RECT 701.000000 473.850000 706.000000 474.150000 ;
        RECT 701.000000 477.850000 706.000000 478.150000 ;
        RECT 701.000000 485.850000 706.000000 486.150000 ;
        RECT 701.000000 489.850000 706.000000 490.150000 ;
        RECT 725.000000 469.850000 735.000000 470.150000 ;
        RECT 725.000000 465.850000 735.000000 466.150000 ;
        RECT 725.000000 457.850000 735.000000 458.150000 ;
        RECT 725.000000 461.850000 735.000000 462.150000 ;
        RECT 725.000000 481.850000 735.000000 482.150000 ;
        RECT 725.000000 477.850000 735.000000 478.150000 ;
        RECT 725.000000 473.850000 735.000000 474.150000 ;
        RECT 725.000000 489.850000 735.000000 490.150000 ;
        RECT 725.000000 485.850000 735.000000 486.150000 ;
        RECT 751.000000 357.850000 756.000000 358.150000 ;
        RECT 751.000000 353.850000 756.000000 354.150000 ;
        RECT 751.000000 349.850000 756.000000 350.150000 ;
        RECT 751.000000 345.850000 756.000000 346.150000 ;
        RECT 751.000000 361.850000 756.000000 362.150000 ;
        RECT 751.000000 365.850000 756.000000 366.150000 ;
        RECT 751.000000 369.850000 756.000000 370.150000 ;
        RECT 751.000000 373.850000 756.000000 374.150000 ;
        RECT 751.000000 377.850000 756.000000 378.150000 ;
        RECT 801.000000 345.850000 806.000000 346.150000 ;
        RECT 801.000000 349.850000 806.000000 350.150000 ;
        RECT 801.000000 353.850000 806.000000 354.150000 ;
        RECT 801.000000 357.850000 806.000000 358.150000 ;
        RECT 801.000000 361.850000 806.000000 362.150000 ;
        RECT 801.000000 365.850000 806.000000 366.150000 ;
        RECT 801.000000 369.850000 806.000000 370.150000 ;
        RECT 801.000000 377.850000 806.000000 378.150000 ;
        RECT 801.000000 373.850000 806.000000 374.150000 ;
        RECT 751.000000 385.850000 756.000000 386.150000 ;
        RECT 751.000000 381.850000 756.000000 382.150000 ;
        RECT 751.000000 393.850000 756.000000 394.150000 ;
        RECT 751.000000 389.850000 756.000000 390.150000 ;
        RECT 751.000000 397.850000 756.000000 398.150000 ;
        RECT 751.000000 401.850000 756.000000 402.150000 ;
        RECT 751.000000 405.850000 756.000000 406.150000 ;
        RECT 751.000000 409.850000 756.000000 410.150000 ;
        RECT 751.000000 413.850000 756.000000 414.150000 ;
        RECT 801.000000 385.850000 806.000000 386.150000 ;
        RECT 801.000000 381.850000 806.000000 382.150000 ;
        RECT 801.000000 393.850000 806.000000 394.150000 ;
        RECT 801.000000 389.850000 806.000000 390.150000 ;
        RECT 801.000000 397.850000 806.000000 398.150000 ;
        RECT 801.000000 405.850000 806.000000 406.150000 ;
        RECT 801.000000 401.850000 806.000000 402.150000 ;
        RECT 801.000000 409.850000 806.000000 410.150000 ;
        RECT 801.000000 413.850000 806.000000 414.150000 ;
        RECT 851.000000 357.850000 856.000000 358.150000 ;
        RECT 851.000000 353.850000 856.000000 354.150000 ;
        RECT 851.000000 349.850000 856.000000 350.150000 ;
        RECT 851.000000 345.850000 856.000000 346.150000 ;
        RECT 851.000000 361.850000 856.000000 362.150000 ;
        RECT 851.000000 365.850000 856.000000 366.150000 ;
        RECT 851.000000 369.850000 856.000000 370.150000 ;
        RECT 851.000000 373.850000 856.000000 374.150000 ;
        RECT 851.000000 377.850000 856.000000 378.150000 ;
        RECT 851.000000 385.850000 856.000000 386.150000 ;
        RECT 851.000000 381.850000 856.000000 382.150000 ;
        RECT 851.000000 397.850000 856.000000 398.150000 ;
        RECT 851.000000 393.850000 856.000000 394.150000 ;
        RECT 851.000000 389.850000 856.000000 390.150000 ;
        RECT 851.000000 413.850000 856.000000 414.150000 ;
        RECT 851.000000 409.850000 856.000000 410.150000 ;
        RECT 851.000000 405.850000 856.000000 406.150000 ;
        RECT 851.000000 401.850000 856.000000 402.150000 ;
        RECT 751.000000 417.850000 756.000000 418.150000 ;
        RECT 751.000000 421.850000 756.000000 422.150000 ;
        RECT 751.000000 425.850000 756.000000 426.150000 ;
        RECT 751.000000 429.850000 756.000000 430.150000 ;
        RECT 751.000000 433.850000 756.000000 434.150000 ;
        RECT 751.000000 437.850000 756.000000 438.150000 ;
        RECT 751.000000 441.850000 756.000000 442.150000 ;
        RECT 801.000000 417.850000 806.000000 418.150000 ;
        RECT 801.000000 421.850000 806.000000 422.150000 ;
        RECT 801.000000 425.850000 806.000000 426.150000 ;
        RECT 801.000000 429.850000 806.000000 430.150000 ;
        RECT 801.000000 433.850000 806.000000 434.150000 ;
        RECT 801.000000 437.850000 806.000000 438.150000 ;
        RECT 801.000000 441.850000 806.000000 442.150000 ;
        RECT 851.000000 417.850000 856.000000 418.150000 ;
        RECT 851.000000 421.850000 856.000000 422.150000 ;
        RECT 851.000000 425.850000 856.000000 426.150000 ;
        RECT 851.000000 433.850000 856.000000 434.150000 ;
        RECT 851.000000 429.850000 856.000000 430.150000 ;
        RECT 851.000000 441.850000 856.000000 442.150000 ;
        RECT 851.000000 437.850000 856.000000 438.150000 ;
        RECT 601.000000 501.850000 606.000000 502.150000 ;
        RECT 601.000000 497.850000 606.000000 498.150000 ;
        RECT 601.000000 493.850000 606.000000 494.150000 ;
        RECT 651.000000 497.850000 656.000000 498.150000 ;
        RECT 651.000000 493.850000 656.000000 494.150000 ;
        RECT 651.000000 501.850000 656.000000 502.150000 ;
        RECT 701.000000 501.850000 706.000000 502.150000 ;
        RECT 701.000000 493.850000 706.000000 494.150000 ;
        RECT 701.000000 497.850000 706.000000 498.150000 ;
        RECT 725.000000 497.850000 735.000000 498.150000 ;
        RECT 725.000000 493.850000 735.000000 494.150000 ;
        RECT 725.000000 501.850000 735.000000 502.150000 ;
        RECT 901.000000 357.850000 906.000000 358.150000 ;
        RECT 901.000000 353.850000 906.000000 354.150000 ;
        RECT 901.000000 349.850000 906.000000 350.150000 ;
        RECT 901.000000 345.850000 906.000000 346.150000 ;
        RECT 901.000000 361.850000 906.000000 362.150000 ;
        RECT 901.000000 365.850000 906.000000 366.150000 ;
        RECT 901.000000 369.850000 906.000000 370.150000 ;
        RECT 901.000000 373.850000 906.000000 374.150000 ;
        RECT 901.000000 377.850000 906.000000 378.150000 ;
        RECT 951.000000 345.850000 956.000000 346.150000 ;
        RECT 951.000000 349.850000 956.000000 350.150000 ;
        RECT 951.000000 353.850000 956.000000 354.150000 ;
        RECT 951.000000 357.850000 956.000000 358.150000 ;
        RECT 951.000000 361.850000 956.000000 362.150000 ;
        RECT 951.000000 365.850000 956.000000 366.150000 ;
        RECT 951.000000 369.850000 956.000000 370.150000 ;
        RECT 951.000000 373.850000 956.000000 374.150000 ;
        RECT 951.000000 377.850000 956.000000 378.150000 ;
        RECT 901.000000 385.850000 906.000000 386.150000 ;
        RECT 901.000000 381.850000 906.000000 382.150000 ;
        RECT 901.000000 393.850000 906.000000 394.150000 ;
        RECT 901.000000 389.850000 906.000000 390.150000 ;
        RECT 901.000000 397.850000 906.000000 398.150000 ;
        RECT 901.000000 405.850000 906.000000 406.150000 ;
        RECT 901.000000 401.850000 906.000000 402.150000 ;
        RECT 901.000000 409.850000 906.000000 410.150000 ;
        RECT 901.000000 413.850000 906.000000 414.150000 ;
        RECT 951.000000 385.850000 956.000000 386.150000 ;
        RECT 951.000000 381.850000 956.000000 382.150000 ;
        RECT 951.000000 389.850000 956.000000 390.150000 ;
        RECT 951.000000 393.850000 956.000000 394.150000 ;
        RECT 951.000000 397.850000 956.000000 398.150000 ;
        RECT 951.000000 405.850000 956.000000 406.150000 ;
        RECT 951.000000 401.850000 956.000000 402.150000 ;
        RECT 951.000000 413.850000 956.000000 414.150000 ;
        RECT 951.000000 409.850000 956.000000 410.150000 ;
        RECT 1001.000000 349.850000 1006.000000 350.150000 ;
        RECT 1001.000000 345.850000 1006.000000 346.150000 ;
        RECT 1001.000000 353.850000 1006.000000 354.150000 ;
        RECT 1001.000000 357.850000 1006.000000 358.150000 ;
        RECT 1001.000000 361.850000 1006.000000 362.150000 ;
        RECT 1001.000000 365.850000 1006.000000 366.150000 ;
        RECT 1001.000000 369.850000 1006.000000 370.150000 ;
        RECT 1001.000000 377.850000 1006.000000 378.150000 ;
        RECT 1001.000000 373.850000 1006.000000 374.150000 ;
        RECT 1001.000000 385.850000 1006.000000 386.150000 ;
        RECT 1001.000000 381.850000 1006.000000 382.150000 ;
        RECT 1001.000000 393.850000 1006.000000 394.150000 ;
        RECT 1001.000000 389.850000 1006.000000 390.150000 ;
        RECT 1001.000000 397.850000 1006.000000 398.150000 ;
        RECT 1001.000000 405.850000 1006.000000 406.150000 ;
        RECT 1001.000000 401.850000 1006.000000 402.150000 ;
        RECT 1001.000000 409.850000 1006.000000 410.150000 ;
        RECT 1001.000000 413.850000 1006.000000 414.150000 ;
        RECT 901.000000 417.850000 906.000000 418.150000 ;
        RECT 901.000000 421.850000 906.000000 422.150000 ;
        RECT 901.000000 425.850000 906.000000 426.150000 ;
        RECT 901.000000 433.850000 906.000000 434.150000 ;
        RECT 901.000000 429.850000 906.000000 430.150000 ;
        RECT 901.000000 437.850000 906.000000 438.150000 ;
        RECT 901.000000 441.850000 906.000000 442.150000 ;
        RECT 951.000000 417.850000 956.000000 418.150000 ;
        RECT 951.000000 421.850000 956.000000 422.150000 ;
        RECT 951.000000 425.850000 956.000000 426.150000 ;
        RECT 951.000000 429.850000 956.000000 430.150000 ;
        RECT 951.000000 433.850000 956.000000 434.150000 ;
        RECT 951.000000 441.850000 956.000000 442.150000 ;
        RECT 951.000000 437.850000 956.000000 438.150000 ;
        RECT 1001.000000 425.850000 1006.000000 426.150000 ;
        RECT 1001.000000 421.850000 1006.000000 422.150000 ;
        RECT 1001.000000 417.850000 1006.000000 418.150000 ;
        RECT 1001.000000 429.850000 1006.000000 430.150000 ;
        RECT 1001.000000 433.850000 1006.000000 434.150000 ;
        RECT 1001.000000 437.850000 1006.000000 438.150000 ;
        RECT 1001.000000 441.850000 1006.000000 442.150000 ;
        RECT 1051.000000 357.850000 1056.000000 358.150000 ;
        RECT 1051.000000 353.850000 1056.000000 354.150000 ;
        RECT 1051.000000 349.850000 1056.000000 350.150000 ;
        RECT 1051.000000 345.850000 1056.000000 346.150000 ;
        RECT 1051.000000 361.850000 1056.000000 362.150000 ;
        RECT 1051.000000 365.850000 1056.000000 366.150000 ;
        RECT 1051.000000 369.850000 1056.000000 370.150000 ;
        RECT 1051.000000 373.850000 1056.000000 374.150000 ;
        RECT 1051.000000 377.850000 1056.000000 378.150000 ;
        RECT 1101.000000 345.850000 1106.000000 346.150000 ;
        RECT 1101.000000 349.850000 1106.000000 350.150000 ;
        RECT 1101.000000 353.850000 1106.000000 354.150000 ;
        RECT 1101.000000 357.850000 1106.000000 358.150000 ;
        RECT 1101.000000 361.850000 1106.000000 362.150000 ;
        RECT 1101.000000 365.850000 1106.000000 366.150000 ;
        RECT 1101.000000 369.850000 1106.000000 370.150000 ;
        RECT 1101.000000 373.850000 1106.000000 374.150000 ;
        RECT 1101.000000 377.850000 1106.000000 378.150000 ;
        RECT 1051.000000 385.850000 1056.000000 386.150000 ;
        RECT 1051.000000 381.850000 1056.000000 382.150000 ;
        RECT 1051.000000 393.850000 1056.000000 394.150000 ;
        RECT 1051.000000 389.850000 1056.000000 390.150000 ;
        RECT 1051.000000 397.850000 1056.000000 398.150000 ;
        RECT 1051.000000 405.850000 1056.000000 406.150000 ;
        RECT 1051.000000 401.850000 1056.000000 402.150000 ;
        RECT 1051.000000 409.850000 1056.000000 410.150000 ;
        RECT 1051.000000 413.850000 1056.000000 414.150000 ;
        RECT 1101.000000 397.850000 1106.000000 398.150000 ;
        RECT 1101.000000 393.850000 1106.000000 394.150000 ;
        RECT 1101.000000 389.850000 1106.000000 390.150000 ;
        RECT 1101.000000 381.850000 1106.000000 382.150000 ;
        RECT 1101.000000 385.850000 1106.000000 386.150000 ;
        RECT 1101.000000 405.850000 1106.000000 406.150000 ;
        RECT 1101.000000 401.850000 1106.000000 402.150000 ;
        RECT 1101.000000 413.850000 1106.000000 414.150000 ;
        RECT 1101.000000 409.850000 1106.000000 410.150000 ;
        RECT 1151.000000 357.850000 1156.000000 358.150000 ;
        RECT 1151.000000 353.850000 1156.000000 354.150000 ;
        RECT 1151.000000 349.850000 1156.000000 350.150000 ;
        RECT 1151.000000 345.850000 1156.000000 346.150000 ;
        RECT 1172.000000 357.850000 1182.000000 358.150000 ;
        RECT 1172.000000 349.850000 1182.000000 350.150000 ;
        RECT 1172.000000 345.850000 1182.000000 346.150000 ;
        RECT 1172.000000 353.850000 1182.000000 354.150000 ;
        RECT 1151.000000 365.850000 1156.000000 366.150000 ;
        RECT 1151.000000 361.850000 1156.000000 362.150000 ;
        RECT 1151.000000 369.850000 1156.000000 370.150000 ;
        RECT 1151.000000 373.850000 1156.000000 374.150000 ;
        RECT 1151.000000 377.850000 1156.000000 378.150000 ;
        RECT 1172.000000 369.850000 1182.000000 370.150000 ;
        RECT 1172.000000 365.850000 1182.000000 366.150000 ;
        RECT 1172.000000 361.850000 1182.000000 362.150000 ;
        RECT 1172.000000 373.850000 1182.000000 374.150000 ;
        RECT 1172.000000 377.850000 1182.000000 378.150000 ;
        RECT 1151.000000 385.850000 1156.000000 386.150000 ;
        RECT 1151.000000 381.850000 1156.000000 382.150000 ;
        RECT 1151.000000 393.850000 1156.000000 394.150000 ;
        RECT 1151.000000 389.850000 1156.000000 390.150000 ;
        RECT 1151.000000 397.850000 1156.000000 398.150000 ;
        RECT 1172.000000 385.850000 1182.000000 386.150000 ;
        RECT 1172.000000 381.850000 1182.000000 382.150000 ;
        RECT 1172.000000 389.850000 1182.000000 390.150000 ;
        RECT 1172.000000 393.850000 1182.000000 394.150000 ;
        RECT 1172.000000 397.850000 1182.000000 398.150000 ;
        RECT 1151.000000 405.850000 1156.000000 406.150000 ;
        RECT 1151.000000 401.850000 1156.000000 402.150000 ;
        RECT 1151.000000 409.850000 1156.000000 410.150000 ;
        RECT 1151.000000 413.850000 1156.000000 414.150000 ;
        RECT 1172.000000 405.850000 1182.000000 406.150000 ;
        RECT 1172.000000 401.850000 1182.000000 402.150000 ;
        RECT 1172.000000 409.850000 1182.000000 410.150000 ;
        RECT 1172.000000 413.850000 1182.000000 414.150000 ;
        RECT 1051.000000 417.850000 1056.000000 418.150000 ;
        RECT 1051.000000 421.850000 1056.000000 422.150000 ;
        RECT 1051.000000 425.850000 1056.000000 426.150000 ;
        RECT 1051.000000 429.850000 1056.000000 430.150000 ;
        RECT 1051.000000 433.850000 1056.000000 434.150000 ;
        RECT 1051.000000 437.850000 1056.000000 438.150000 ;
        RECT 1051.000000 441.850000 1056.000000 442.150000 ;
        RECT 1101.000000 433.850000 1106.000000 434.150000 ;
        RECT 1101.000000 429.850000 1106.000000 430.150000 ;
        RECT 1101.000000 425.850000 1106.000000 426.150000 ;
        RECT 1101.000000 421.850000 1106.000000 422.150000 ;
        RECT 1101.000000 417.850000 1106.000000 418.150000 ;
        RECT 1101.000000 441.850000 1106.000000 442.150000 ;
        RECT 1101.000000 437.850000 1106.000000 438.150000 ;
        RECT 1151.000000 417.850000 1156.000000 418.150000 ;
        RECT 1151.000000 421.850000 1156.000000 422.150000 ;
        RECT 1151.000000 425.850000 1156.000000 426.150000 ;
        RECT 1151.000000 429.850000 1156.000000 430.150000 ;
        RECT 1151.000000 433.850000 1156.000000 434.150000 ;
        RECT 1172.000000 417.850000 1182.000000 418.150000 ;
        RECT 1172.000000 421.850000 1182.000000 422.150000 ;
        RECT 1172.000000 425.850000 1182.000000 426.150000 ;
        RECT 1172.000000 429.850000 1182.000000 430.150000 ;
        RECT 1172.000000 433.850000 1182.000000 434.150000 ;
        RECT 1151.000000 437.850000 1156.000000 438.150000 ;
        RECT 1151.000000 441.850000 1156.000000 442.150000 ;
        RECT 1151.000000 453.850000 1156.000000 454.150000 ;
        RECT 1151.000000 449.850000 1156.000000 450.150000 ;
        RECT 1151.000000 445.850000 1156.000000 446.150000 ;
        RECT 1172.000000 437.850000 1182.000000 438.150000 ;
        RECT 1172.000000 441.850000 1182.000000 442.150000 ;
        RECT 1151.000000 461.850000 1156.000000 462.150000 ;
        RECT 1151.000000 457.850000 1156.000000 458.150000 ;
        RECT 1151.000000 465.850000 1156.000000 466.150000 ;
        RECT 1151.000000 469.850000 1156.000000 470.150000 ;
        RECT 1151.000000 481.850000 1156.000000 482.150000 ;
        RECT 1151.000000 477.850000 1156.000000 478.150000 ;
        RECT 1151.000000 473.850000 1156.000000 474.150000 ;
        RECT 1151.000000 489.850000 1156.000000 490.150000 ;
        RECT 1151.000000 485.850000 1156.000000 486.150000 ;
        RECT 1151.000000 493.850000 1156.000000 494.150000 ;
        RECT 1151.000000 497.850000 1156.000000 498.150000 ;
        RECT 1151.000000 505.850000 1156.000000 506.150000 ;
        RECT 1151.000000 501.850000 1156.000000 502.150000 ;
        RECT 1151.000000 509.850000 1156.000000 510.150000 ;
        RECT 1151.000000 513.850000 1156.000000 514.150000 ;
        RECT 1151.000000 517.850000 1156.000000 518.150000 ;
        RECT 1151.000000 521.850000 1156.000000 522.150000 ;
        RECT 1151.000000 525.850000 1156.000000 526.150000 ;
        RECT 1151.000000 533.850000 1156.000000 534.150000 ;
        RECT 1151.000000 529.850000 1156.000000 530.150000 ;
        RECT 1151.000000 545.850000 1156.000000 546.150000 ;
        RECT 1151.000000 537.850000 1156.000000 538.150000 ;
        RECT 1151.000000 541.850000 1156.000000 542.150000 ;
        RECT 1151.000000 553.850000 1156.000000 554.150000 ;
        RECT 1151.000000 549.850000 1156.000000 550.150000 ;
        RECT 1151.000000 561.850000 1156.000000 562.150000 ;
        RECT 1151.000000 557.850000 1156.000000 558.150000 ;
        RECT 1151.000000 565.850000 1156.000000 566.150000 ;
        RECT 1151.000000 569.850000 1156.000000 570.150000 ;
        RECT 1151.000000 573.850000 1156.000000 574.150000 ;
        RECT 1151.000000 577.850000 1156.000000 578.150000 ;
        RECT 1151.000000 581.850000 1156.000000 582.150000 ;
        RECT 1151.000000 589.850000 1156.000000 590.150000 ;
        RECT 1151.000000 585.850000 1156.000000 586.150000 ;
        RECT 1151.000000 593.850000 1156.000000 594.150000 ;
        RECT 1151.000000 597.850000 1156.000000 598.150000 ;
        RECT 1151.000000 601.850000 1156.000000 602.150000 ;
        RECT 1151.000000 609.850000 1156.000000 610.150000 ;
        RECT 1151.000000 605.850000 1156.000000 606.150000 ;
        RECT 1151.000000 613.850000 1156.000000 614.150000 ;
        RECT 1151.000000 617.850000 1156.000000 618.150000 ;
        RECT 1151.000000 621.850000 1156.000000 622.150000 ;
        RECT 1151.000000 625.850000 1156.000000 626.150000 ;
        RECT 1151.000000 629.850000 1156.000000 630.150000 ;
        RECT 1151.000000 637.850000 1156.000000 638.150000 ;
        RECT 1151.000000 633.850000 1156.000000 634.150000 ;
        RECT 601.000000 657.850000 606.000000 658.150000 ;
        RECT 601.000000 673.850000 606.000000 674.150000 ;
        RECT 601.000000 669.850000 606.000000 670.150000 ;
        RECT 601.000000 665.850000 606.000000 666.150000 ;
        RECT 601.000000 661.850000 606.000000 662.150000 ;
        RECT 651.000000 657.850000 656.000000 658.150000 ;
        RECT 651.000000 665.850000 656.000000 666.150000 ;
        RECT 651.000000 661.850000 656.000000 662.150000 ;
        RECT 651.000000 673.850000 656.000000 674.150000 ;
        RECT 651.000000 669.850000 656.000000 670.150000 ;
        RECT 601.000000 677.850000 606.000000 678.150000 ;
        RECT 601.000000 681.850000 606.000000 682.150000 ;
        RECT 651.000000 677.850000 656.000000 678.150000 ;
        RECT 651.000000 681.850000 656.000000 682.150000 ;
        RECT 1151.000000 657.850000 1156.000000 658.150000 ;
        RECT 1151.000000 641.850000 1156.000000 642.150000 ;
        RECT 1151.000000 645.850000 1156.000000 646.150000 ;
        RECT 1151.000000 649.850000 1156.000000 650.150000 ;
        RECT 1151.000000 653.850000 1156.000000 654.150000 ;
        RECT 1151.000000 665.850000 1156.000000 666.150000 ;
        RECT 1151.000000 661.850000 1156.000000 662.150000 ;
        RECT 1151.000000 669.850000 1156.000000 670.150000 ;
        RECT 1151.000000 673.850000 1156.000000 674.150000 ;
        RECT 1151.000000 681.850000 1156.000000 682.150000 ;
        RECT 1151.000000 677.850000 1156.000000 678.150000 ;
      LAYER M3 ;
        RECT 4.000000 5.850000 14.000000 6.150000 ;
        RECT 51.000000 5.850000 56.000000 6.150000 ;
        RECT 51.000000 1.850000 56.000000 2.150000 ;
        RECT 101.000000 1.850000 106.000000 2.150000 ;
        RECT 101.000000 5.850000 106.000000 6.150000 ;
        RECT 151.000000 1.850000 156.000000 2.150000 ;
        RECT 151.000000 5.850000 156.000000 6.150000 ;
        RECT 201.000000 1.850000 206.000000 2.150000 ;
        RECT 201.000000 5.850000 206.000000 6.150000 ;
        RECT 251.000000 1.850000 256.000000 2.150000 ;
        RECT 251.000000 5.850000 256.000000 6.150000 ;
        RECT 301.000000 1.850000 306.000000 2.150000 ;
        RECT 301.000000 5.850000 306.000000 6.150000 ;
        RECT 351.000000 1.850000 356.000000 2.150000 ;
        RECT 351.000000 5.850000 356.000000 6.150000 ;
        RECT 401.000000 1.850000 406.000000 2.150000 ;
        RECT 401.000000 5.850000 406.000000 6.150000 ;
        RECT 451.000000 1.850000 456.000000 2.150000 ;
        RECT 451.000000 5.850000 456.000000 6.150000 ;
        RECT 501.000000 1.850000 506.000000 2.150000 ;
        RECT 501.000000 5.850000 506.000000 6.150000 ;
        RECT 551.000000 1.850000 556.000000 2.150000 ;
        RECT 551.000000 5.850000 556.000000 6.150000 ;
        RECT 4.000000 265.850000 14.000000 266.150000 ;
        RECT 4.000000 261.850000 14.000000 262.150000 ;
        RECT 51.000000 265.850000 56.000000 266.150000 ;
        RECT 51.000000 261.850000 56.000000 262.150000 ;
        RECT 101.000000 265.850000 106.000000 266.150000 ;
        RECT 101.000000 261.850000 106.000000 262.150000 ;
        RECT 51.000000 305.850000 56.000000 306.150000 ;
        RECT 4.000000 305.850000 14.000000 306.150000 ;
        RECT 4.000000 285.850000 14.000000 286.150000 ;
        RECT 4.000000 281.850000 14.000000 282.150000 ;
        RECT 4.000000 269.850000 14.000000 270.150000 ;
        RECT 4.000000 273.850000 14.000000 274.150000 ;
        RECT 4.000000 277.850000 14.000000 278.150000 ;
        RECT 4.000000 289.850000 14.000000 290.150000 ;
        RECT 4.000000 293.850000 14.000000 294.150000 ;
        RECT 4.000000 297.850000 14.000000 298.150000 ;
        RECT 4.000000 301.850000 14.000000 302.150000 ;
        RECT 51.000000 269.850000 56.000000 270.150000 ;
        RECT 51.000000 273.850000 56.000000 274.150000 ;
        RECT 51.000000 277.850000 56.000000 278.150000 ;
        RECT 51.000000 281.850000 56.000000 282.150000 ;
        RECT 51.000000 285.850000 56.000000 286.150000 ;
        RECT 51.000000 301.850000 56.000000 302.150000 ;
        RECT 51.000000 297.850000 56.000000 298.150000 ;
        RECT 51.000000 293.850000 56.000000 294.150000 ;
        RECT 51.000000 289.850000 56.000000 290.150000 ;
        RECT 4.000000 321.850000 14.000000 322.150000 ;
        RECT 4.000000 309.850000 14.000000 310.150000 ;
        RECT 4.000000 313.850000 14.000000 314.150000 ;
        RECT 4.000000 317.850000 14.000000 318.150000 ;
        RECT 4.000000 325.850000 14.000000 326.150000 ;
        RECT 4.000000 329.850000 14.000000 330.150000 ;
        RECT 4.000000 333.850000 14.000000 334.150000 ;
        RECT 4.000000 337.850000 14.000000 338.150000 ;
        RECT 4.000000 341.850000 14.000000 342.150000 ;
        RECT 51.000000 313.850000 56.000000 314.150000 ;
        RECT 51.000000 309.850000 56.000000 310.150000 ;
        RECT 51.000000 317.850000 56.000000 318.150000 ;
        RECT 51.000000 321.850000 56.000000 322.150000 ;
        RECT 51.000000 341.850000 56.000000 342.150000 ;
        RECT 51.000000 337.850000 56.000000 338.150000 ;
        RECT 51.000000 333.850000 56.000000 334.150000 ;
        RECT 51.000000 329.850000 56.000000 330.150000 ;
        RECT 51.000000 325.850000 56.000000 326.150000 ;
        RECT 101.000000 305.850000 106.000000 306.150000 ;
        RECT 101.000000 269.850000 106.000000 270.150000 ;
        RECT 101.000000 273.850000 106.000000 274.150000 ;
        RECT 101.000000 277.850000 106.000000 278.150000 ;
        RECT 101.000000 281.850000 106.000000 282.150000 ;
        RECT 101.000000 285.850000 106.000000 286.150000 ;
        RECT 101.000000 301.850000 106.000000 302.150000 ;
        RECT 101.000000 297.850000 106.000000 298.150000 ;
        RECT 101.000000 293.850000 106.000000 294.150000 ;
        RECT 101.000000 289.850000 106.000000 290.150000 ;
        RECT 101.000000 321.850000 106.000000 322.150000 ;
        RECT 101.000000 317.850000 106.000000 318.150000 ;
        RECT 101.000000 313.850000 106.000000 314.150000 ;
        RECT 101.000000 309.850000 106.000000 310.150000 ;
        RECT 101.000000 325.850000 106.000000 326.150000 ;
        RECT 101.000000 329.850000 106.000000 330.150000 ;
        RECT 101.000000 333.850000 106.000000 334.150000 ;
        RECT 101.000000 337.850000 106.000000 338.150000 ;
        RECT 101.000000 341.850000 106.000000 342.150000 ;
        RECT 151.000000 261.850000 156.000000 262.150000 ;
        RECT 151.000000 265.850000 156.000000 266.150000 ;
        RECT 201.000000 265.850000 206.000000 266.150000 ;
        RECT 201.000000 261.850000 206.000000 262.150000 ;
        RECT 251.000000 265.850000 256.000000 266.150000 ;
        RECT 251.000000 261.850000 256.000000 262.150000 ;
        RECT 201.000000 305.850000 206.000000 306.150000 ;
        RECT 151.000000 305.850000 156.000000 306.150000 ;
        RECT 151.000000 277.850000 156.000000 278.150000 ;
        RECT 151.000000 273.850000 156.000000 274.150000 ;
        RECT 151.000000 269.850000 156.000000 270.150000 ;
        RECT 151.000000 281.850000 156.000000 282.150000 ;
        RECT 151.000000 285.850000 156.000000 286.150000 ;
        RECT 151.000000 289.850000 156.000000 290.150000 ;
        RECT 151.000000 293.850000 156.000000 294.150000 ;
        RECT 151.000000 301.850000 156.000000 302.150000 ;
        RECT 151.000000 297.850000 156.000000 298.150000 ;
        RECT 201.000000 269.850000 206.000000 270.150000 ;
        RECT 201.000000 273.850000 206.000000 274.150000 ;
        RECT 201.000000 277.850000 206.000000 278.150000 ;
        RECT 201.000000 281.850000 206.000000 282.150000 ;
        RECT 201.000000 285.850000 206.000000 286.150000 ;
        RECT 201.000000 301.850000 206.000000 302.150000 ;
        RECT 201.000000 297.850000 206.000000 298.150000 ;
        RECT 201.000000 293.850000 206.000000 294.150000 ;
        RECT 201.000000 289.850000 206.000000 290.150000 ;
        RECT 151.000000 313.850000 156.000000 314.150000 ;
        RECT 151.000000 309.850000 156.000000 310.150000 ;
        RECT 151.000000 321.850000 156.000000 322.150000 ;
        RECT 151.000000 317.850000 156.000000 318.150000 ;
        RECT 151.000000 329.850000 156.000000 330.150000 ;
        RECT 151.000000 325.850000 156.000000 326.150000 ;
        RECT 151.000000 333.850000 156.000000 334.150000 ;
        RECT 151.000000 337.850000 156.000000 338.150000 ;
        RECT 151.000000 341.850000 156.000000 342.150000 ;
        RECT 201.000000 313.850000 206.000000 314.150000 ;
        RECT 201.000000 309.850000 206.000000 310.150000 ;
        RECT 201.000000 317.850000 206.000000 318.150000 ;
        RECT 201.000000 321.850000 206.000000 322.150000 ;
        RECT 201.000000 341.850000 206.000000 342.150000 ;
        RECT 201.000000 337.850000 206.000000 338.150000 ;
        RECT 201.000000 333.850000 206.000000 334.150000 ;
        RECT 201.000000 329.850000 206.000000 330.150000 ;
        RECT 201.000000 325.850000 206.000000 326.150000 ;
        RECT 251.000000 305.850000 256.000000 306.150000 ;
        RECT 251.000000 269.850000 256.000000 270.150000 ;
        RECT 251.000000 273.850000 256.000000 274.150000 ;
        RECT 251.000000 277.850000 256.000000 278.150000 ;
        RECT 251.000000 281.850000 256.000000 282.150000 ;
        RECT 251.000000 285.850000 256.000000 286.150000 ;
        RECT 251.000000 293.850000 256.000000 294.150000 ;
        RECT 251.000000 289.850000 256.000000 290.150000 ;
        RECT 251.000000 297.850000 256.000000 298.150000 ;
        RECT 251.000000 301.850000 256.000000 302.150000 ;
        RECT 251.000000 309.850000 256.000000 310.150000 ;
        RECT 251.000000 313.850000 256.000000 314.150000 ;
        RECT 251.000000 321.850000 256.000000 322.150000 ;
        RECT 251.000000 317.850000 256.000000 318.150000 ;
        RECT 251.000000 325.850000 256.000000 326.150000 ;
        RECT 251.000000 329.850000 256.000000 330.150000 ;
        RECT 251.000000 333.850000 256.000000 334.150000 ;
        RECT 251.000000 337.850000 256.000000 338.150000 ;
        RECT 251.000000 341.850000 256.000000 342.150000 ;
        RECT 301.000000 265.850000 306.000000 266.150000 ;
        RECT 301.000000 261.850000 306.000000 262.150000 ;
        RECT 351.000000 265.850000 356.000000 266.150000 ;
        RECT 351.000000 261.850000 356.000000 262.150000 ;
        RECT 401.000000 261.850000 406.000000 262.150000 ;
        RECT 401.000000 265.850000 406.000000 266.150000 ;
        RECT 301.000000 305.850000 306.000000 306.150000 ;
        RECT 351.000000 305.850000 356.000000 306.150000 ;
        RECT 301.000000 277.850000 306.000000 278.150000 ;
        RECT 301.000000 269.850000 306.000000 270.150000 ;
        RECT 301.000000 273.850000 306.000000 274.150000 ;
        RECT 301.000000 281.850000 306.000000 282.150000 ;
        RECT 301.000000 285.850000 306.000000 286.150000 ;
        RECT 301.000000 293.850000 306.000000 294.150000 ;
        RECT 301.000000 289.850000 306.000000 290.150000 ;
        RECT 301.000000 301.850000 306.000000 302.150000 ;
        RECT 301.000000 297.850000 306.000000 298.150000 ;
        RECT 351.000000 269.850000 356.000000 270.150000 ;
        RECT 351.000000 273.850000 356.000000 274.150000 ;
        RECT 351.000000 277.850000 356.000000 278.150000 ;
        RECT 351.000000 281.850000 356.000000 282.150000 ;
        RECT 351.000000 285.850000 356.000000 286.150000 ;
        RECT 351.000000 289.850000 356.000000 290.150000 ;
        RECT 351.000000 293.850000 356.000000 294.150000 ;
        RECT 351.000000 297.850000 356.000000 298.150000 ;
        RECT 351.000000 301.850000 356.000000 302.150000 ;
        RECT 301.000000 313.850000 306.000000 314.150000 ;
        RECT 301.000000 309.850000 306.000000 310.150000 ;
        RECT 301.000000 317.850000 306.000000 318.150000 ;
        RECT 301.000000 321.850000 306.000000 322.150000 ;
        RECT 301.000000 329.850000 306.000000 330.150000 ;
        RECT 301.000000 325.850000 306.000000 326.150000 ;
        RECT 301.000000 341.850000 306.000000 342.150000 ;
        RECT 301.000000 337.850000 306.000000 338.150000 ;
        RECT 301.000000 333.850000 306.000000 334.150000 ;
        RECT 351.000000 313.850000 356.000000 314.150000 ;
        RECT 351.000000 309.850000 356.000000 310.150000 ;
        RECT 351.000000 317.850000 356.000000 318.150000 ;
        RECT 351.000000 321.850000 356.000000 322.150000 ;
        RECT 351.000000 341.850000 356.000000 342.150000 ;
        RECT 351.000000 337.850000 356.000000 338.150000 ;
        RECT 351.000000 333.850000 356.000000 334.150000 ;
        RECT 351.000000 329.850000 356.000000 330.150000 ;
        RECT 351.000000 325.850000 356.000000 326.150000 ;
        RECT 401.000000 305.850000 406.000000 306.150000 ;
        RECT 401.000000 273.850000 406.000000 274.150000 ;
        RECT 401.000000 269.850000 406.000000 270.150000 ;
        RECT 401.000000 277.850000 406.000000 278.150000 ;
        RECT 401.000000 281.850000 406.000000 282.150000 ;
        RECT 401.000000 285.850000 406.000000 286.150000 ;
        RECT 401.000000 293.850000 406.000000 294.150000 ;
        RECT 401.000000 289.850000 406.000000 290.150000 ;
        RECT 401.000000 297.850000 406.000000 298.150000 ;
        RECT 401.000000 301.850000 406.000000 302.150000 ;
        RECT 401.000000 309.850000 406.000000 310.150000 ;
        RECT 401.000000 313.850000 406.000000 314.150000 ;
        RECT 401.000000 317.850000 406.000000 318.150000 ;
        RECT 401.000000 321.850000 406.000000 322.150000 ;
        RECT 401.000000 329.850000 406.000000 330.150000 ;
        RECT 401.000000 325.850000 406.000000 326.150000 ;
        RECT 401.000000 333.850000 406.000000 334.150000 ;
        RECT 401.000000 337.850000 406.000000 338.150000 ;
        RECT 401.000000 341.850000 406.000000 342.150000 ;
        RECT 451.000000 265.850000 456.000000 266.150000 ;
        RECT 451.000000 261.850000 456.000000 262.150000 ;
        RECT 501.000000 261.850000 506.000000 262.150000 ;
        RECT 501.000000 265.850000 506.000000 266.150000 ;
        RECT 551.000000 265.850000 556.000000 266.150000 ;
        RECT 551.000000 261.850000 556.000000 262.150000 ;
        RECT 501.000000 305.850000 506.000000 306.150000 ;
        RECT 451.000000 277.850000 456.000000 278.150000 ;
        RECT 451.000000 273.850000 456.000000 274.150000 ;
        RECT 451.000000 269.850000 456.000000 270.150000 ;
        RECT 451.000000 285.850000 456.000000 286.150000 ;
        RECT 451.000000 281.850000 456.000000 282.150000 ;
        RECT 451.000000 293.850000 456.000000 294.150000 ;
        RECT 451.000000 289.850000 456.000000 290.150000 ;
        RECT 451.000000 297.850000 456.000000 298.150000 ;
        RECT 501.000000 277.850000 506.000000 278.150000 ;
        RECT 501.000000 269.850000 506.000000 270.150000 ;
        RECT 501.000000 273.850000 506.000000 274.150000 ;
        RECT 501.000000 281.850000 506.000000 282.150000 ;
        RECT 501.000000 285.850000 506.000000 286.150000 ;
        RECT 501.000000 289.850000 506.000000 290.150000 ;
        RECT 501.000000 293.850000 506.000000 294.150000 ;
        RECT 501.000000 301.850000 506.000000 302.150000 ;
        RECT 501.000000 297.850000 506.000000 298.150000 ;
        RECT 451.000000 316.105000 456.000000 317.105000 ;
        RECT 451.000000 321.850000 456.000000 322.150000 ;
        RECT 451.000000 333.850000 456.000000 334.150000 ;
        RECT 451.000000 329.850000 456.000000 330.150000 ;
        RECT 451.000000 325.850000 456.000000 326.150000 ;
        RECT 451.000000 337.850000 456.000000 338.150000 ;
        RECT 451.000000 341.850000 456.000000 342.150000 ;
        RECT 501.000000 313.850000 506.000000 314.150000 ;
        RECT 501.000000 309.850000 506.000000 310.150000 ;
        RECT 501.000000 317.850000 506.000000 318.150000 ;
        RECT 501.000000 321.850000 506.000000 322.150000 ;
        RECT 501.000000 329.850000 506.000000 330.150000 ;
        RECT 501.000000 325.850000 506.000000 326.150000 ;
        RECT 501.000000 333.850000 506.000000 334.150000 ;
        RECT 501.000000 337.850000 506.000000 338.150000 ;
        RECT 501.000000 341.850000 506.000000 342.150000 ;
        RECT 551.000000 305.850000 556.000000 306.150000 ;
        RECT 551.000000 277.850000 556.000000 278.150000 ;
        RECT 551.000000 269.850000 556.000000 270.150000 ;
        RECT 551.000000 273.850000 556.000000 274.150000 ;
        RECT 551.000000 281.850000 556.000000 282.150000 ;
        RECT 551.000000 285.850000 556.000000 286.150000 ;
        RECT 551.000000 301.850000 556.000000 302.150000 ;
        RECT 551.000000 297.850000 556.000000 298.150000 ;
        RECT 551.000000 293.850000 556.000000 294.150000 ;
        RECT 551.000000 289.850000 556.000000 290.150000 ;
        RECT 551.000000 309.850000 556.000000 310.150000 ;
        RECT 551.000000 313.850000 556.000000 314.150000 ;
        RECT 551.000000 317.850000 556.000000 318.150000 ;
        RECT 551.000000 321.850000 556.000000 322.150000 ;
        RECT 551.000000 325.850000 556.000000 326.150000 ;
        RECT 551.000000 329.850000 556.000000 330.150000 ;
        RECT 551.000000 333.850000 556.000000 334.150000 ;
        RECT 551.000000 337.850000 556.000000 338.150000 ;
        RECT 551.000000 341.850000 556.000000 342.150000 ;
        RECT 601.000000 1.850000 606.000000 2.150000 ;
        RECT 601.000000 5.850000 606.000000 6.150000 ;
        RECT 651.000000 1.850000 656.000000 2.150000 ;
        RECT 651.000000 5.850000 656.000000 6.150000 ;
        RECT 701.000000 1.850000 706.000000 2.150000 ;
        RECT 701.000000 5.850000 706.000000 6.150000 ;
        RECT 751.000000 1.850000 756.000000 2.150000 ;
        RECT 751.000000 5.850000 756.000000 6.150000 ;
        RECT 801.000000 1.850000 806.000000 2.150000 ;
        RECT 801.000000 5.850000 806.000000 6.150000 ;
        RECT 851.000000 1.850000 856.000000 2.150000 ;
        RECT 851.000000 5.850000 856.000000 6.150000 ;
        RECT 901.000000 1.850000 906.000000 2.150000 ;
        RECT 901.000000 5.850000 906.000000 6.150000 ;
        RECT 951.000000 1.850000 956.000000 2.150000 ;
        RECT 951.000000 5.850000 956.000000 6.150000 ;
        RECT 1001.000000 1.850000 1006.000000 2.150000 ;
        RECT 1001.000000 5.850000 1006.000000 6.150000 ;
        RECT 1051.000000 1.850000 1056.000000 2.150000 ;
        RECT 1051.000000 5.850000 1056.000000 6.150000 ;
        RECT 1101.000000 1.850000 1106.000000 2.150000 ;
        RECT 1101.000000 5.850000 1106.000000 6.150000 ;
        RECT 1151.000000 5.850000 1156.000000 6.150000 ;
        RECT 1172.000000 5.850000 1182.000000 6.150000 ;
        RECT 1151.000000 1.850000 1156.000000 2.150000 ;
        RECT 1172.000000 17.850000 1182.000000 18.150000 ;
        RECT 1172.000000 13.850000 1182.000000 14.150000 ;
        RECT 1172.000000 9.850000 1182.000000 10.150000 ;
        RECT 1172.000000 21.850000 1182.000000 22.150000 ;
        RECT 1172.000000 25.850000 1182.000000 26.150000 ;
        RECT 1172.000000 33.850000 1182.000000 34.150000 ;
        RECT 1172.000000 29.850000 1182.000000 30.150000 ;
        RECT 1172.000000 41.850000 1182.000000 42.150000 ;
        RECT 1172.000000 37.850000 1182.000000 38.150000 ;
        RECT 1172.000000 45.850000 1182.000000 46.150000 ;
        RECT 601.000000 265.850000 606.000000 266.150000 ;
        RECT 601.000000 261.850000 606.000000 262.150000 ;
        RECT 651.000000 261.850000 656.000000 262.150000 ;
        RECT 651.000000 265.850000 656.000000 266.150000 ;
        RECT 701.000000 265.850000 706.000000 266.150000 ;
        RECT 701.000000 261.850000 706.000000 262.150000 ;
        RECT 601.000000 305.850000 606.000000 306.150000 ;
        RECT 651.000000 305.850000 656.000000 306.150000 ;
        RECT 601.000000 277.850000 606.000000 278.150000 ;
        RECT 601.000000 269.850000 606.000000 270.150000 ;
        RECT 601.000000 273.850000 606.000000 274.150000 ;
        RECT 601.000000 281.850000 606.000000 282.150000 ;
        RECT 601.000000 285.850000 606.000000 286.150000 ;
        RECT 601.000000 289.850000 606.000000 290.150000 ;
        RECT 601.000000 293.850000 606.000000 294.150000 ;
        RECT 601.000000 297.850000 606.000000 298.150000 ;
        RECT 601.000000 301.850000 606.000000 302.150000 ;
        RECT 651.000000 277.850000 656.000000 278.150000 ;
        RECT 651.000000 273.850000 656.000000 274.150000 ;
        RECT 651.000000 269.850000 656.000000 270.150000 ;
        RECT 651.000000 281.850000 656.000000 282.150000 ;
        RECT 651.000000 285.850000 656.000000 286.150000 ;
        RECT 651.000000 289.850000 656.000000 290.150000 ;
        RECT 651.000000 293.850000 656.000000 294.150000 ;
        RECT 651.000000 301.850000 656.000000 302.150000 ;
        RECT 651.000000 297.850000 656.000000 298.150000 ;
        RECT 601.000000 321.850000 606.000000 322.150000 ;
        RECT 601.000000 317.850000 606.000000 318.150000 ;
        RECT 601.000000 309.850000 606.000000 310.150000 ;
        RECT 601.000000 313.850000 606.000000 314.150000 ;
        RECT 601.000000 325.850000 606.000000 326.150000 ;
        RECT 601.000000 329.850000 606.000000 330.150000 ;
        RECT 601.000000 333.850000 606.000000 334.150000 ;
        RECT 601.000000 337.850000 606.000000 338.150000 ;
        RECT 601.000000 341.850000 606.000000 342.150000 ;
        RECT 651.000000 313.850000 656.000000 314.150000 ;
        RECT 651.000000 309.850000 656.000000 310.150000 ;
        RECT 651.000000 321.850000 656.000000 322.150000 ;
        RECT 651.000000 317.850000 656.000000 318.150000 ;
        RECT 651.000000 329.850000 656.000000 330.150000 ;
        RECT 651.000000 325.850000 656.000000 326.150000 ;
        RECT 651.000000 333.850000 656.000000 334.150000 ;
        RECT 651.000000 337.850000 656.000000 338.150000 ;
        RECT 651.000000 341.850000 656.000000 342.150000 ;
        RECT 701.000000 305.850000 706.000000 306.150000 ;
        RECT 701.000000 285.850000 706.000000 286.150000 ;
        RECT 701.000000 281.850000 706.000000 282.150000 ;
        RECT 701.000000 277.850000 706.000000 278.150000 ;
        RECT 701.000000 273.850000 706.000000 274.150000 ;
        RECT 701.000000 269.850000 706.000000 270.150000 ;
        RECT 701.000000 301.850000 706.000000 302.150000 ;
        RECT 701.000000 297.850000 706.000000 298.150000 ;
        RECT 701.000000 293.850000 706.000000 294.150000 ;
        RECT 701.000000 289.850000 706.000000 290.150000 ;
        RECT 701.000000 309.850000 706.000000 310.150000 ;
        RECT 701.000000 313.850000 706.000000 314.150000 ;
        RECT 701.000000 317.850000 706.000000 318.150000 ;
        RECT 701.000000 321.850000 706.000000 322.150000 ;
        RECT 701.000000 325.850000 706.000000 326.150000 ;
        RECT 701.000000 329.850000 706.000000 330.150000 ;
        RECT 701.000000 333.850000 706.000000 334.150000 ;
        RECT 701.000000 337.850000 706.000000 338.150000 ;
        RECT 701.000000 341.850000 706.000000 342.150000 ;
        RECT 751.000000 261.850000 756.000000 262.150000 ;
        RECT 751.000000 265.850000 756.000000 266.150000 ;
        RECT 801.000000 261.850000 806.000000 262.150000 ;
        RECT 801.000000 265.850000 806.000000 266.150000 ;
        RECT 851.000000 265.850000 856.000000 266.150000 ;
        RECT 851.000000 261.850000 856.000000 262.150000 ;
        RECT 801.000000 305.850000 806.000000 306.150000 ;
        RECT 751.000000 305.850000 756.000000 306.150000 ;
        RECT 751.000000 285.850000 756.000000 286.150000 ;
        RECT 751.000000 281.850000 756.000000 282.150000 ;
        RECT 751.000000 269.850000 756.000000 270.150000 ;
        RECT 751.000000 273.850000 756.000000 274.150000 ;
        RECT 751.000000 277.850000 756.000000 278.150000 ;
        RECT 751.000000 289.850000 756.000000 290.150000 ;
        RECT 751.000000 293.850000 756.000000 294.150000 ;
        RECT 751.000000 297.850000 756.000000 298.150000 ;
        RECT 751.000000 301.850000 756.000000 302.150000 ;
        RECT 801.000000 277.850000 806.000000 278.150000 ;
        RECT 801.000000 269.850000 806.000000 270.150000 ;
        RECT 801.000000 273.850000 806.000000 274.150000 ;
        RECT 801.000000 281.850000 806.000000 282.150000 ;
        RECT 801.000000 285.850000 806.000000 286.150000 ;
        RECT 801.000000 289.850000 806.000000 290.150000 ;
        RECT 801.000000 293.850000 806.000000 294.150000 ;
        RECT 801.000000 301.850000 806.000000 302.150000 ;
        RECT 801.000000 297.850000 806.000000 298.150000 ;
        RECT 751.000000 321.850000 756.000000 322.150000 ;
        RECT 751.000000 309.850000 756.000000 310.150000 ;
        RECT 751.000000 313.850000 756.000000 314.150000 ;
        RECT 751.000000 317.850000 756.000000 318.150000 ;
        RECT 751.000000 325.850000 756.000000 326.150000 ;
        RECT 751.000000 329.850000 756.000000 330.150000 ;
        RECT 751.000000 333.850000 756.000000 334.150000 ;
        RECT 751.000000 337.850000 756.000000 338.150000 ;
        RECT 751.000000 341.850000 756.000000 342.150000 ;
        RECT 801.000000 313.850000 806.000000 314.150000 ;
        RECT 801.000000 309.850000 806.000000 310.150000 ;
        RECT 801.000000 321.850000 806.000000 322.150000 ;
        RECT 801.000000 317.850000 806.000000 318.150000 ;
        RECT 801.000000 329.850000 806.000000 330.150000 ;
        RECT 801.000000 325.850000 806.000000 326.150000 ;
        RECT 801.000000 333.850000 806.000000 334.150000 ;
        RECT 801.000000 337.850000 806.000000 338.150000 ;
        RECT 801.000000 341.850000 806.000000 342.150000 ;
        RECT 851.000000 305.850000 856.000000 306.150000 ;
        RECT 851.000000 285.850000 856.000000 286.150000 ;
        RECT 851.000000 281.850000 856.000000 282.150000 ;
        RECT 851.000000 277.850000 856.000000 278.150000 ;
        RECT 851.000000 273.850000 856.000000 274.150000 ;
        RECT 851.000000 269.850000 856.000000 270.150000 ;
        RECT 851.000000 301.850000 856.000000 302.150000 ;
        RECT 851.000000 297.850000 856.000000 298.150000 ;
        RECT 851.000000 293.850000 856.000000 294.150000 ;
        RECT 851.000000 289.850000 856.000000 290.150000 ;
        RECT 851.000000 309.850000 856.000000 310.150000 ;
        RECT 851.000000 313.850000 856.000000 314.150000 ;
        RECT 851.000000 317.850000 856.000000 318.150000 ;
        RECT 851.000000 321.850000 856.000000 322.150000 ;
        RECT 851.000000 325.850000 856.000000 326.150000 ;
        RECT 851.000000 329.850000 856.000000 330.150000 ;
        RECT 851.000000 333.850000 856.000000 334.150000 ;
        RECT 851.000000 337.850000 856.000000 338.150000 ;
        RECT 851.000000 341.850000 856.000000 342.150000 ;
        RECT 1172.000000 61.850000 1182.000000 62.150000 ;
        RECT 1172.000000 57.850000 1182.000000 58.150000 ;
        RECT 1172.000000 53.850000 1182.000000 54.150000 ;
        RECT 1172.000000 49.850000 1182.000000 50.150000 ;
        RECT 1172.000000 73.850000 1182.000000 74.150000 ;
        RECT 1172.000000 69.850000 1182.000000 70.150000 ;
        RECT 1172.000000 65.850000 1182.000000 66.150000 ;
        RECT 1172.000000 77.850000 1182.000000 78.150000 ;
        RECT 1172.000000 81.850000 1182.000000 82.150000 ;
        RECT 1172.000000 101.850000 1182.000000 102.150000 ;
        RECT 1172.000000 85.850000 1182.000000 86.150000 ;
        RECT 1172.000000 89.850000 1182.000000 90.150000 ;
        RECT 1172.000000 93.850000 1182.000000 94.150000 ;
        RECT 1172.000000 97.850000 1182.000000 98.150000 ;
        RECT 1172.000000 117.850000 1182.000000 118.150000 ;
        RECT 1172.000000 113.850000 1182.000000 114.150000 ;
        RECT 1172.000000 105.850000 1182.000000 106.150000 ;
        RECT 1172.000000 109.850000 1182.000000 110.150000 ;
        RECT 1151.000000 133.850000 1156.000000 134.150000 ;
        RECT 1172.000000 129.850000 1182.000000 130.150000 ;
        RECT 1172.000000 125.850000 1182.000000 126.150000 ;
        RECT 1172.000000 121.850000 1182.000000 122.150000 ;
        RECT 1172.000000 133.850000 1182.000000 134.150000 ;
        RECT 1172.000000 137.850000 1182.000000 138.150000 ;
        RECT 1172.000000 141.850000 1182.000000 142.150000 ;
        RECT 1172.000000 145.850000 1182.000000 146.150000 ;
        RECT 1172.000000 149.850000 1182.000000 150.150000 ;
        RECT 1172.000000 153.850000 1182.000000 154.150000 ;
        RECT 1172.000000 165.850000 1182.000000 166.150000 ;
        RECT 1172.000000 161.850000 1182.000000 162.150000 ;
        RECT 1172.000000 157.850000 1182.000000 158.150000 ;
        RECT 1172.000000 169.850000 1182.000000 170.150000 ;
        RECT 1172.000000 173.850000 1182.000000 174.150000 ;
        RECT 1172.000000 177.850000 1182.000000 178.150000 ;
        RECT 1172.000000 181.850000 1182.000000 182.150000 ;
        RECT 1172.000000 185.850000 1182.000000 186.150000 ;
        RECT 1172.000000 189.850000 1182.000000 190.150000 ;
        RECT 1172.000000 193.850000 1182.000000 194.150000 ;
        RECT 901.000000 261.850000 906.000000 262.150000 ;
        RECT 901.000000 265.850000 906.000000 266.150000 ;
        RECT 951.000000 265.850000 956.000000 266.150000 ;
        RECT 951.000000 261.850000 956.000000 262.150000 ;
        RECT 1001.000000 261.850000 1006.000000 262.150000 ;
        RECT 1001.000000 265.850000 1006.000000 266.150000 ;
        RECT 951.000000 305.850000 956.000000 306.150000 ;
        RECT 901.000000 305.850000 906.000000 306.150000 ;
        RECT 901.000000 285.850000 906.000000 286.150000 ;
        RECT 901.000000 281.850000 906.000000 282.150000 ;
        RECT 901.000000 269.850000 906.000000 270.150000 ;
        RECT 901.000000 273.850000 906.000000 274.150000 ;
        RECT 901.000000 277.850000 906.000000 278.150000 ;
        RECT 901.000000 289.850000 906.000000 290.150000 ;
        RECT 901.000000 293.850000 906.000000 294.150000 ;
        RECT 901.000000 297.850000 906.000000 298.150000 ;
        RECT 901.000000 301.850000 906.000000 302.150000 ;
        RECT 951.000000 269.850000 956.000000 270.150000 ;
        RECT 951.000000 273.850000 956.000000 274.150000 ;
        RECT 951.000000 277.850000 956.000000 278.150000 ;
        RECT 951.000000 281.850000 956.000000 282.150000 ;
        RECT 951.000000 285.850000 956.000000 286.150000 ;
        RECT 951.000000 301.850000 956.000000 302.150000 ;
        RECT 951.000000 297.850000 956.000000 298.150000 ;
        RECT 951.000000 293.850000 956.000000 294.150000 ;
        RECT 951.000000 289.850000 956.000000 290.150000 ;
        RECT 901.000000 321.850000 906.000000 322.150000 ;
        RECT 901.000000 309.850000 906.000000 310.150000 ;
        RECT 901.000000 313.850000 906.000000 314.150000 ;
        RECT 901.000000 317.850000 906.000000 318.150000 ;
        RECT 901.000000 325.850000 906.000000 326.150000 ;
        RECT 901.000000 329.850000 906.000000 330.150000 ;
        RECT 901.000000 333.850000 906.000000 334.150000 ;
        RECT 901.000000 337.850000 906.000000 338.150000 ;
        RECT 901.000000 341.850000 906.000000 342.150000 ;
        RECT 951.000000 313.850000 956.000000 314.150000 ;
        RECT 951.000000 309.850000 956.000000 310.150000 ;
        RECT 951.000000 317.850000 956.000000 318.150000 ;
        RECT 951.000000 321.850000 956.000000 322.150000 ;
        RECT 951.000000 325.850000 956.000000 326.150000 ;
        RECT 951.000000 329.850000 956.000000 330.150000 ;
        RECT 951.000000 333.850000 956.000000 334.150000 ;
        RECT 951.000000 337.850000 956.000000 338.150000 ;
        RECT 951.000000 341.850000 956.000000 342.150000 ;
        RECT 1001.000000 305.850000 1006.000000 306.150000 ;
        RECT 1001.000000 277.850000 1006.000000 278.150000 ;
        RECT 1001.000000 269.850000 1006.000000 270.150000 ;
        RECT 1001.000000 273.850000 1006.000000 274.150000 ;
        RECT 1001.000000 281.850000 1006.000000 282.150000 ;
        RECT 1001.000000 285.850000 1006.000000 286.150000 ;
        RECT 1001.000000 289.850000 1006.000000 290.150000 ;
        RECT 1001.000000 293.850000 1006.000000 294.150000 ;
        RECT 1001.000000 301.850000 1006.000000 302.150000 ;
        RECT 1001.000000 297.850000 1006.000000 298.150000 ;
        RECT 1001.000000 313.850000 1006.000000 314.150000 ;
        RECT 1001.000000 309.850000 1006.000000 310.150000 ;
        RECT 1001.000000 317.850000 1006.000000 318.150000 ;
        RECT 1001.000000 321.850000 1006.000000 322.150000 ;
        RECT 1001.000000 329.850000 1006.000000 330.150000 ;
        RECT 1001.000000 325.850000 1006.000000 326.150000 ;
        RECT 1001.000000 333.850000 1006.000000 334.150000 ;
        RECT 1001.000000 337.850000 1006.000000 338.150000 ;
        RECT 1001.000000 341.850000 1006.000000 342.150000 ;
        RECT 1051.000000 261.850000 1056.000000 262.150000 ;
        RECT 1051.000000 265.850000 1056.000000 266.150000 ;
        RECT 1101.000000 265.850000 1106.000000 266.150000 ;
        RECT 1101.000000 261.850000 1106.000000 262.150000 ;
        RECT 1172.000000 197.850000 1182.000000 198.150000 ;
        RECT 1172.000000 201.850000 1182.000000 202.150000 ;
        RECT 1172.000000 205.850000 1182.000000 206.150000 ;
        RECT 1172.000000 209.850000 1182.000000 210.150000 ;
        RECT 1172.000000 221.850000 1182.000000 222.150000 ;
        RECT 1172.000000 217.850000 1182.000000 218.150000 ;
        RECT 1172.000000 213.850000 1182.000000 214.150000 ;
        RECT 1172.000000 225.850000 1182.000000 226.150000 ;
        RECT 1172.000000 229.850000 1182.000000 230.150000 ;
        RECT 1172.000000 237.850000 1182.000000 238.150000 ;
        RECT 1172.000000 233.850000 1182.000000 234.150000 ;
        RECT 1172.000000 241.850000 1182.000000 242.150000 ;
        RECT 1172.000000 245.850000 1182.000000 246.150000 ;
        RECT 1172.000000 249.850000 1182.000000 250.150000 ;
        RECT 1151.000000 257.850000 1156.000000 258.150000 ;
        RECT 1151.000000 265.850000 1156.000000 266.150000 ;
        RECT 1151.000000 261.850000 1156.000000 262.150000 ;
        RECT 1172.000000 265.850000 1182.000000 266.150000 ;
        RECT 1172.000000 253.850000 1182.000000 254.150000 ;
        RECT 1172.000000 257.850000 1182.000000 258.150000 ;
        RECT 1172.000000 261.850000 1182.000000 262.150000 ;
        RECT 1101.000000 305.850000 1106.000000 306.150000 ;
        RECT 1051.000000 305.850000 1056.000000 306.150000 ;
        RECT 1051.000000 285.850000 1056.000000 286.150000 ;
        RECT 1051.000000 281.850000 1056.000000 282.150000 ;
        RECT 1051.000000 273.850000 1056.000000 274.150000 ;
        RECT 1051.000000 269.850000 1056.000000 270.150000 ;
        RECT 1051.000000 277.850000 1056.000000 278.150000 ;
        RECT 1051.000000 289.850000 1056.000000 290.150000 ;
        RECT 1051.000000 293.850000 1056.000000 294.150000 ;
        RECT 1051.000000 297.850000 1056.000000 298.150000 ;
        RECT 1051.000000 301.850000 1056.000000 302.150000 ;
        RECT 1101.000000 269.850000 1106.000000 270.150000 ;
        RECT 1101.000000 273.850000 1106.000000 274.150000 ;
        RECT 1101.000000 277.850000 1106.000000 278.150000 ;
        RECT 1101.000000 281.850000 1106.000000 282.150000 ;
        RECT 1101.000000 285.850000 1106.000000 286.150000 ;
        RECT 1101.000000 301.850000 1106.000000 302.150000 ;
        RECT 1101.000000 297.850000 1106.000000 298.150000 ;
        RECT 1101.000000 293.850000 1106.000000 294.150000 ;
        RECT 1101.000000 289.850000 1106.000000 290.150000 ;
        RECT 1051.000000 321.850000 1056.000000 322.150000 ;
        RECT 1051.000000 309.850000 1056.000000 310.150000 ;
        RECT 1051.000000 313.850000 1056.000000 314.150000 ;
        RECT 1051.000000 317.850000 1056.000000 318.150000 ;
        RECT 1051.000000 325.850000 1056.000000 326.150000 ;
        RECT 1051.000000 329.850000 1056.000000 330.150000 ;
        RECT 1051.000000 333.850000 1056.000000 334.150000 ;
        RECT 1051.000000 337.850000 1056.000000 338.150000 ;
        RECT 1051.000000 341.850000 1056.000000 342.150000 ;
        RECT 1101.000000 313.850000 1106.000000 314.150000 ;
        RECT 1101.000000 309.850000 1106.000000 310.150000 ;
        RECT 1101.000000 317.850000 1106.000000 318.150000 ;
        RECT 1101.000000 321.850000 1106.000000 322.150000 ;
        RECT 1101.000000 325.850000 1106.000000 326.150000 ;
        RECT 1101.000000 329.850000 1106.000000 330.150000 ;
        RECT 1101.000000 333.850000 1106.000000 334.150000 ;
        RECT 1101.000000 337.850000 1106.000000 338.150000 ;
        RECT 1101.000000 341.850000 1106.000000 342.150000 ;
        RECT 1151.000000 305.850000 1156.000000 306.150000 ;
        RECT 1172.000000 305.850000 1182.000000 306.150000 ;
        RECT 1151.000000 277.850000 1156.000000 278.150000 ;
        RECT 1151.000000 269.850000 1156.000000 270.150000 ;
        RECT 1151.000000 273.850000 1156.000000 274.150000 ;
        RECT 1151.000000 281.850000 1156.000000 282.150000 ;
        RECT 1151.000000 285.850000 1156.000000 286.150000 ;
        RECT 1172.000000 277.850000 1182.000000 278.150000 ;
        RECT 1172.000000 269.850000 1182.000000 270.150000 ;
        RECT 1172.000000 273.850000 1182.000000 274.150000 ;
        RECT 1172.000000 281.850000 1182.000000 282.150000 ;
        RECT 1172.000000 285.850000 1182.000000 286.150000 ;
        RECT 1151.000000 301.850000 1156.000000 302.150000 ;
        RECT 1151.000000 297.850000 1156.000000 298.150000 ;
        RECT 1151.000000 289.850000 1156.000000 290.150000 ;
        RECT 1151.000000 293.850000 1156.000000 294.150000 ;
        RECT 1172.000000 301.850000 1182.000000 302.150000 ;
        RECT 1172.000000 289.850000 1182.000000 290.150000 ;
        RECT 1172.000000 293.850000 1182.000000 294.150000 ;
        RECT 1172.000000 297.850000 1182.000000 298.150000 ;
        RECT 1151.000000 321.850000 1156.000000 322.150000 ;
        RECT 1151.000000 317.850000 1156.000000 318.150000 ;
        RECT 1151.000000 309.850000 1156.000000 310.150000 ;
        RECT 1151.000000 313.850000 1156.000000 314.150000 ;
        RECT 1172.000000 321.850000 1182.000000 322.150000 ;
        RECT 1172.000000 309.850000 1182.000000 310.150000 ;
        RECT 1172.000000 313.850000 1182.000000 314.150000 ;
        RECT 1172.000000 317.850000 1182.000000 318.150000 ;
        RECT 1151.000000 329.850000 1156.000000 330.150000 ;
        RECT 1151.000000 325.850000 1156.000000 326.150000 ;
        RECT 1151.000000 333.850000 1156.000000 334.150000 ;
        RECT 1151.000000 337.850000 1156.000000 338.150000 ;
        RECT 1151.000000 341.850000 1156.000000 342.150000 ;
        RECT 1172.000000 329.850000 1182.000000 330.150000 ;
        RECT 1172.000000 325.850000 1182.000000 326.150000 ;
        RECT 1172.000000 333.850000 1182.000000 334.150000 ;
        RECT 1172.000000 337.850000 1182.000000 338.150000 ;
        RECT 1172.000000 341.850000 1182.000000 342.150000 ;
        RECT 4.000000 357.850000 14.000000 358.150000 ;
        RECT 4.000000 353.850000 14.000000 354.150000 ;
        RECT 4.000000 345.850000 14.000000 346.150000 ;
        RECT 4.000000 349.850000 14.000000 350.150000 ;
        RECT 4.000000 369.850000 14.000000 370.150000 ;
        RECT 4.000000 365.850000 14.000000 366.150000 ;
        RECT 4.000000 361.850000 14.000000 362.150000 ;
        RECT 4.000000 377.850000 14.000000 378.150000 ;
        RECT 4.000000 373.850000 14.000000 374.150000 ;
        RECT 51.000000 354.445000 56.000000 354.745000 ;
        RECT 51.000000 345.850000 56.000000 346.150000 ;
        RECT 51.000000 369.850000 56.000000 370.150000 ;
        RECT 51.000000 365.850000 56.000000 366.150000 ;
        RECT 51.000000 361.850000 56.000000 362.150000 ;
        RECT 51.000000 373.850000 56.000000 374.150000 ;
        RECT 51.000000 377.850000 56.000000 378.150000 ;
        RECT 4.000000 397.850000 14.000000 398.150000 ;
        RECT 4.000000 393.850000 14.000000 394.150000 ;
        RECT 4.000000 389.850000 14.000000 390.150000 ;
        RECT 4.000000 381.850000 14.000000 382.150000 ;
        RECT 4.000000 385.850000 14.000000 386.150000 ;
        RECT 4.000000 401.850000 14.000000 402.150000 ;
        RECT 4.000000 405.850000 14.000000 406.150000 ;
        RECT 4.000000 409.850000 14.000000 410.150000 ;
        RECT 4.000000 413.850000 14.000000 414.150000 ;
        RECT 51.000000 385.850000 56.000000 386.150000 ;
        RECT 51.000000 381.850000 56.000000 382.150000 ;
        RECT 51.000000 389.850000 56.000000 390.150000 ;
        RECT 51.000000 393.850000 56.000000 394.150000 ;
        RECT 51.000000 397.850000 56.000000 398.150000 ;
        RECT 51.000000 413.850000 56.000000 414.150000 ;
        RECT 51.000000 409.850000 56.000000 410.150000 ;
        RECT 51.000000 405.850000 56.000000 406.150000 ;
        RECT 51.000000 401.850000 56.000000 402.150000 ;
        RECT 101.000000 345.850000 106.000000 346.150000 ;
        RECT 101.000000 349.850000 106.000000 350.150000 ;
        RECT 101.000000 353.850000 106.000000 354.150000 ;
        RECT 101.000000 357.850000 106.000000 358.150000 ;
        RECT 101.000000 361.850000 106.000000 362.150000 ;
        RECT 101.000000 365.850000 106.000000 366.150000 ;
        RECT 101.000000 369.850000 106.000000 370.150000 ;
        RECT 101.000000 373.850000 106.000000 374.150000 ;
        RECT 101.000000 377.850000 106.000000 378.150000 ;
        RECT 101.000000 381.850000 106.000000 382.150000 ;
        RECT 101.000000 385.850000 106.000000 386.150000 ;
        RECT 101.000000 389.850000 106.000000 390.150000 ;
        RECT 101.000000 393.850000 106.000000 394.150000 ;
        RECT 101.000000 397.850000 106.000000 398.150000 ;
        RECT 101.000000 413.850000 106.000000 414.150000 ;
        RECT 101.000000 409.850000 106.000000 410.150000 ;
        RECT 101.000000 405.850000 106.000000 406.150000 ;
        RECT 101.000000 401.850000 106.000000 402.150000 ;
        RECT 4.000000 433.850000 14.000000 434.150000 ;
        RECT 4.000000 429.850000 14.000000 430.150000 ;
        RECT 4.000000 417.850000 14.000000 418.150000 ;
        RECT 4.000000 421.850000 14.000000 422.150000 ;
        RECT 4.000000 425.850000 14.000000 426.150000 ;
        RECT 4.000000 437.850000 14.000000 438.150000 ;
        RECT 4.000000 441.850000 14.000000 442.150000 ;
        RECT 4.000000 445.850000 14.000000 446.150000 ;
        RECT 4.000000 449.850000 14.000000 450.150000 ;
        RECT 4.000000 453.850000 14.000000 454.150000 ;
        RECT 51.000000 417.850000 56.000000 418.150000 ;
        RECT 51.000000 421.850000 56.000000 422.150000 ;
        RECT 51.000000 425.850000 56.000000 426.150000 ;
        RECT 51.000000 429.850000 56.000000 430.150000 ;
        RECT 51.000000 433.850000 56.000000 434.150000 ;
        RECT 51.000000 453.850000 56.000000 454.150000 ;
        RECT 51.000000 449.850000 56.000000 450.150000 ;
        RECT 51.000000 445.850000 56.000000 446.150000 ;
        RECT 51.000000 441.850000 56.000000 442.150000 ;
        RECT 51.000000 437.850000 56.000000 438.150000 ;
        RECT 4.000000 469.850000 14.000000 470.150000 ;
        RECT 4.000000 457.850000 14.000000 458.150000 ;
        RECT 4.000000 461.850000 14.000000 462.150000 ;
        RECT 4.000000 465.850000 14.000000 466.150000 ;
        RECT 4.000000 473.850000 14.000000 474.150000 ;
        RECT 4.000000 477.850000 14.000000 478.150000 ;
        RECT 4.000000 481.850000 14.000000 482.150000 ;
        RECT 4.000000 485.850000 14.000000 486.150000 ;
        RECT 4.000000 489.850000 14.000000 490.150000 ;
        RECT 51.000000 461.850000 56.000000 462.150000 ;
        RECT 51.000000 457.850000 56.000000 458.150000 ;
        RECT 51.000000 465.850000 56.000000 466.150000 ;
        RECT 51.000000 469.850000 56.000000 470.150000 ;
        RECT 51.000000 489.850000 56.000000 490.150000 ;
        RECT 51.000000 485.850000 56.000000 486.150000 ;
        RECT 51.000000 481.850000 56.000000 482.150000 ;
        RECT 51.000000 477.850000 56.000000 478.150000 ;
        RECT 51.000000 473.850000 56.000000 474.150000 ;
        RECT 101.000000 417.850000 106.000000 418.150000 ;
        RECT 101.000000 421.850000 106.000000 422.150000 ;
        RECT 101.000000 425.850000 106.000000 426.150000 ;
        RECT 101.000000 429.850000 106.000000 430.150000 ;
        RECT 101.000000 433.850000 106.000000 434.150000 ;
        RECT 101.000000 437.850000 106.000000 438.150000 ;
        RECT 101.000000 441.850000 106.000000 442.150000 ;
        RECT 101.000000 445.850000 106.000000 446.150000 ;
        RECT 101.000000 449.850000 106.000000 450.150000 ;
        RECT 101.000000 453.850000 106.000000 454.150000 ;
        RECT 101.000000 469.850000 106.000000 470.150000 ;
        RECT 101.000000 465.850000 106.000000 466.150000 ;
        RECT 101.000000 461.850000 106.000000 462.150000 ;
        RECT 101.000000 457.850000 106.000000 458.150000 ;
        RECT 101.000000 473.850000 106.000000 474.150000 ;
        RECT 101.000000 477.850000 106.000000 478.150000 ;
        RECT 101.000000 481.850000 106.000000 482.150000 ;
        RECT 101.000000 485.850000 106.000000 486.150000 ;
        RECT 101.000000 489.850000 106.000000 490.150000 ;
        RECT 151.000000 349.850000 156.000000 350.150000 ;
        RECT 151.000000 345.850000 156.000000 346.150000 ;
        RECT 151.000000 353.850000 156.000000 354.150000 ;
        RECT 151.000000 357.850000 156.000000 358.150000 ;
        RECT 151.000000 361.850000 156.000000 362.150000 ;
        RECT 151.000000 365.850000 156.000000 366.150000 ;
        RECT 151.000000 369.850000 156.000000 370.150000 ;
        RECT 151.000000 377.850000 156.000000 378.150000 ;
        RECT 151.000000 373.850000 156.000000 374.150000 ;
        RECT 201.000000 349.850000 206.000000 350.150000 ;
        RECT 201.000000 345.850000 206.000000 346.150000 ;
        RECT 201.000000 353.850000 206.000000 354.150000 ;
        RECT 201.000000 357.850000 206.000000 358.150000 ;
        RECT 201.000000 361.850000 206.000000 362.150000 ;
        RECT 201.000000 365.850000 206.000000 366.150000 ;
        RECT 201.000000 369.850000 206.000000 370.150000 ;
        RECT 201.000000 373.850000 206.000000 374.150000 ;
        RECT 201.000000 377.850000 206.000000 378.150000 ;
        RECT 151.000000 385.850000 156.000000 386.150000 ;
        RECT 151.000000 381.850000 156.000000 382.150000 ;
        RECT 151.000000 393.850000 156.000000 394.150000 ;
        RECT 151.000000 389.850000 156.000000 390.150000 ;
        RECT 151.000000 397.850000 156.000000 398.150000 ;
        RECT 151.000000 401.850000 156.000000 402.150000 ;
        RECT 201.000000 381.850000 206.000000 382.150000 ;
        RECT 201.000000 385.850000 206.000000 386.150000 ;
        RECT 201.000000 397.850000 206.000000 398.150000 ;
        RECT 201.000000 393.850000 206.000000 394.150000 ;
        RECT 201.000000 389.850000 206.000000 390.150000 ;
        RECT 201.000000 413.850000 206.000000 414.150000 ;
        RECT 201.000000 409.850000 206.000000 410.150000 ;
        RECT 201.000000 405.850000 206.000000 406.150000 ;
        RECT 201.000000 401.850000 206.000000 402.150000 ;
        RECT 251.000000 345.850000 256.000000 346.150000 ;
        RECT 251.000000 349.850000 256.000000 350.150000 ;
        RECT 251.000000 353.850000 256.000000 354.150000 ;
        RECT 251.000000 357.850000 256.000000 358.150000 ;
        RECT 251.000000 369.850000 256.000000 370.150000 ;
        RECT 251.000000 365.850000 256.000000 366.150000 ;
        RECT 251.000000 361.850000 256.000000 362.150000 ;
        RECT 251.000000 373.850000 256.000000 374.150000 ;
        RECT 251.000000 377.850000 256.000000 378.150000 ;
        RECT 251.000000 381.850000 256.000000 382.150000 ;
        RECT 251.000000 385.850000 256.000000 386.150000 ;
        RECT 251.000000 397.850000 256.000000 398.150000 ;
        RECT 251.000000 393.850000 256.000000 394.150000 ;
        RECT 251.000000 389.850000 256.000000 390.150000 ;
        RECT 251.000000 401.850000 256.000000 402.150000 ;
        RECT 151.000000 453.850000 156.000000 454.150000 ;
        RECT 201.000000 425.850000 206.000000 426.150000 ;
        RECT 201.000000 421.850000 206.000000 422.150000 ;
        RECT 201.000000 417.850000 206.000000 418.150000 ;
        RECT 201.000000 429.850000 206.000000 430.150000 ;
        RECT 201.000000 433.850000 206.000000 434.150000 ;
        RECT 201.000000 453.850000 206.000000 454.150000 ;
        RECT 201.000000 449.850000 206.000000 450.150000 ;
        RECT 201.000000 445.850000 206.000000 446.150000 ;
        RECT 201.000000 441.850000 206.000000 442.150000 ;
        RECT 201.000000 437.850000 206.000000 438.150000 ;
        RECT 151.000000 461.850000 156.000000 462.150000 ;
        RECT 151.000000 457.850000 156.000000 458.150000 ;
        RECT 151.000000 469.850000 156.000000 470.150000 ;
        RECT 151.000000 465.850000 156.000000 466.150000 ;
        RECT 151.000000 481.850000 156.000000 482.150000 ;
        RECT 151.000000 477.850000 156.000000 478.150000 ;
        RECT 151.000000 473.850000 156.000000 474.150000 ;
        RECT 151.000000 489.850000 156.000000 490.150000 ;
        RECT 151.000000 485.850000 156.000000 486.150000 ;
        RECT 201.000000 461.850000 206.000000 462.150000 ;
        RECT 201.000000 457.850000 206.000000 458.150000 ;
        RECT 201.000000 465.850000 206.000000 466.150000 ;
        RECT 201.000000 469.850000 206.000000 470.150000 ;
        RECT 201.000000 489.850000 206.000000 490.150000 ;
        RECT 201.000000 485.850000 206.000000 486.150000 ;
        RECT 201.000000 481.850000 206.000000 482.150000 ;
        RECT 201.000000 477.850000 206.000000 478.150000 ;
        RECT 201.000000 473.850000 206.000000 474.150000 ;
        RECT 251.000000 453.850000 256.000000 454.150000 ;
        RECT 251.000000 457.850000 256.000000 458.150000 ;
        RECT 251.000000 461.850000 256.000000 462.150000 ;
        RECT 251.000000 465.850000 256.000000 466.150000 ;
        RECT 251.000000 469.850000 256.000000 470.150000 ;
        RECT 251.000000 481.850000 256.000000 482.150000 ;
        RECT 251.000000 473.850000 256.000000 474.150000 ;
        RECT 251.000000 477.850000 256.000000 478.150000 ;
        RECT 251.000000 485.850000 256.000000 486.150000 ;
        RECT 251.000000 489.850000 256.000000 490.150000 ;
        RECT 4.000000 505.850000 14.000000 506.150000 ;
        RECT 4.000000 497.850000 14.000000 498.150000 ;
        RECT 4.000000 493.850000 14.000000 494.150000 ;
        RECT 4.000000 501.850000 14.000000 502.150000 ;
        RECT 4.000000 513.850000 14.000000 514.150000 ;
        RECT 4.000000 509.850000 14.000000 510.150000 ;
        RECT 51.000000 493.850000 56.000000 494.150000 ;
        RECT 51.000000 497.850000 56.000000 498.150000 ;
        RECT 51.000000 501.850000 56.000000 502.150000 ;
        RECT 51.000000 505.850000 56.000000 506.150000 ;
        RECT 51.000000 513.850000 56.000000 514.150000 ;
        RECT 51.000000 509.850000 56.000000 510.150000 ;
        RECT 101.000000 505.850000 106.000000 506.150000 ;
        RECT 101.000000 501.850000 106.000000 502.150000 ;
        RECT 101.000000 497.850000 106.000000 498.150000 ;
        RECT 101.000000 493.850000 106.000000 494.150000 ;
        RECT 101.000000 513.850000 106.000000 514.150000 ;
        RECT 101.000000 509.850000 106.000000 510.150000 ;
        RECT 151.000000 493.850000 156.000000 494.150000 ;
        RECT 151.000000 497.850000 156.000000 498.150000 ;
        RECT 151.000000 501.850000 156.000000 502.150000 ;
        RECT 151.000000 505.850000 156.000000 506.150000 ;
        RECT 151.000000 513.850000 156.000000 514.150000 ;
        RECT 151.000000 509.850000 156.000000 510.150000 ;
        RECT 201.000000 497.850000 206.000000 498.150000 ;
        RECT 201.000000 493.850000 206.000000 494.150000 ;
        RECT 201.000000 501.850000 206.000000 502.150000 ;
        RECT 201.000000 505.850000 206.000000 506.150000 ;
        RECT 201.000000 513.850000 206.000000 514.150000 ;
        RECT 201.000000 509.850000 206.000000 510.150000 ;
        RECT 251.000000 493.850000 256.000000 494.150000 ;
        RECT 251.000000 497.850000 256.000000 498.150000 ;
        RECT 251.000000 505.850000 256.000000 506.150000 ;
        RECT 251.000000 501.850000 256.000000 502.150000 ;
        RECT 251.000000 513.850000 256.000000 514.150000 ;
        RECT 251.000000 509.850000 256.000000 510.150000 ;
        RECT 301.000000 345.850000 306.000000 346.150000 ;
        RECT 301.000000 349.850000 306.000000 350.150000 ;
        RECT 301.000000 353.850000 306.000000 354.150000 ;
        RECT 301.000000 357.850000 306.000000 358.150000 ;
        RECT 301.000000 369.850000 306.000000 370.150000 ;
        RECT 301.000000 365.850000 306.000000 366.150000 ;
        RECT 301.000000 361.850000 306.000000 362.150000 ;
        RECT 301.000000 377.850000 306.000000 378.150000 ;
        RECT 301.000000 373.850000 306.000000 374.150000 ;
        RECT 351.000000 345.850000 356.000000 346.150000 ;
        RECT 351.000000 349.850000 356.000000 350.150000 ;
        RECT 351.000000 353.850000 356.000000 354.150000 ;
        RECT 351.000000 357.850000 356.000000 358.150000 ;
        RECT 351.000000 361.850000 356.000000 362.150000 ;
        RECT 351.000000 365.850000 356.000000 366.150000 ;
        RECT 351.000000 369.850000 356.000000 370.150000 ;
        RECT 351.000000 373.850000 356.000000 374.150000 ;
        RECT 351.000000 377.850000 356.000000 378.150000 ;
        RECT 301.000000 385.850000 306.000000 386.150000 ;
        RECT 301.000000 381.850000 306.000000 382.150000 ;
        RECT 301.000000 389.850000 306.000000 390.150000 ;
        RECT 301.000000 393.850000 306.000000 394.150000 ;
        RECT 301.000000 397.850000 306.000000 398.150000 ;
        RECT 301.000000 405.850000 306.000000 406.150000 ;
        RECT 301.000000 401.850000 306.000000 402.150000 ;
        RECT 301.000000 409.850000 306.000000 410.150000 ;
        RECT 301.000000 413.850000 306.000000 414.150000 ;
        RECT 351.000000 381.850000 356.000000 382.150000 ;
        RECT 351.000000 385.850000 356.000000 386.150000 ;
        RECT 351.000000 397.850000 356.000000 398.150000 ;
        RECT 351.000000 393.850000 356.000000 394.150000 ;
        RECT 351.000000 389.850000 356.000000 390.150000 ;
        RECT 351.000000 413.850000 356.000000 414.150000 ;
        RECT 351.000000 409.850000 356.000000 410.150000 ;
        RECT 351.000000 405.850000 356.000000 406.150000 ;
        RECT 351.000000 401.850000 356.000000 402.150000 ;
        RECT 401.000000 345.850000 406.000000 346.150000 ;
        RECT 401.000000 349.850000 406.000000 350.150000 ;
        RECT 401.000000 353.850000 406.000000 354.150000 ;
        RECT 401.000000 357.850000 406.000000 358.150000 ;
        RECT 401.000000 365.850000 406.000000 366.150000 ;
        RECT 401.000000 361.850000 406.000000 362.150000 ;
        RECT 401.000000 369.850000 406.000000 370.150000 ;
        RECT 401.000000 373.850000 406.000000 374.150000 ;
        RECT 401.000000 377.850000 406.000000 378.150000 ;
        RECT 401.000000 381.850000 406.000000 382.150000 ;
        RECT 401.000000 385.850000 406.000000 386.150000 ;
        RECT 401.000000 393.850000 406.000000 394.150000 ;
        RECT 401.000000 389.850000 406.000000 390.150000 ;
        RECT 401.000000 397.850000 406.000000 398.150000 ;
        RECT 401.000000 401.850000 406.000000 402.150000 ;
        RECT 401.000000 405.850000 406.000000 406.150000 ;
        RECT 401.000000 409.850000 406.000000 410.150000 ;
        RECT 401.000000 413.850000 406.000000 414.150000 ;
        RECT 301.000000 425.850000 306.000000 426.150000 ;
        RECT 301.000000 417.850000 306.000000 418.150000 ;
        RECT 301.000000 421.850000 306.000000 422.150000 ;
        RECT 301.000000 429.850000 306.000000 430.150000 ;
        RECT 301.000000 433.850000 306.000000 434.150000 ;
        RECT 301.000000 441.850000 306.000000 442.150000 ;
        RECT 301.000000 437.850000 306.000000 438.150000 ;
        RECT 301.000000 453.850000 306.000000 454.150000 ;
        RECT 301.000000 449.850000 306.000000 450.150000 ;
        RECT 301.000000 445.850000 306.000000 446.150000 ;
        RECT 351.000000 425.850000 356.000000 426.150000 ;
        RECT 351.000000 421.850000 356.000000 422.150000 ;
        RECT 351.000000 417.850000 356.000000 418.150000 ;
        RECT 351.000000 433.850000 356.000000 434.150000 ;
        RECT 351.000000 429.850000 356.000000 430.150000 ;
        RECT 351.000000 453.850000 356.000000 454.150000 ;
        RECT 351.000000 449.850000 356.000000 450.150000 ;
        RECT 351.000000 445.850000 356.000000 446.150000 ;
        RECT 351.000000 441.850000 356.000000 442.150000 ;
        RECT 351.000000 437.850000 356.000000 438.150000 ;
        RECT 301.000000 457.850000 306.000000 458.150000 ;
        RECT 301.000000 461.850000 306.000000 462.150000 ;
        RECT 301.000000 465.850000 306.000000 466.150000 ;
        RECT 301.000000 469.850000 306.000000 470.150000 ;
        RECT 301.000000 481.850000 306.000000 482.150000 ;
        RECT 301.000000 477.850000 306.000000 478.150000 ;
        RECT 301.000000 473.850000 306.000000 474.150000 ;
        RECT 301.000000 489.850000 306.000000 490.150000 ;
        RECT 301.000000 485.850000 306.000000 486.150000 ;
        RECT 351.000000 461.850000 356.000000 462.150000 ;
        RECT 351.000000 457.850000 356.000000 458.150000 ;
        RECT 351.000000 465.850000 356.000000 466.150000 ;
        RECT 351.000000 469.850000 356.000000 470.150000 ;
        RECT 351.000000 481.850000 356.000000 482.150000 ;
        RECT 351.000000 473.850000 356.000000 474.150000 ;
        RECT 351.000000 477.850000 356.000000 478.150000 ;
        RECT 351.000000 485.850000 356.000000 486.150000 ;
        RECT 351.000000 489.850000 356.000000 490.150000 ;
        RECT 401.000000 417.850000 406.000000 418.150000 ;
        RECT 401.000000 421.850000 406.000000 422.150000 ;
        RECT 401.000000 425.850000 406.000000 426.150000 ;
        RECT 401.000000 433.850000 406.000000 434.150000 ;
        RECT 401.000000 429.850000 406.000000 430.150000 ;
        RECT 401.000000 441.850000 406.000000 442.150000 ;
        RECT 401.000000 437.850000 406.000000 438.150000 ;
        RECT 401.000000 445.850000 406.000000 446.150000 ;
        RECT 401.000000 453.850000 406.000000 454.150000 ;
        RECT 401.000000 449.850000 406.000000 450.150000 ;
        RECT 401.000000 457.850000 406.000000 458.150000 ;
        RECT 401.000000 461.850000 406.000000 462.150000 ;
        RECT 401.000000 465.850000 406.000000 466.150000 ;
        RECT 401.000000 469.850000 406.000000 470.150000 ;
        RECT 401.000000 481.850000 406.000000 482.150000 ;
        RECT 401.000000 473.850000 406.000000 474.150000 ;
        RECT 401.000000 477.850000 406.000000 478.150000 ;
        RECT 401.000000 485.850000 406.000000 486.150000 ;
        RECT 401.000000 489.850000 406.000000 490.150000 ;
        RECT 451.000000 345.850000 456.000000 346.150000 ;
        RECT 451.000000 366.105000 456.000000 367.105000 ;
        RECT 451.000000 369.850000 456.000000 370.150000 ;
        RECT 451.000000 373.850000 456.000000 374.150000 ;
        RECT 451.000000 377.850000 456.000000 378.150000 ;
        RECT 501.000000 345.850000 506.000000 346.150000 ;
        RECT 501.000000 349.850000 506.000000 350.150000 ;
        RECT 501.000000 353.850000 506.000000 354.150000 ;
        RECT 501.000000 357.850000 506.000000 358.150000 ;
        RECT 501.000000 365.850000 506.000000 366.150000 ;
        RECT 501.000000 361.850000 506.000000 362.150000 ;
        RECT 501.000000 369.850000 506.000000 370.150000 ;
        RECT 501.000000 377.850000 506.000000 378.150000 ;
        RECT 501.000000 373.850000 506.000000 374.150000 ;
        RECT 451.000000 381.850000 456.000000 382.150000 ;
        RECT 451.000000 385.850000 456.000000 386.150000 ;
        RECT 451.000000 397.850000 456.000000 398.150000 ;
        RECT 451.000000 393.850000 456.000000 394.150000 ;
        RECT 451.000000 389.850000 456.000000 390.150000 ;
        RECT 451.000000 416.105000 456.000000 417.105000 ;
        RECT 501.000000 385.850000 506.000000 386.150000 ;
        RECT 501.000000 381.850000 506.000000 382.150000 ;
        RECT 501.000000 393.850000 506.000000 394.150000 ;
        RECT 501.000000 389.850000 506.000000 390.150000 ;
        RECT 501.000000 397.850000 506.000000 398.150000 ;
        RECT 501.000000 401.850000 506.000000 402.150000 ;
        RECT 501.000000 405.850000 506.000000 406.150000 ;
        RECT 501.000000 409.850000 506.000000 410.150000 ;
        RECT 501.000000 413.850000 506.000000 414.150000 ;
        RECT 551.000000 357.850000 556.000000 358.150000 ;
        RECT 551.000000 353.850000 556.000000 354.150000 ;
        RECT 551.000000 349.850000 556.000000 350.150000 ;
        RECT 551.000000 345.850000 556.000000 346.150000 ;
        RECT 551.000000 361.850000 556.000000 362.150000 ;
        RECT 551.000000 365.850000 556.000000 366.150000 ;
        RECT 551.000000 369.850000 556.000000 370.150000 ;
        RECT 551.000000 373.850000 556.000000 374.150000 ;
        RECT 551.000000 377.850000 556.000000 378.150000 ;
        RECT 551.000000 385.850000 556.000000 386.150000 ;
        RECT 551.000000 381.850000 556.000000 382.150000 ;
        RECT 551.000000 397.850000 556.000000 398.150000 ;
        RECT 551.000000 393.850000 556.000000 394.150000 ;
        RECT 551.000000 389.850000 556.000000 390.150000 ;
        RECT 551.000000 413.850000 556.000000 414.150000 ;
        RECT 551.000000 409.850000 556.000000 410.150000 ;
        RECT 551.000000 405.850000 556.000000 406.150000 ;
        RECT 551.000000 401.850000 556.000000 402.150000 ;
        RECT 451.000000 425.850000 456.000000 426.150000 ;
        RECT 451.000000 421.850000 456.000000 422.150000 ;
        RECT 451.000000 429.850000 456.000000 430.150000 ;
        RECT 451.000000 433.850000 456.000000 434.150000 ;
        RECT 451.000000 441.850000 456.000000 442.150000 ;
        RECT 451.000000 437.850000 456.000000 438.150000 ;
        RECT 451.000000 453.850000 456.000000 454.150000 ;
        RECT 451.000000 449.850000 456.000000 450.150000 ;
        RECT 451.000000 445.850000 456.000000 446.150000 ;
        RECT 501.000000 417.850000 506.000000 418.150000 ;
        RECT 501.000000 421.850000 506.000000 422.150000 ;
        RECT 501.000000 425.850000 506.000000 426.150000 ;
        RECT 501.000000 429.850000 506.000000 430.150000 ;
        RECT 501.000000 433.850000 506.000000 434.150000 ;
        RECT 501.000000 437.850000 506.000000 438.150000 ;
        RECT 501.000000 441.850000 506.000000 442.150000 ;
        RECT 501.000000 445.850000 506.000000 446.150000 ;
        RECT 501.000000 449.850000 506.000000 450.150000 ;
        RECT 501.000000 453.850000 506.000000 454.150000 ;
        RECT 451.000000 461.850000 456.000000 462.150000 ;
        RECT 451.000000 457.850000 456.000000 458.150000 ;
        RECT 451.000000 465.850000 456.000000 466.150000 ;
        RECT 451.000000 469.850000 456.000000 470.150000 ;
        RECT 451.000000 481.850000 456.000000 482.150000 ;
        RECT 451.000000 477.850000 456.000000 478.150000 ;
        RECT 451.000000 473.850000 456.000000 474.150000 ;
        RECT 451.000000 489.850000 456.000000 490.150000 ;
        RECT 451.000000 485.850000 456.000000 486.150000 ;
        RECT 501.000000 457.850000 506.000000 458.150000 ;
        RECT 501.000000 461.850000 506.000000 462.150000 ;
        RECT 501.000000 465.850000 506.000000 466.150000 ;
        RECT 501.000000 469.850000 506.000000 470.150000 ;
        RECT 501.000000 481.850000 506.000000 482.150000 ;
        RECT 501.000000 473.850000 506.000000 474.150000 ;
        RECT 501.000000 477.850000 506.000000 478.150000 ;
        RECT 501.000000 485.850000 506.000000 486.150000 ;
        RECT 501.000000 489.850000 506.000000 490.150000 ;
        RECT 551.000000 429.850000 556.000000 430.150000 ;
        RECT 551.000000 425.850000 556.000000 426.150000 ;
        RECT 551.000000 417.850000 556.000000 418.150000 ;
        RECT 551.000000 421.850000 556.000000 422.150000 ;
        RECT 551.000000 433.850000 556.000000 434.150000 ;
        RECT 551.000000 437.850000 556.000000 438.150000 ;
        RECT 551.000000 441.850000 556.000000 442.150000 ;
        RECT 551.000000 445.850000 556.000000 446.150000 ;
        RECT 551.000000 449.850000 556.000000 450.150000 ;
        RECT 551.000000 453.850000 556.000000 454.150000 ;
        RECT 551.000000 457.850000 556.000000 458.150000 ;
        RECT 551.000000 461.850000 556.000000 462.150000 ;
        RECT 551.000000 465.850000 556.000000 466.150000 ;
        RECT 551.000000 469.850000 556.000000 470.150000 ;
        RECT 551.000000 481.850000 556.000000 482.150000 ;
        RECT 551.000000 473.850000 556.000000 474.150000 ;
        RECT 551.000000 477.850000 556.000000 478.150000 ;
        RECT 551.000000 485.850000 556.000000 486.150000 ;
        RECT 551.000000 489.850000 556.000000 490.150000 ;
        RECT 301.000000 497.850000 306.000000 498.150000 ;
        RECT 301.000000 493.850000 306.000000 494.150000 ;
        RECT 301.000000 501.850000 306.000000 502.150000 ;
        RECT 301.000000 505.850000 306.000000 506.150000 ;
        RECT 301.000000 517.850000 306.000000 518.150000 ;
        RECT 301.000000 513.850000 306.000000 514.150000 ;
        RECT 301.000000 509.850000 306.000000 510.150000 ;
        RECT 351.000000 493.850000 356.000000 494.150000 ;
        RECT 351.000000 497.850000 356.000000 498.150000 ;
        RECT 351.000000 505.850000 356.000000 506.150000 ;
        RECT 351.000000 501.850000 356.000000 502.150000 ;
        RECT 351.000000 509.850000 356.000000 510.150000 ;
        RECT 351.000000 513.850000 356.000000 514.150000 ;
        RECT 351.000000 517.850000 356.000000 518.150000 ;
        RECT 351.000000 521.850000 356.000000 522.150000 ;
        RECT 351.000000 525.850000 356.000000 526.150000 ;
        RECT 351.000000 537.850000 356.000000 538.150000 ;
        RECT 351.000000 533.850000 356.000000 534.150000 ;
        RECT 351.000000 529.850000 356.000000 530.150000 ;
        RECT 351.000000 541.850000 356.000000 542.150000 ;
        RECT 351.000000 545.850000 356.000000 546.150000 ;
        RECT 351.000000 561.850000 356.000000 562.150000 ;
        RECT 351.000000 557.850000 356.000000 558.150000 ;
        RECT 351.000000 553.850000 356.000000 554.150000 ;
        RECT 351.000000 549.850000 356.000000 550.150000 ;
        RECT 375.000000 493.850000 385.000000 494.150000 ;
        RECT 375.000000 497.850000 385.000000 498.150000 ;
        RECT 375.000000 501.850000 385.000000 502.150000 ;
        RECT 375.000000 505.850000 385.000000 506.150000 ;
        RECT 401.000000 493.850000 406.000000 494.150000 ;
        RECT 401.000000 497.850000 406.000000 498.150000 ;
        RECT 401.000000 501.850000 406.000000 502.150000 ;
        RECT 375.000000 509.850000 385.000000 510.150000 ;
        RECT 375.000000 513.850000 385.000000 514.150000 ;
        RECT 375.000000 517.850000 385.000000 518.150000 ;
        RECT 375.000000 521.850000 385.000000 522.150000 ;
        RECT 375.000000 525.850000 385.000000 526.150000 ;
        RECT 375.000000 545.850000 385.000000 546.150000 ;
        RECT 375.000000 541.850000 385.000000 542.150000 ;
        RECT 375.000000 537.850000 385.000000 538.150000 ;
        RECT 375.000000 533.850000 385.000000 534.150000 ;
        RECT 375.000000 529.850000 385.000000 530.150000 ;
        RECT 375.000000 561.850000 385.000000 562.150000 ;
        RECT 375.000000 557.850000 385.000000 558.150000 ;
        RECT 375.000000 553.850000 385.000000 554.150000 ;
        RECT 375.000000 549.850000 385.000000 550.150000 ;
        RECT 351.000000 565.850000 356.000000 566.150000 ;
        RECT 351.000000 569.850000 356.000000 570.150000 ;
        RECT 351.000000 573.850000 356.000000 574.150000 ;
        RECT 351.000000 577.850000 356.000000 578.150000 ;
        RECT 351.000000 581.850000 356.000000 582.150000 ;
        RECT 351.000000 601.850000 356.000000 602.150000 ;
        RECT 351.000000 597.850000 356.000000 598.150000 ;
        RECT 351.000000 593.850000 356.000000 594.150000 ;
        RECT 351.000000 589.850000 356.000000 590.150000 ;
        RECT 351.000000 585.850000 356.000000 586.150000 ;
        RECT 351.000000 609.850000 356.000000 610.150000 ;
        RECT 351.000000 605.850000 356.000000 606.150000 ;
        RECT 351.000000 613.850000 356.000000 614.150000 ;
        RECT 351.000000 617.850000 356.000000 618.150000 ;
        RECT 351.000000 621.850000 356.000000 622.150000 ;
        RECT 351.000000 625.850000 356.000000 626.150000 ;
        RECT 351.000000 629.850000 356.000000 630.150000 ;
        RECT 351.000000 633.850000 356.000000 634.150000 ;
        RECT 351.000000 637.850000 356.000000 638.150000 ;
        RECT 375.000000 565.850000 385.000000 566.150000 ;
        RECT 375.000000 569.850000 385.000000 570.150000 ;
        RECT 375.000000 573.850000 385.000000 574.150000 ;
        RECT 375.000000 577.850000 385.000000 578.150000 ;
        RECT 375.000000 581.850000 385.000000 582.150000 ;
        RECT 375.000000 585.850000 385.000000 586.150000 ;
        RECT 375.000000 589.850000 385.000000 590.150000 ;
        RECT 375.000000 593.850000 385.000000 594.150000 ;
        RECT 375.000000 597.850000 385.000000 598.150000 ;
        RECT 375.000000 601.850000 385.000000 602.150000 ;
        RECT 375.000000 617.850000 385.000000 618.150000 ;
        RECT 375.000000 613.850000 385.000000 614.150000 ;
        RECT 375.000000 609.850000 385.000000 610.150000 ;
        RECT 375.000000 605.850000 385.000000 606.150000 ;
        RECT 375.000000 621.850000 385.000000 622.150000 ;
        RECT 375.000000 625.850000 385.000000 626.150000 ;
        RECT 375.000000 629.850000 385.000000 630.150000 ;
        RECT 375.000000 633.850000 385.000000 634.150000 ;
        RECT 375.000000 637.850000 385.000000 638.150000 ;
        RECT 451.000000 493.850000 456.000000 494.150000 ;
        RECT 451.000000 497.850000 456.000000 498.150000 ;
        RECT 451.000000 501.850000 456.000000 502.150000 ;
        RECT 501.000000 493.850000 506.000000 494.150000 ;
        RECT 501.000000 497.850000 506.000000 498.150000 ;
        RECT 501.000000 501.850000 506.000000 502.150000 ;
        RECT 551.000000 493.850000 556.000000 494.150000 ;
        RECT 551.000000 497.850000 556.000000 498.150000 ;
        RECT 551.000000 501.850000 556.000000 502.150000 ;
        RECT 351.000000 657.850000 356.000000 658.150000 ;
        RECT 351.000000 641.850000 356.000000 642.150000 ;
        RECT 351.000000 645.850000 356.000000 646.150000 ;
        RECT 351.000000 649.850000 356.000000 650.150000 ;
        RECT 351.000000 653.850000 356.000000 654.150000 ;
        RECT 351.000000 673.850000 356.000000 674.150000 ;
        RECT 351.000000 669.850000 356.000000 670.150000 ;
        RECT 351.000000 665.850000 356.000000 666.150000 ;
        RECT 351.000000 661.850000 356.000000 662.150000 ;
        RECT 301.000000 681.850000 306.000000 682.150000 ;
        RECT 301.000000 677.850000 306.000000 678.150000 ;
        RECT 351.000000 677.850000 356.000000 678.150000 ;
        RECT 351.000000 681.850000 356.000000 682.150000 ;
        RECT 375.000000 657.850000 385.000000 658.150000 ;
        RECT 401.000000 657.850000 406.000000 658.150000 ;
        RECT 375.000000 641.850000 385.000000 642.150000 ;
        RECT 375.000000 645.850000 385.000000 646.150000 ;
        RECT 375.000000 649.850000 385.000000 650.150000 ;
        RECT 375.000000 653.850000 385.000000 654.150000 ;
        RECT 375.000000 665.850000 385.000000 666.150000 ;
        RECT 375.000000 661.850000 385.000000 662.150000 ;
        RECT 375.000000 669.850000 385.000000 670.150000 ;
        RECT 375.000000 673.850000 385.000000 674.150000 ;
        RECT 401.000000 665.850000 406.000000 666.150000 ;
        RECT 401.000000 661.850000 406.000000 662.150000 ;
        RECT 401.000000 669.850000 406.000000 670.150000 ;
        RECT 401.000000 673.850000 406.000000 674.150000 ;
        RECT 401.000000 677.850000 406.000000 678.150000 ;
        RECT 375.000000 677.850000 385.000000 678.150000 ;
        RECT 401.000000 681.850000 406.000000 682.150000 ;
        RECT 375.000000 681.850000 385.000000 682.150000 ;
        RECT 451.000000 657.850000 456.000000 658.150000 ;
        RECT 451.000000 673.850000 456.000000 674.150000 ;
        RECT 451.000000 669.850000 456.000000 670.150000 ;
        RECT 451.000000 665.850000 456.000000 666.150000 ;
        RECT 451.000000 661.850000 456.000000 662.150000 ;
        RECT 501.000000 657.850000 506.000000 658.150000 ;
        RECT 501.000000 661.850000 506.000000 662.150000 ;
        RECT 501.000000 665.850000 506.000000 666.150000 ;
        RECT 501.000000 673.850000 506.000000 674.150000 ;
        RECT 501.000000 669.850000 506.000000 670.150000 ;
        RECT 451.000000 677.850000 456.000000 678.150000 ;
        RECT 451.000000 681.850000 456.000000 682.150000 ;
        RECT 501.000000 677.850000 506.000000 678.150000 ;
        RECT 501.000000 681.850000 506.000000 682.150000 ;
        RECT 551.000000 657.850000 556.000000 658.150000 ;
        RECT 551.000000 661.850000 556.000000 662.150000 ;
        RECT 551.000000 665.850000 556.000000 666.150000 ;
        RECT 551.000000 669.850000 556.000000 670.150000 ;
        RECT 551.000000 673.850000 556.000000 674.150000 ;
        RECT 551.000000 681.850000 556.000000 682.150000 ;
        RECT 551.000000 677.850000 556.000000 678.150000 ;
        RECT 601.000000 357.850000 606.000000 358.150000 ;
        RECT 601.000000 353.850000 606.000000 354.150000 ;
        RECT 601.000000 349.850000 606.000000 350.150000 ;
        RECT 601.000000 345.850000 606.000000 346.150000 ;
        RECT 601.000000 361.850000 606.000000 362.150000 ;
        RECT 601.000000 365.850000 606.000000 366.150000 ;
        RECT 601.000000 369.850000 606.000000 370.150000 ;
        RECT 601.000000 373.850000 606.000000 374.150000 ;
        RECT 601.000000 377.850000 606.000000 378.150000 ;
        RECT 651.000000 349.850000 656.000000 350.150000 ;
        RECT 651.000000 345.850000 656.000000 346.150000 ;
        RECT 651.000000 353.850000 656.000000 354.150000 ;
        RECT 651.000000 357.850000 656.000000 358.150000 ;
        RECT 651.000000 361.850000 656.000000 362.150000 ;
        RECT 651.000000 365.850000 656.000000 366.150000 ;
        RECT 651.000000 369.850000 656.000000 370.150000 ;
        RECT 651.000000 377.850000 656.000000 378.150000 ;
        RECT 651.000000 373.850000 656.000000 374.150000 ;
        RECT 601.000000 385.850000 606.000000 386.150000 ;
        RECT 601.000000 381.850000 606.000000 382.150000 ;
        RECT 601.000000 389.850000 606.000000 390.150000 ;
        RECT 601.000000 393.850000 606.000000 394.150000 ;
        RECT 601.000000 397.850000 606.000000 398.150000 ;
        RECT 601.000000 405.850000 606.000000 406.150000 ;
        RECT 601.000000 401.850000 606.000000 402.150000 ;
        RECT 601.000000 413.850000 606.000000 414.150000 ;
        RECT 601.000000 409.850000 606.000000 410.150000 ;
        RECT 651.000000 385.850000 656.000000 386.150000 ;
        RECT 651.000000 381.850000 656.000000 382.150000 ;
        RECT 651.000000 393.850000 656.000000 394.150000 ;
        RECT 651.000000 389.850000 656.000000 390.150000 ;
        RECT 651.000000 397.850000 656.000000 398.150000 ;
        RECT 651.000000 405.850000 656.000000 406.150000 ;
        RECT 651.000000 401.850000 656.000000 402.150000 ;
        RECT 651.000000 409.850000 656.000000 410.150000 ;
        RECT 651.000000 413.850000 656.000000 414.150000 ;
        RECT 701.000000 357.850000 706.000000 358.150000 ;
        RECT 701.000000 353.850000 706.000000 354.150000 ;
        RECT 701.000000 349.850000 706.000000 350.150000 ;
        RECT 701.000000 345.850000 706.000000 346.150000 ;
        RECT 701.000000 361.850000 706.000000 362.150000 ;
        RECT 701.000000 365.850000 706.000000 366.150000 ;
        RECT 701.000000 369.850000 706.000000 370.150000 ;
        RECT 701.000000 373.850000 706.000000 374.150000 ;
        RECT 701.000000 377.850000 706.000000 378.150000 ;
        RECT 701.000000 385.850000 706.000000 386.150000 ;
        RECT 701.000000 381.850000 706.000000 382.150000 ;
        RECT 701.000000 397.850000 706.000000 398.150000 ;
        RECT 701.000000 393.850000 706.000000 394.150000 ;
        RECT 701.000000 389.850000 706.000000 390.150000 ;
        RECT 701.000000 413.850000 706.000000 414.150000 ;
        RECT 701.000000 409.850000 706.000000 410.150000 ;
        RECT 701.000000 405.850000 706.000000 406.150000 ;
        RECT 701.000000 401.850000 706.000000 402.150000 ;
        RECT 601.000000 417.850000 606.000000 418.150000 ;
        RECT 601.000000 421.850000 606.000000 422.150000 ;
        RECT 601.000000 425.850000 606.000000 426.150000 ;
        RECT 601.000000 429.850000 606.000000 430.150000 ;
        RECT 601.000000 433.850000 606.000000 434.150000 ;
        RECT 601.000000 441.850000 606.000000 442.150000 ;
        RECT 601.000000 437.850000 606.000000 438.150000 ;
        RECT 601.000000 453.850000 606.000000 454.150000 ;
        RECT 601.000000 449.850000 606.000000 450.150000 ;
        RECT 601.000000 445.850000 606.000000 446.150000 ;
        RECT 651.000000 417.850000 656.000000 418.150000 ;
        RECT 651.000000 425.850000 656.000000 426.150000 ;
        RECT 651.000000 421.850000 656.000000 422.150000 ;
        RECT 651.000000 429.850000 656.000000 430.150000 ;
        RECT 651.000000 433.850000 656.000000 434.150000 ;
        RECT 651.000000 437.850000 656.000000 438.150000 ;
        RECT 651.000000 441.850000 656.000000 442.150000 ;
        RECT 651.000000 445.850000 656.000000 446.150000 ;
        RECT 651.000000 449.850000 656.000000 450.150000 ;
        RECT 651.000000 453.850000 656.000000 454.150000 ;
        RECT 601.000000 469.850000 606.000000 470.150000 ;
        RECT 601.000000 465.850000 606.000000 466.150000 ;
        RECT 601.000000 457.850000 606.000000 458.150000 ;
        RECT 601.000000 461.850000 606.000000 462.150000 ;
        RECT 601.000000 481.850000 606.000000 482.150000 ;
        RECT 601.000000 477.850000 606.000000 478.150000 ;
        RECT 601.000000 473.850000 606.000000 474.150000 ;
        RECT 601.000000 489.850000 606.000000 490.150000 ;
        RECT 601.000000 485.850000 606.000000 486.150000 ;
        RECT 651.000000 461.850000 656.000000 462.150000 ;
        RECT 651.000000 457.850000 656.000000 458.150000 ;
        RECT 651.000000 469.850000 656.000000 470.150000 ;
        RECT 651.000000 465.850000 656.000000 466.150000 ;
        RECT 651.000000 481.850000 656.000000 482.150000 ;
        RECT 651.000000 477.850000 656.000000 478.150000 ;
        RECT 651.000000 473.850000 656.000000 474.150000 ;
        RECT 651.000000 489.850000 656.000000 490.150000 ;
        RECT 651.000000 485.850000 656.000000 486.150000 ;
        RECT 701.000000 425.850000 706.000000 426.150000 ;
        RECT 701.000000 421.850000 706.000000 422.150000 ;
        RECT 701.000000 417.850000 706.000000 418.150000 ;
        RECT 701.000000 429.850000 706.000000 430.150000 ;
        RECT 701.000000 433.850000 706.000000 434.150000 ;
        RECT 701.000000 437.850000 706.000000 438.150000 ;
        RECT 701.000000 441.850000 706.000000 442.150000 ;
        RECT 701.000000 445.850000 706.000000 446.150000 ;
        RECT 701.000000 449.850000 706.000000 450.150000 ;
        RECT 701.000000 453.850000 706.000000 454.150000 ;
        RECT 725.000000 433.850000 735.000000 434.150000 ;
        RECT 725.000000 437.850000 735.000000 438.150000 ;
        RECT 725.000000 441.850000 735.000000 442.150000 ;
        RECT 725.000000 453.850000 735.000000 454.150000 ;
        RECT 725.000000 449.850000 735.000000 450.150000 ;
        RECT 725.000000 445.850000 735.000000 446.150000 ;
        RECT 701.000000 457.850000 706.000000 458.150000 ;
        RECT 701.000000 461.850000 706.000000 462.150000 ;
        RECT 701.000000 465.850000 706.000000 466.150000 ;
        RECT 701.000000 469.850000 706.000000 470.150000 ;
        RECT 701.000000 481.850000 706.000000 482.150000 ;
        RECT 701.000000 473.850000 706.000000 474.150000 ;
        RECT 701.000000 477.850000 706.000000 478.150000 ;
        RECT 701.000000 485.850000 706.000000 486.150000 ;
        RECT 701.000000 489.850000 706.000000 490.150000 ;
        RECT 725.000000 469.850000 735.000000 470.150000 ;
        RECT 725.000000 457.850000 735.000000 458.150000 ;
        RECT 725.000000 461.850000 735.000000 462.150000 ;
        RECT 725.000000 465.850000 735.000000 466.150000 ;
        RECT 725.000000 481.850000 735.000000 482.150000 ;
        RECT 725.000000 477.850000 735.000000 478.150000 ;
        RECT 725.000000 473.850000 735.000000 474.150000 ;
        RECT 725.000000 489.850000 735.000000 490.150000 ;
        RECT 725.000000 485.850000 735.000000 486.150000 ;
        RECT 751.000000 357.850000 756.000000 358.150000 ;
        RECT 751.000000 353.850000 756.000000 354.150000 ;
        RECT 751.000000 349.850000 756.000000 350.150000 ;
        RECT 751.000000 345.850000 756.000000 346.150000 ;
        RECT 751.000000 361.850000 756.000000 362.150000 ;
        RECT 751.000000 365.850000 756.000000 366.150000 ;
        RECT 751.000000 369.850000 756.000000 370.150000 ;
        RECT 751.000000 373.850000 756.000000 374.150000 ;
        RECT 751.000000 377.850000 756.000000 378.150000 ;
        RECT 801.000000 349.850000 806.000000 350.150000 ;
        RECT 801.000000 345.850000 806.000000 346.150000 ;
        RECT 801.000000 353.850000 806.000000 354.150000 ;
        RECT 801.000000 357.850000 806.000000 358.150000 ;
        RECT 801.000000 361.850000 806.000000 362.150000 ;
        RECT 801.000000 365.850000 806.000000 366.150000 ;
        RECT 801.000000 369.850000 806.000000 370.150000 ;
        RECT 801.000000 377.850000 806.000000 378.150000 ;
        RECT 801.000000 373.850000 806.000000 374.150000 ;
        RECT 751.000000 385.850000 756.000000 386.150000 ;
        RECT 751.000000 381.850000 756.000000 382.150000 ;
        RECT 751.000000 397.850000 756.000000 398.150000 ;
        RECT 751.000000 393.850000 756.000000 394.150000 ;
        RECT 751.000000 389.850000 756.000000 390.150000 ;
        RECT 751.000000 401.850000 756.000000 402.150000 ;
        RECT 751.000000 405.850000 756.000000 406.150000 ;
        RECT 751.000000 409.850000 756.000000 410.150000 ;
        RECT 751.000000 413.850000 756.000000 414.150000 ;
        RECT 801.000000 385.850000 806.000000 386.150000 ;
        RECT 801.000000 381.850000 806.000000 382.150000 ;
        RECT 801.000000 393.850000 806.000000 394.150000 ;
        RECT 801.000000 389.850000 806.000000 390.150000 ;
        RECT 801.000000 397.850000 806.000000 398.150000 ;
        RECT 801.000000 405.850000 806.000000 406.150000 ;
        RECT 801.000000 401.850000 806.000000 402.150000 ;
        RECT 801.000000 409.850000 806.000000 410.150000 ;
        RECT 801.000000 413.850000 806.000000 414.150000 ;
        RECT 851.000000 357.850000 856.000000 358.150000 ;
        RECT 851.000000 353.850000 856.000000 354.150000 ;
        RECT 851.000000 349.850000 856.000000 350.150000 ;
        RECT 851.000000 345.850000 856.000000 346.150000 ;
        RECT 851.000000 361.850000 856.000000 362.150000 ;
        RECT 851.000000 365.850000 856.000000 366.150000 ;
        RECT 851.000000 369.850000 856.000000 370.150000 ;
        RECT 851.000000 373.850000 856.000000 374.150000 ;
        RECT 851.000000 377.850000 856.000000 378.150000 ;
        RECT 851.000000 385.850000 856.000000 386.150000 ;
        RECT 851.000000 381.850000 856.000000 382.150000 ;
        RECT 851.000000 397.850000 856.000000 398.150000 ;
        RECT 851.000000 393.850000 856.000000 394.150000 ;
        RECT 851.000000 389.850000 856.000000 390.150000 ;
        RECT 851.000000 413.850000 856.000000 414.150000 ;
        RECT 851.000000 409.850000 856.000000 410.150000 ;
        RECT 851.000000 405.850000 856.000000 406.150000 ;
        RECT 851.000000 401.850000 856.000000 402.150000 ;
        RECT 751.000000 417.850000 756.000000 418.150000 ;
        RECT 751.000000 421.850000 756.000000 422.150000 ;
        RECT 751.000000 425.850000 756.000000 426.150000 ;
        RECT 751.000000 429.850000 756.000000 430.150000 ;
        RECT 751.000000 433.850000 756.000000 434.150000 ;
        RECT 751.000000 437.850000 756.000000 438.150000 ;
        RECT 751.000000 441.850000 756.000000 442.150000 ;
        RECT 801.000000 417.850000 806.000000 418.150000 ;
        RECT 801.000000 421.850000 806.000000 422.150000 ;
        RECT 801.000000 425.850000 806.000000 426.150000 ;
        RECT 801.000000 429.850000 806.000000 430.150000 ;
        RECT 801.000000 433.850000 806.000000 434.150000 ;
        RECT 801.000000 437.850000 806.000000 438.150000 ;
        RECT 801.000000 441.850000 806.000000 442.150000 ;
        RECT 851.000000 417.850000 856.000000 418.150000 ;
        RECT 851.000000 421.850000 856.000000 422.150000 ;
        RECT 851.000000 425.850000 856.000000 426.150000 ;
        RECT 851.000000 429.850000 856.000000 430.150000 ;
        RECT 851.000000 433.850000 856.000000 434.150000 ;
        RECT 851.000000 441.850000 856.000000 442.150000 ;
        RECT 851.000000 437.850000 856.000000 438.150000 ;
        RECT 601.000000 501.850000 606.000000 502.150000 ;
        RECT 601.000000 497.850000 606.000000 498.150000 ;
        RECT 601.000000 493.850000 606.000000 494.150000 ;
        RECT 651.000000 493.850000 656.000000 494.150000 ;
        RECT 651.000000 497.850000 656.000000 498.150000 ;
        RECT 651.000000 501.850000 656.000000 502.150000 ;
        RECT 701.000000 501.850000 706.000000 502.150000 ;
        RECT 701.000000 493.850000 706.000000 494.150000 ;
        RECT 701.000000 497.850000 706.000000 498.150000 ;
        RECT 725.000000 501.850000 735.000000 502.150000 ;
        RECT 725.000000 497.850000 735.000000 498.150000 ;
        RECT 725.000000 493.850000 735.000000 494.150000 ;
        RECT 901.000000 357.850000 906.000000 358.150000 ;
        RECT 901.000000 353.850000 906.000000 354.150000 ;
        RECT 901.000000 349.850000 906.000000 350.150000 ;
        RECT 901.000000 345.850000 906.000000 346.150000 ;
        RECT 901.000000 361.850000 906.000000 362.150000 ;
        RECT 901.000000 365.850000 906.000000 366.150000 ;
        RECT 901.000000 369.850000 906.000000 370.150000 ;
        RECT 901.000000 373.850000 906.000000 374.150000 ;
        RECT 901.000000 377.850000 906.000000 378.150000 ;
        RECT 951.000000 345.850000 956.000000 346.150000 ;
        RECT 951.000000 349.850000 956.000000 350.150000 ;
        RECT 951.000000 353.850000 956.000000 354.150000 ;
        RECT 951.000000 357.850000 956.000000 358.150000 ;
        RECT 951.000000 361.850000 956.000000 362.150000 ;
        RECT 951.000000 365.850000 956.000000 366.150000 ;
        RECT 951.000000 369.850000 956.000000 370.150000 ;
        RECT 951.000000 373.850000 956.000000 374.150000 ;
        RECT 951.000000 377.850000 956.000000 378.150000 ;
        RECT 901.000000 385.850000 906.000000 386.150000 ;
        RECT 901.000000 381.850000 906.000000 382.150000 ;
        RECT 901.000000 393.850000 906.000000 394.150000 ;
        RECT 901.000000 389.850000 906.000000 390.150000 ;
        RECT 901.000000 397.850000 906.000000 398.150000 ;
        RECT 901.000000 405.850000 906.000000 406.150000 ;
        RECT 901.000000 401.850000 906.000000 402.150000 ;
        RECT 901.000000 409.850000 906.000000 410.150000 ;
        RECT 901.000000 413.850000 906.000000 414.150000 ;
        RECT 951.000000 385.850000 956.000000 386.150000 ;
        RECT 951.000000 381.850000 956.000000 382.150000 ;
        RECT 951.000000 389.850000 956.000000 390.150000 ;
        RECT 951.000000 393.850000 956.000000 394.150000 ;
        RECT 951.000000 397.850000 956.000000 398.150000 ;
        RECT 951.000000 405.850000 956.000000 406.150000 ;
        RECT 951.000000 401.850000 956.000000 402.150000 ;
        RECT 951.000000 413.850000 956.000000 414.150000 ;
        RECT 951.000000 409.850000 956.000000 410.150000 ;
        RECT 1001.000000 349.850000 1006.000000 350.150000 ;
        RECT 1001.000000 345.850000 1006.000000 346.150000 ;
        RECT 1001.000000 353.850000 1006.000000 354.150000 ;
        RECT 1001.000000 357.850000 1006.000000 358.150000 ;
        RECT 1001.000000 361.850000 1006.000000 362.150000 ;
        RECT 1001.000000 365.850000 1006.000000 366.150000 ;
        RECT 1001.000000 369.850000 1006.000000 370.150000 ;
        RECT 1001.000000 377.850000 1006.000000 378.150000 ;
        RECT 1001.000000 373.850000 1006.000000 374.150000 ;
        RECT 1001.000000 385.850000 1006.000000 386.150000 ;
        RECT 1001.000000 381.850000 1006.000000 382.150000 ;
        RECT 1001.000000 393.850000 1006.000000 394.150000 ;
        RECT 1001.000000 389.850000 1006.000000 390.150000 ;
        RECT 1001.000000 397.850000 1006.000000 398.150000 ;
        RECT 1001.000000 405.850000 1006.000000 406.150000 ;
        RECT 1001.000000 401.850000 1006.000000 402.150000 ;
        RECT 1001.000000 409.850000 1006.000000 410.150000 ;
        RECT 1001.000000 413.850000 1006.000000 414.150000 ;
        RECT 901.000000 417.850000 906.000000 418.150000 ;
        RECT 901.000000 425.850000 906.000000 426.150000 ;
        RECT 901.000000 421.850000 906.000000 422.150000 ;
        RECT 901.000000 429.850000 906.000000 430.150000 ;
        RECT 901.000000 433.850000 906.000000 434.150000 ;
        RECT 901.000000 437.850000 906.000000 438.150000 ;
        RECT 901.000000 441.850000 906.000000 442.150000 ;
        RECT 951.000000 417.850000 956.000000 418.150000 ;
        RECT 951.000000 421.850000 956.000000 422.150000 ;
        RECT 951.000000 425.850000 956.000000 426.150000 ;
        RECT 951.000000 429.850000 956.000000 430.150000 ;
        RECT 951.000000 433.850000 956.000000 434.150000 ;
        RECT 951.000000 441.850000 956.000000 442.150000 ;
        RECT 951.000000 437.850000 956.000000 438.150000 ;
        RECT 1001.000000 425.850000 1006.000000 426.150000 ;
        RECT 1001.000000 421.850000 1006.000000 422.150000 ;
        RECT 1001.000000 417.850000 1006.000000 418.150000 ;
        RECT 1001.000000 433.850000 1006.000000 434.150000 ;
        RECT 1001.000000 429.850000 1006.000000 430.150000 ;
        RECT 1001.000000 437.850000 1006.000000 438.150000 ;
        RECT 1001.000000 441.850000 1006.000000 442.150000 ;
        RECT 1051.000000 357.850000 1056.000000 358.150000 ;
        RECT 1051.000000 353.850000 1056.000000 354.150000 ;
        RECT 1051.000000 349.850000 1056.000000 350.150000 ;
        RECT 1051.000000 345.850000 1056.000000 346.150000 ;
        RECT 1051.000000 361.850000 1056.000000 362.150000 ;
        RECT 1051.000000 365.850000 1056.000000 366.150000 ;
        RECT 1051.000000 369.850000 1056.000000 370.150000 ;
        RECT 1051.000000 373.850000 1056.000000 374.150000 ;
        RECT 1051.000000 377.850000 1056.000000 378.150000 ;
        RECT 1101.000000 345.850000 1106.000000 346.150000 ;
        RECT 1101.000000 349.850000 1106.000000 350.150000 ;
        RECT 1101.000000 353.850000 1106.000000 354.150000 ;
        RECT 1101.000000 357.850000 1106.000000 358.150000 ;
        RECT 1101.000000 361.850000 1106.000000 362.150000 ;
        RECT 1101.000000 365.850000 1106.000000 366.150000 ;
        RECT 1101.000000 369.850000 1106.000000 370.150000 ;
        RECT 1101.000000 373.850000 1106.000000 374.150000 ;
        RECT 1101.000000 377.850000 1106.000000 378.150000 ;
        RECT 1051.000000 385.850000 1056.000000 386.150000 ;
        RECT 1051.000000 381.850000 1056.000000 382.150000 ;
        RECT 1051.000000 393.850000 1056.000000 394.150000 ;
        RECT 1051.000000 389.850000 1056.000000 390.150000 ;
        RECT 1051.000000 397.850000 1056.000000 398.150000 ;
        RECT 1051.000000 405.850000 1056.000000 406.150000 ;
        RECT 1051.000000 401.850000 1056.000000 402.150000 ;
        RECT 1051.000000 409.850000 1056.000000 410.150000 ;
        RECT 1051.000000 413.850000 1056.000000 414.150000 ;
        RECT 1101.000000 397.850000 1106.000000 398.150000 ;
        RECT 1101.000000 393.850000 1106.000000 394.150000 ;
        RECT 1101.000000 389.850000 1106.000000 390.150000 ;
        RECT 1101.000000 381.850000 1106.000000 382.150000 ;
        RECT 1101.000000 385.850000 1106.000000 386.150000 ;
        RECT 1101.000000 405.850000 1106.000000 406.150000 ;
        RECT 1101.000000 401.850000 1106.000000 402.150000 ;
        RECT 1101.000000 413.850000 1106.000000 414.150000 ;
        RECT 1101.000000 409.850000 1106.000000 410.150000 ;
        RECT 1151.000000 357.850000 1156.000000 358.150000 ;
        RECT 1151.000000 353.850000 1156.000000 354.150000 ;
        RECT 1151.000000 349.850000 1156.000000 350.150000 ;
        RECT 1151.000000 345.850000 1156.000000 346.150000 ;
        RECT 1172.000000 357.850000 1182.000000 358.150000 ;
        RECT 1172.000000 353.850000 1182.000000 354.150000 ;
        RECT 1172.000000 349.850000 1182.000000 350.150000 ;
        RECT 1172.000000 345.850000 1182.000000 346.150000 ;
        RECT 1151.000000 365.850000 1156.000000 366.150000 ;
        RECT 1151.000000 361.850000 1156.000000 362.150000 ;
        RECT 1151.000000 369.850000 1156.000000 370.150000 ;
        RECT 1151.000000 373.850000 1156.000000 374.150000 ;
        RECT 1151.000000 377.850000 1156.000000 378.150000 ;
        RECT 1172.000000 369.850000 1182.000000 370.150000 ;
        RECT 1172.000000 365.850000 1182.000000 366.150000 ;
        RECT 1172.000000 361.850000 1182.000000 362.150000 ;
        RECT 1172.000000 373.850000 1182.000000 374.150000 ;
        RECT 1172.000000 377.850000 1182.000000 378.150000 ;
        RECT 1151.000000 385.850000 1156.000000 386.150000 ;
        RECT 1151.000000 381.850000 1156.000000 382.150000 ;
        RECT 1151.000000 393.850000 1156.000000 394.150000 ;
        RECT 1151.000000 389.850000 1156.000000 390.150000 ;
        RECT 1151.000000 397.850000 1156.000000 398.150000 ;
        RECT 1172.000000 385.850000 1182.000000 386.150000 ;
        RECT 1172.000000 381.850000 1182.000000 382.150000 ;
        RECT 1172.000000 389.850000 1182.000000 390.150000 ;
        RECT 1172.000000 393.850000 1182.000000 394.150000 ;
        RECT 1172.000000 397.850000 1182.000000 398.150000 ;
        RECT 1151.000000 405.850000 1156.000000 406.150000 ;
        RECT 1151.000000 401.850000 1156.000000 402.150000 ;
        RECT 1151.000000 409.850000 1156.000000 410.150000 ;
        RECT 1151.000000 413.850000 1156.000000 414.150000 ;
        RECT 1172.000000 405.850000 1182.000000 406.150000 ;
        RECT 1172.000000 401.850000 1182.000000 402.150000 ;
        RECT 1172.000000 409.850000 1182.000000 410.150000 ;
        RECT 1172.000000 413.850000 1182.000000 414.150000 ;
        RECT 1051.000000 425.850000 1056.000000 426.150000 ;
        RECT 1051.000000 417.850000 1056.000000 418.150000 ;
        RECT 1051.000000 421.850000 1056.000000 422.150000 ;
        RECT 1051.000000 429.850000 1056.000000 430.150000 ;
        RECT 1051.000000 433.850000 1056.000000 434.150000 ;
        RECT 1051.000000 437.850000 1056.000000 438.150000 ;
        RECT 1051.000000 441.850000 1056.000000 442.150000 ;
        RECT 1101.000000 433.850000 1106.000000 434.150000 ;
        RECT 1101.000000 429.850000 1106.000000 430.150000 ;
        RECT 1101.000000 425.850000 1106.000000 426.150000 ;
        RECT 1101.000000 421.850000 1106.000000 422.150000 ;
        RECT 1101.000000 417.850000 1106.000000 418.150000 ;
        RECT 1101.000000 441.850000 1106.000000 442.150000 ;
        RECT 1101.000000 437.850000 1106.000000 438.150000 ;
        RECT 1151.000000 417.850000 1156.000000 418.150000 ;
        RECT 1151.000000 421.850000 1156.000000 422.150000 ;
        RECT 1151.000000 425.850000 1156.000000 426.150000 ;
        RECT 1151.000000 429.850000 1156.000000 430.150000 ;
        RECT 1151.000000 433.850000 1156.000000 434.150000 ;
        RECT 1172.000000 425.850000 1182.000000 426.150000 ;
        RECT 1172.000000 417.850000 1182.000000 418.150000 ;
        RECT 1172.000000 421.850000 1182.000000 422.150000 ;
        RECT 1172.000000 429.850000 1182.000000 430.150000 ;
        RECT 1172.000000 433.850000 1182.000000 434.150000 ;
        RECT 1151.000000 437.850000 1156.000000 438.150000 ;
        RECT 1151.000000 441.850000 1156.000000 442.150000 ;
        RECT 1151.000000 453.850000 1156.000000 454.150000 ;
        RECT 1151.000000 449.850000 1156.000000 450.150000 ;
        RECT 1151.000000 445.850000 1156.000000 446.150000 ;
        RECT 1172.000000 437.850000 1182.000000 438.150000 ;
        RECT 1172.000000 441.850000 1182.000000 442.150000 ;
        RECT 1151.000000 461.850000 1156.000000 462.150000 ;
        RECT 1151.000000 457.850000 1156.000000 458.150000 ;
        RECT 1151.000000 465.850000 1156.000000 466.150000 ;
        RECT 1151.000000 469.850000 1156.000000 470.150000 ;
        RECT 1151.000000 481.850000 1156.000000 482.150000 ;
        RECT 1151.000000 477.850000 1156.000000 478.150000 ;
        RECT 1151.000000 473.850000 1156.000000 474.150000 ;
        RECT 1151.000000 489.850000 1156.000000 490.150000 ;
        RECT 1151.000000 485.850000 1156.000000 486.150000 ;
        RECT 1151.000000 493.850000 1156.000000 494.150000 ;
        RECT 1151.000000 497.850000 1156.000000 498.150000 ;
        RECT 1151.000000 505.850000 1156.000000 506.150000 ;
        RECT 1151.000000 501.850000 1156.000000 502.150000 ;
        RECT 1151.000000 509.850000 1156.000000 510.150000 ;
        RECT 1151.000000 513.850000 1156.000000 514.150000 ;
        RECT 1151.000000 517.850000 1156.000000 518.150000 ;
        RECT 1151.000000 521.850000 1156.000000 522.150000 ;
        RECT 1151.000000 525.850000 1156.000000 526.150000 ;
        RECT 1151.000000 533.850000 1156.000000 534.150000 ;
        RECT 1151.000000 529.850000 1156.000000 530.150000 ;
        RECT 1151.000000 545.850000 1156.000000 546.150000 ;
        RECT 1151.000000 537.850000 1156.000000 538.150000 ;
        RECT 1151.000000 541.850000 1156.000000 542.150000 ;
        RECT 1151.000000 553.850000 1156.000000 554.150000 ;
        RECT 1151.000000 549.850000 1156.000000 550.150000 ;
        RECT 1151.000000 561.850000 1156.000000 562.150000 ;
        RECT 1151.000000 557.850000 1156.000000 558.150000 ;
        RECT 1151.000000 565.850000 1156.000000 566.150000 ;
        RECT 1151.000000 569.850000 1156.000000 570.150000 ;
        RECT 1151.000000 573.850000 1156.000000 574.150000 ;
        RECT 1151.000000 577.850000 1156.000000 578.150000 ;
        RECT 1151.000000 581.850000 1156.000000 582.150000 ;
        RECT 1151.000000 589.850000 1156.000000 590.150000 ;
        RECT 1151.000000 585.850000 1156.000000 586.150000 ;
        RECT 1151.000000 593.850000 1156.000000 594.150000 ;
        RECT 1151.000000 597.850000 1156.000000 598.150000 ;
        RECT 1151.000000 601.850000 1156.000000 602.150000 ;
        RECT 1151.000000 609.850000 1156.000000 610.150000 ;
        RECT 1151.000000 605.850000 1156.000000 606.150000 ;
        RECT 1151.000000 613.850000 1156.000000 614.150000 ;
        RECT 1151.000000 617.850000 1156.000000 618.150000 ;
        RECT 1151.000000 621.850000 1156.000000 622.150000 ;
        RECT 1151.000000 625.850000 1156.000000 626.150000 ;
        RECT 1151.000000 629.850000 1156.000000 630.150000 ;
        RECT 1151.000000 637.850000 1156.000000 638.150000 ;
        RECT 1151.000000 633.850000 1156.000000 634.150000 ;
        RECT 601.000000 657.850000 606.000000 658.150000 ;
        RECT 601.000000 673.850000 606.000000 674.150000 ;
        RECT 601.000000 669.850000 606.000000 670.150000 ;
        RECT 601.000000 665.850000 606.000000 666.150000 ;
        RECT 601.000000 661.850000 606.000000 662.150000 ;
        RECT 651.000000 657.850000 656.000000 658.150000 ;
        RECT 651.000000 661.850000 656.000000 662.150000 ;
        RECT 651.000000 665.850000 656.000000 666.150000 ;
        RECT 651.000000 673.850000 656.000000 674.150000 ;
        RECT 651.000000 669.850000 656.000000 670.150000 ;
        RECT 601.000000 677.850000 606.000000 678.150000 ;
        RECT 601.000000 681.850000 606.000000 682.150000 ;
        RECT 651.000000 677.850000 656.000000 678.150000 ;
        RECT 651.000000 681.850000 656.000000 682.150000 ;
        RECT 1151.000000 657.850000 1156.000000 658.150000 ;
        RECT 1151.000000 641.850000 1156.000000 642.150000 ;
        RECT 1151.000000 645.850000 1156.000000 646.150000 ;
        RECT 1151.000000 653.850000 1156.000000 654.150000 ;
        RECT 1151.000000 649.850000 1156.000000 650.150000 ;
        RECT 1151.000000 665.850000 1156.000000 666.150000 ;
        RECT 1151.000000 661.850000 1156.000000 662.150000 ;
        RECT 1151.000000 669.850000 1156.000000 670.150000 ;
        RECT 1151.000000 673.850000 1156.000000 674.150000 ;
        RECT 1151.000000 681.850000 1156.000000 682.150000 ;
        RECT 1151.000000 677.850000 1156.000000 678.150000 ;
    END
# end of P/G power stripe data as pin

  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M7 ;
        RECT 60.000000 0.000000 65.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 60.000000 681.000000 65.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 110.000000 0.000000 115.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 110.000000 681.000000 115.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 160.000000 0.000000 165.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 210.000000 0.000000 215.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 260.000000 0.000000 265.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 260.000000 681.000000 265.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 310.000000 0.000000 315.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 310.000000 681.000000 315.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 360.000000 0.000000 365.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 360.000000 681.000000 365.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 410.000000 0.000000 415.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 410.000000 501.000000 415.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 410.000000 656.000000 415.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 410.000000 681.000000 415.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 460.000000 0.000000 465.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 460.000000 501.000000 465.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 460.000000 656.000000 465.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 460.000000 681.000000 465.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 510.000000 0.000000 515.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 510.000000 501.000000 515.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 510.000000 656.000000 515.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 510.000000 681.000000 515.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 560.000000 0.000000 565.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 560.000000 501.000000 565.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 560.000000 656.000000 565.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 560.000000 681.000000 565.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 610.000000 0.000000 615.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 610.000000 501.000000 615.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 610.000000 656.000000 615.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 610.000000 681.000000 615.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 660.000000 0.000000 665.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 660.000000 501.000000 665.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 660.000000 656.000000 665.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 660.000000 681.000000 665.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 710.000000 0.000000 715.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 710.000000 501.000000 715.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 760.000000 0.000000 765.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 760.000000 441.000000 765.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 810.000000 0.000000 815.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 810.000000 441.000000 815.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 860.000000 0.000000 865.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 860.000000 441.000000 865.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 910.000000 0.000000 915.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 910.000000 441.000000 915.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 960.000000 0.000000 965.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 960.000000 441.000000 965.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1010.000000 0.000000 1015.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1010.000000 441.000000 1015.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1060.000000 0.000000 1065.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1060.000000 441.000000 1065.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1110.000000 0.000000 1115.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1110.000000 441.000000 1115.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1160.000000 0.000000 1165.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1160.000000 681.000000 1165.000000 686.000000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER M2 ;
        RECT 60.000000 3.850000 65.000000 4.150000 ;
        RECT 60.000000 7.850000 65.000000 8.150000 ;
        RECT 110.000000 7.850000 115.000000 8.150000 ;
        RECT 110.000000 3.850000 115.000000 4.150000 ;
        RECT 160.000000 7.850000 165.000000 8.150000 ;
        RECT 160.000000 3.850000 165.000000 4.150000 ;
        RECT 210.000000 7.850000 215.000000 8.150000 ;
        RECT 210.000000 3.850000 215.000000 4.150000 ;
        RECT 260.000000 7.850000 265.000000 8.150000 ;
        RECT 260.000000 3.850000 265.000000 4.150000 ;
        RECT 310.000000 7.850000 315.000000 8.150000 ;
        RECT 310.000000 3.850000 315.000000 4.150000 ;
        RECT 360.000000 7.850000 365.000000 8.150000 ;
        RECT 360.000000 3.850000 365.000000 4.150000 ;
        RECT 410.000000 7.850000 415.000000 8.150000 ;
        RECT 410.000000 3.850000 415.000000 4.150000 ;
        RECT 460.000000 7.850000 465.000000 8.150000 ;
        RECT 460.000000 3.850000 465.000000 4.150000 ;
        RECT 510.000000 7.850000 515.000000 8.150000 ;
        RECT 510.000000 3.850000 515.000000 4.150000 ;
        RECT 560.000000 3.850000 565.000000 4.150000 ;
        RECT 560.000000 7.850000 565.000000 8.150000 ;
        RECT 18.000000 267.850000 28.000000 268.150000 ;
        RECT 18.000000 259.850000 28.000000 260.150000 ;
        RECT 18.000000 263.850000 28.000000 264.150000 ;
        RECT 60.000000 267.850000 65.000000 268.150000 ;
        RECT 60.000000 263.850000 65.000000 264.150000 ;
        RECT 60.000000 259.850000 65.000000 260.150000 ;
        RECT 110.000000 267.850000 115.000000 268.150000 ;
        RECT 110.000000 259.850000 115.000000 260.150000 ;
        RECT 110.000000 263.850000 115.000000 264.150000 ;
        RECT 18.000000 283.850000 28.000000 284.150000 ;
        RECT 18.000000 279.850000 28.000000 280.150000 ;
        RECT 18.000000 275.850000 28.000000 276.150000 ;
        RECT 18.000000 271.850000 28.000000 272.150000 ;
        RECT 18.000000 287.850000 28.000000 288.150000 ;
        RECT 18.000000 291.850000 28.000000 292.150000 ;
        RECT 18.000000 295.850000 28.000000 296.150000 ;
        RECT 18.000000 299.850000 28.000000 300.150000 ;
        RECT 18.000000 303.850000 28.000000 304.150000 ;
        RECT 60.000000 283.850000 65.000000 284.150000 ;
        RECT 60.000000 279.850000 65.000000 280.150000 ;
        RECT 60.000000 275.850000 65.000000 276.150000 ;
        RECT 60.000000 271.850000 65.000000 272.150000 ;
        RECT 60.000000 287.850000 65.000000 288.150000 ;
        RECT 60.000000 291.850000 65.000000 292.150000 ;
        RECT 60.000000 295.850000 65.000000 296.150000 ;
        RECT 60.000000 299.850000 65.000000 300.150000 ;
        RECT 60.000000 303.850000 65.000000 304.150000 ;
        RECT 18.000000 307.850000 28.000000 308.150000 ;
        RECT 18.000000 311.850000 28.000000 312.150000 ;
        RECT 18.000000 315.850000 28.000000 316.150000 ;
        RECT 18.000000 319.850000 28.000000 320.150000 ;
        RECT 18.000000 323.850000 28.000000 324.150000 ;
        RECT 18.000000 339.850000 28.000000 340.150000 ;
        RECT 18.000000 335.850000 28.000000 336.150000 ;
        RECT 18.000000 331.850000 28.000000 332.150000 ;
        RECT 18.000000 327.850000 28.000000 328.150000 ;
        RECT 60.000000 307.850000 65.000000 308.150000 ;
        RECT 60.000000 311.850000 65.000000 312.150000 ;
        RECT 60.000000 315.850000 65.000000 316.150000 ;
        RECT 60.000000 319.850000 65.000000 320.150000 ;
        RECT 60.000000 323.850000 65.000000 324.150000 ;
        RECT 60.000000 339.850000 65.000000 340.150000 ;
        RECT 60.000000 335.850000 65.000000 336.150000 ;
        RECT 60.000000 331.850000 65.000000 332.150000 ;
        RECT 60.000000 327.850000 65.000000 328.150000 ;
        RECT 110.000000 271.850000 115.000000 272.150000 ;
        RECT 110.000000 275.850000 115.000000 276.150000 ;
        RECT 110.000000 279.850000 115.000000 280.150000 ;
        RECT 110.000000 283.850000 115.000000 284.150000 ;
        RECT 110.000000 287.850000 115.000000 288.150000 ;
        RECT 110.000000 291.850000 115.000000 292.150000 ;
        RECT 110.000000 295.850000 115.000000 296.150000 ;
        RECT 110.000000 299.850000 115.000000 300.150000 ;
        RECT 110.000000 303.850000 115.000000 304.150000 ;
        RECT 110.000000 311.850000 115.000000 312.150000 ;
        RECT 110.000000 307.850000 115.000000 308.150000 ;
        RECT 110.000000 323.850000 115.000000 324.150000 ;
        RECT 110.000000 319.850000 115.000000 320.150000 ;
        RECT 110.000000 315.850000 115.000000 316.150000 ;
        RECT 110.000000 339.850000 115.000000 340.150000 ;
        RECT 110.000000 335.850000 115.000000 336.150000 ;
        RECT 110.000000 331.850000 115.000000 332.150000 ;
        RECT 110.000000 327.850000 115.000000 328.150000 ;
        RECT 160.000000 259.850000 165.000000 260.150000 ;
        RECT 160.000000 263.850000 165.000000 264.150000 ;
        RECT 160.000000 267.850000 165.000000 268.150000 ;
        RECT 210.000000 267.850000 215.000000 268.150000 ;
        RECT 210.000000 263.850000 215.000000 264.150000 ;
        RECT 210.000000 259.850000 215.000000 260.150000 ;
        RECT 260.000000 267.850000 265.000000 268.150000 ;
        RECT 260.000000 259.850000 265.000000 260.150000 ;
        RECT 260.000000 263.850000 265.000000 264.150000 ;
        RECT 160.000000 275.850000 165.000000 276.150000 ;
        RECT 160.000000 271.850000 165.000000 272.150000 ;
        RECT 160.000000 283.850000 165.000000 284.150000 ;
        RECT 160.000000 279.850000 165.000000 280.150000 ;
        RECT 160.000000 287.850000 165.000000 288.150000 ;
        RECT 160.000000 291.850000 165.000000 292.150000 ;
        RECT 160.000000 295.850000 165.000000 296.150000 ;
        RECT 160.000000 303.850000 165.000000 304.150000 ;
        RECT 160.000000 299.850000 165.000000 300.150000 ;
        RECT 210.000000 271.850000 215.000000 272.150000 ;
        RECT 210.000000 275.850000 215.000000 276.150000 ;
        RECT 210.000000 279.850000 215.000000 280.150000 ;
        RECT 210.000000 283.850000 215.000000 284.150000 ;
        RECT 210.000000 287.850000 215.000000 288.150000 ;
        RECT 210.000000 291.850000 215.000000 292.150000 ;
        RECT 210.000000 295.850000 215.000000 296.150000 ;
        RECT 210.000000 299.850000 215.000000 300.150000 ;
        RECT 210.000000 303.850000 215.000000 304.150000 ;
        RECT 160.000000 311.850000 165.000000 312.150000 ;
        RECT 160.000000 307.850000 165.000000 308.150000 ;
        RECT 160.000000 315.850000 165.000000 316.150000 ;
        RECT 160.000000 319.850000 165.000000 320.150000 ;
        RECT 160.000000 323.850000 165.000000 324.150000 ;
        RECT 160.000000 331.850000 165.000000 332.150000 ;
        RECT 160.000000 327.850000 165.000000 328.150000 ;
        RECT 160.000000 335.850000 165.000000 336.150000 ;
        RECT 160.000000 339.850000 165.000000 340.150000 ;
        RECT 210.000000 307.850000 215.000000 308.150000 ;
        RECT 210.000000 311.850000 215.000000 312.150000 ;
        RECT 210.000000 315.850000 215.000000 316.150000 ;
        RECT 210.000000 319.850000 215.000000 320.150000 ;
        RECT 210.000000 323.850000 215.000000 324.150000 ;
        RECT 210.000000 327.850000 215.000000 328.150000 ;
        RECT 210.000000 331.850000 215.000000 332.150000 ;
        RECT 210.000000 335.850000 215.000000 336.150000 ;
        RECT 210.000000 339.850000 215.000000 340.150000 ;
        RECT 260.000000 271.850000 265.000000 272.150000 ;
        RECT 260.000000 275.850000 265.000000 276.150000 ;
        RECT 260.000000 279.850000 265.000000 280.150000 ;
        RECT 260.000000 283.850000 265.000000 284.150000 ;
        RECT 260.000000 295.850000 265.000000 296.150000 ;
        RECT 260.000000 291.850000 265.000000 292.150000 ;
        RECT 260.000000 287.850000 265.000000 288.150000 ;
        RECT 260.000000 303.850000 265.000000 304.150000 ;
        RECT 260.000000 299.850000 265.000000 300.150000 ;
        RECT 260.000000 323.850000 265.000000 324.150000 ;
        RECT 260.000000 319.850000 265.000000 320.150000 ;
        RECT 260.000000 315.850000 265.000000 316.150000 ;
        RECT 260.000000 311.850000 265.000000 312.150000 ;
        RECT 260.000000 307.850000 265.000000 308.150000 ;
        RECT 260.000000 327.850000 265.000000 328.150000 ;
        RECT 260.000000 331.850000 265.000000 332.150000 ;
        RECT 260.000000 335.850000 265.000000 336.150000 ;
        RECT 260.000000 339.850000 265.000000 340.150000 ;
        RECT 310.000000 263.850000 315.000000 264.150000 ;
        RECT 310.000000 259.850000 315.000000 260.150000 ;
        RECT 310.000000 267.850000 315.000000 268.150000 ;
        RECT 360.000000 259.850000 365.000000 260.150000 ;
        RECT 360.000000 263.850000 365.000000 264.150000 ;
        RECT 360.000000 267.850000 365.000000 268.150000 ;
        RECT 410.000000 259.850000 415.000000 260.150000 ;
        RECT 410.000000 263.850000 415.000000 264.150000 ;
        RECT 410.000000 267.850000 415.000000 268.150000 ;
        RECT 310.000000 275.850000 315.000000 276.150000 ;
        RECT 310.000000 271.850000 315.000000 272.150000 ;
        RECT 310.000000 279.850000 315.000000 280.150000 ;
        RECT 310.000000 283.850000 315.000000 284.150000 ;
        RECT 310.000000 287.850000 315.000000 288.150000 ;
        RECT 310.000000 291.850000 315.000000 292.150000 ;
        RECT 310.000000 295.850000 315.000000 296.150000 ;
        RECT 310.000000 303.850000 315.000000 304.150000 ;
        RECT 310.000000 299.850000 315.000000 300.150000 ;
        RECT 360.000000 283.850000 365.000000 284.150000 ;
        RECT 360.000000 279.850000 365.000000 280.150000 ;
        RECT 360.000000 275.850000 365.000000 276.150000 ;
        RECT 360.000000 271.850000 365.000000 272.150000 ;
        RECT 360.000000 287.850000 365.000000 288.150000 ;
        RECT 360.000000 291.850000 365.000000 292.150000 ;
        RECT 360.000000 295.850000 365.000000 296.150000 ;
        RECT 360.000000 299.850000 365.000000 300.150000 ;
        RECT 360.000000 303.850000 365.000000 304.150000 ;
        RECT 310.000000 311.850000 315.000000 312.150000 ;
        RECT 310.000000 307.850000 315.000000 308.150000 ;
        RECT 310.000000 315.850000 315.000000 316.150000 ;
        RECT 310.000000 319.850000 315.000000 320.150000 ;
        RECT 310.000000 323.850000 315.000000 324.150000 ;
        RECT 310.000000 327.850000 315.000000 328.150000 ;
        RECT 310.000000 331.850000 315.000000 332.150000 ;
        RECT 310.000000 335.850000 315.000000 336.150000 ;
        RECT 310.000000 339.850000 315.000000 340.150000 ;
        RECT 360.000000 307.850000 365.000000 308.150000 ;
        RECT 360.000000 311.850000 365.000000 312.150000 ;
        RECT 360.000000 315.850000 365.000000 316.150000 ;
        RECT 360.000000 319.850000 365.000000 320.150000 ;
        RECT 360.000000 323.850000 365.000000 324.150000 ;
        RECT 360.000000 327.850000 365.000000 328.150000 ;
        RECT 360.000000 331.850000 365.000000 332.150000 ;
        RECT 360.000000 335.850000 365.000000 336.150000 ;
        RECT 360.000000 339.850000 365.000000 340.150000 ;
        RECT 410.000000 271.850000 415.000000 272.150000 ;
        RECT 410.000000 275.850000 415.000000 276.150000 ;
        RECT 410.000000 283.850000 415.000000 284.150000 ;
        RECT 410.000000 279.850000 415.000000 280.150000 ;
        RECT 410.000000 295.850000 415.000000 296.150000 ;
        RECT 410.000000 291.850000 415.000000 292.150000 ;
        RECT 410.000000 287.850000 415.000000 288.150000 ;
        RECT 410.000000 299.850000 415.000000 300.150000 ;
        RECT 410.000000 303.850000 415.000000 304.150000 ;
        RECT 410.000000 323.850000 415.000000 324.150000 ;
        RECT 410.000000 319.850000 415.000000 320.150000 ;
        RECT 410.000000 315.850000 415.000000 316.150000 ;
        RECT 410.000000 311.850000 415.000000 312.150000 ;
        RECT 410.000000 307.850000 415.000000 308.150000 ;
        RECT 410.000000 327.850000 415.000000 328.150000 ;
        RECT 410.000000 331.850000 415.000000 332.150000 ;
        RECT 410.000000 335.850000 415.000000 336.150000 ;
        RECT 410.000000 339.850000 415.000000 340.150000 ;
        RECT 460.000000 259.850000 465.000000 260.150000 ;
        RECT 460.000000 263.850000 465.000000 264.150000 ;
        RECT 460.000000 267.850000 465.000000 268.150000 ;
        RECT 510.000000 259.850000 515.000000 260.150000 ;
        RECT 510.000000 263.850000 515.000000 264.150000 ;
        RECT 510.000000 267.850000 515.000000 268.150000 ;
        RECT 560.000000 263.850000 565.000000 264.150000 ;
        RECT 560.000000 259.850000 565.000000 260.150000 ;
        RECT 560.000000 267.850000 565.000000 268.150000 ;
        RECT 460.000000 283.850000 465.000000 284.150000 ;
        RECT 460.000000 279.850000 465.000000 280.150000 ;
        RECT 460.000000 275.850000 465.000000 276.150000 ;
        RECT 460.000000 271.850000 465.000000 272.150000 ;
        RECT 460.000000 287.850000 465.000000 288.150000 ;
        RECT 460.000000 291.850000 465.000000 292.150000 ;
        RECT 460.000000 295.850000 465.000000 296.150000 ;
        RECT 510.000000 275.850000 515.000000 276.150000 ;
        RECT 510.000000 271.850000 515.000000 272.150000 ;
        RECT 510.000000 283.850000 515.000000 284.150000 ;
        RECT 510.000000 279.850000 515.000000 280.150000 ;
        RECT 510.000000 291.850000 515.000000 292.150000 ;
        RECT 510.000000 287.850000 515.000000 288.150000 ;
        RECT 510.000000 295.850000 515.000000 296.150000 ;
        RECT 510.000000 303.850000 515.000000 304.150000 ;
        RECT 510.000000 299.850000 515.000000 300.150000 ;
        RECT 460.000000 319.850000 465.000000 320.150000 ;
        RECT 460.000000 323.850000 465.000000 324.150000 ;
        RECT 460.000000 339.850000 465.000000 340.150000 ;
        RECT 460.000000 335.850000 465.000000 336.150000 ;
        RECT 460.000000 331.850000 465.000000 332.150000 ;
        RECT 460.000000 327.850000 465.000000 328.150000 ;
        RECT 510.000000 311.850000 515.000000 312.150000 ;
        RECT 510.000000 307.850000 515.000000 308.150000 ;
        RECT 510.000000 315.850000 515.000000 316.150000 ;
        RECT 510.000000 319.850000 515.000000 320.150000 ;
        RECT 510.000000 323.850000 515.000000 324.150000 ;
        RECT 510.000000 331.850000 515.000000 332.150000 ;
        RECT 510.000000 327.850000 515.000000 328.150000 ;
        RECT 510.000000 335.850000 515.000000 336.150000 ;
        RECT 510.000000 339.850000 515.000000 340.150000 ;
        RECT 560.000000 271.850000 565.000000 272.150000 ;
        RECT 560.000000 275.850000 565.000000 276.150000 ;
        RECT 560.000000 279.850000 565.000000 280.150000 ;
        RECT 560.000000 283.850000 565.000000 284.150000 ;
        RECT 560.000000 291.850000 565.000000 292.150000 ;
        RECT 560.000000 287.850000 565.000000 288.150000 ;
        RECT 560.000000 295.850000 565.000000 296.150000 ;
        RECT 560.000000 303.850000 565.000000 304.150000 ;
        RECT 560.000000 299.850000 565.000000 300.150000 ;
        RECT 560.000000 323.850000 565.000000 324.150000 ;
        RECT 560.000000 319.850000 565.000000 320.150000 ;
        RECT 560.000000 315.850000 565.000000 316.150000 ;
        RECT 560.000000 311.850000 565.000000 312.150000 ;
        RECT 560.000000 307.850000 565.000000 308.150000 ;
        RECT 560.000000 339.850000 565.000000 340.150000 ;
        RECT 560.000000 335.850000 565.000000 336.150000 ;
        RECT 560.000000 331.850000 565.000000 332.150000 ;
        RECT 560.000000 327.850000 565.000000 328.150000 ;
        RECT 610.000000 3.850000 615.000000 4.150000 ;
        RECT 610.000000 7.850000 615.000000 8.150000 ;
        RECT 660.000000 7.850000 665.000000 8.150000 ;
        RECT 660.000000 3.850000 665.000000 4.150000 ;
        RECT 710.000000 7.850000 715.000000 8.150000 ;
        RECT 710.000000 3.850000 715.000000 4.150000 ;
        RECT 760.000000 7.850000 765.000000 8.150000 ;
        RECT 760.000000 3.850000 765.000000 4.150000 ;
        RECT 810.000000 7.850000 815.000000 8.150000 ;
        RECT 810.000000 3.850000 815.000000 4.150000 ;
        RECT 860.000000 7.850000 865.000000 8.150000 ;
        RECT 860.000000 3.850000 865.000000 4.150000 ;
        RECT 960.000000 7.850000 965.000000 8.150000 ;
        RECT 960.000000 3.850000 965.000000 4.150000 ;
        RECT 910.000000 7.850000 915.000000 8.150000 ;
        RECT 910.000000 3.850000 915.000000 4.150000 ;
        RECT 1010.000000 7.850000 1015.000000 8.150000 ;
        RECT 1010.000000 3.850000 1015.000000 4.150000 ;
        RECT 1110.000000 7.850000 1115.000000 8.150000 ;
        RECT 1110.000000 3.850000 1115.000000 4.150000 ;
        RECT 1060.000000 7.850000 1065.000000 8.150000 ;
        RECT 1060.000000 3.850000 1065.000000 4.150000 ;
        RECT 1160.000000 3.850000 1165.000000 4.150000 ;
        RECT 1160.000000 7.850000 1165.000000 8.150000 ;
        RECT 1158.000000 27.850000 1168.000000 28.150000 ;
        RECT 1158.000000 23.850000 1168.000000 24.150000 ;
        RECT 1158.000000 19.850000 1168.000000 20.150000 ;
        RECT 1160.000000 15.850000 1165.000000 16.150000 ;
        RECT 1160.000000 11.850000 1165.000000 12.150000 ;
        RECT 1158.000000 31.850000 1168.000000 32.150000 ;
        RECT 1158.000000 35.850000 1168.000000 36.150000 ;
        RECT 1158.000000 43.850000 1168.000000 44.150000 ;
        RECT 1158.000000 39.850000 1168.000000 40.150000 ;
        RECT 610.000000 263.850000 615.000000 264.150000 ;
        RECT 610.000000 259.850000 615.000000 260.150000 ;
        RECT 610.000000 267.850000 615.000000 268.150000 ;
        RECT 660.000000 259.850000 665.000000 260.150000 ;
        RECT 660.000000 263.850000 665.000000 264.150000 ;
        RECT 660.000000 267.850000 665.000000 268.150000 ;
        RECT 710.000000 267.850000 715.000000 268.150000 ;
        RECT 710.000000 259.850000 715.000000 260.150000 ;
        RECT 710.000000 263.850000 715.000000 264.150000 ;
        RECT 610.000000 283.850000 615.000000 284.150000 ;
        RECT 610.000000 279.850000 615.000000 280.150000 ;
        RECT 610.000000 275.850000 615.000000 276.150000 ;
        RECT 610.000000 271.850000 615.000000 272.150000 ;
        RECT 610.000000 287.850000 615.000000 288.150000 ;
        RECT 610.000000 291.850000 615.000000 292.150000 ;
        RECT 610.000000 295.850000 615.000000 296.150000 ;
        RECT 610.000000 299.850000 615.000000 300.150000 ;
        RECT 610.000000 303.850000 615.000000 304.150000 ;
        RECT 660.000000 275.850000 665.000000 276.150000 ;
        RECT 660.000000 271.850000 665.000000 272.150000 ;
        RECT 660.000000 283.850000 665.000000 284.150000 ;
        RECT 660.000000 279.850000 665.000000 280.150000 ;
        RECT 660.000000 287.850000 665.000000 288.150000 ;
        RECT 660.000000 291.850000 665.000000 292.150000 ;
        RECT 660.000000 295.850000 665.000000 296.150000 ;
        RECT 660.000000 303.850000 665.000000 304.150000 ;
        RECT 660.000000 299.850000 665.000000 300.150000 ;
        RECT 610.000000 307.850000 615.000000 308.150000 ;
        RECT 610.000000 311.850000 615.000000 312.150000 ;
        RECT 610.000000 315.850000 615.000000 316.150000 ;
        RECT 610.000000 319.850000 615.000000 320.150000 ;
        RECT 610.000000 323.850000 615.000000 324.150000 ;
        RECT 610.000000 339.850000 615.000000 340.150000 ;
        RECT 610.000000 335.850000 615.000000 336.150000 ;
        RECT 610.000000 331.850000 615.000000 332.150000 ;
        RECT 610.000000 327.850000 615.000000 328.150000 ;
        RECT 660.000000 311.850000 665.000000 312.150000 ;
        RECT 660.000000 307.850000 665.000000 308.150000 ;
        RECT 660.000000 315.850000 665.000000 316.150000 ;
        RECT 660.000000 319.850000 665.000000 320.150000 ;
        RECT 660.000000 323.850000 665.000000 324.150000 ;
        RECT 660.000000 331.850000 665.000000 332.150000 ;
        RECT 660.000000 327.850000 665.000000 328.150000 ;
        RECT 660.000000 335.850000 665.000000 336.150000 ;
        RECT 660.000000 339.850000 665.000000 340.150000 ;
        RECT 710.000000 271.850000 715.000000 272.150000 ;
        RECT 710.000000 275.850000 715.000000 276.150000 ;
        RECT 710.000000 279.850000 715.000000 280.150000 ;
        RECT 710.000000 283.850000 715.000000 284.150000 ;
        RECT 710.000000 287.850000 715.000000 288.150000 ;
        RECT 710.000000 291.850000 715.000000 292.150000 ;
        RECT 710.000000 295.850000 715.000000 296.150000 ;
        RECT 710.000000 299.850000 715.000000 300.150000 ;
        RECT 710.000000 303.850000 715.000000 304.150000 ;
        RECT 710.000000 323.850000 715.000000 324.150000 ;
        RECT 710.000000 319.850000 715.000000 320.150000 ;
        RECT 710.000000 315.850000 715.000000 316.150000 ;
        RECT 710.000000 311.850000 715.000000 312.150000 ;
        RECT 710.000000 307.850000 715.000000 308.150000 ;
        RECT 710.000000 339.850000 715.000000 340.150000 ;
        RECT 710.000000 335.850000 715.000000 336.150000 ;
        RECT 710.000000 331.850000 715.000000 332.150000 ;
        RECT 710.000000 327.850000 715.000000 328.150000 ;
        RECT 760.000000 267.850000 765.000000 268.150000 ;
        RECT 760.000000 263.850000 765.000000 264.150000 ;
        RECT 760.000000 259.850000 765.000000 260.150000 ;
        RECT 810.000000 259.850000 815.000000 260.150000 ;
        RECT 810.000000 263.850000 815.000000 264.150000 ;
        RECT 810.000000 267.850000 815.000000 268.150000 ;
        RECT 860.000000 267.850000 865.000000 268.150000 ;
        RECT 860.000000 259.850000 865.000000 260.150000 ;
        RECT 860.000000 263.850000 865.000000 264.150000 ;
        RECT 760.000000 283.850000 765.000000 284.150000 ;
        RECT 760.000000 279.850000 765.000000 280.150000 ;
        RECT 760.000000 275.850000 765.000000 276.150000 ;
        RECT 760.000000 271.850000 765.000000 272.150000 ;
        RECT 760.000000 287.850000 765.000000 288.150000 ;
        RECT 760.000000 291.850000 765.000000 292.150000 ;
        RECT 760.000000 295.850000 765.000000 296.150000 ;
        RECT 760.000000 299.850000 765.000000 300.150000 ;
        RECT 760.000000 303.850000 765.000000 304.150000 ;
        RECT 810.000000 275.850000 815.000000 276.150000 ;
        RECT 810.000000 271.850000 815.000000 272.150000 ;
        RECT 810.000000 283.850000 815.000000 284.150000 ;
        RECT 810.000000 279.850000 815.000000 280.150000 ;
        RECT 810.000000 287.850000 815.000000 288.150000 ;
        RECT 810.000000 291.850000 815.000000 292.150000 ;
        RECT 810.000000 295.850000 815.000000 296.150000 ;
        RECT 810.000000 303.850000 815.000000 304.150000 ;
        RECT 810.000000 299.850000 815.000000 300.150000 ;
        RECT 760.000000 307.850000 765.000000 308.150000 ;
        RECT 760.000000 311.850000 765.000000 312.150000 ;
        RECT 760.000000 315.850000 765.000000 316.150000 ;
        RECT 760.000000 319.850000 765.000000 320.150000 ;
        RECT 760.000000 323.850000 765.000000 324.150000 ;
        RECT 760.000000 339.850000 765.000000 340.150000 ;
        RECT 760.000000 335.850000 765.000000 336.150000 ;
        RECT 760.000000 331.850000 765.000000 332.150000 ;
        RECT 760.000000 327.850000 765.000000 328.150000 ;
        RECT 810.000000 311.850000 815.000000 312.150000 ;
        RECT 810.000000 307.850000 815.000000 308.150000 ;
        RECT 810.000000 315.850000 815.000000 316.150000 ;
        RECT 810.000000 319.850000 815.000000 320.150000 ;
        RECT 810.000000 323.850000 815.000000 324.150000 ;
        RECT 810.000000 331.850000 815.000000 332.150000 ;
        RECT 810.000000 327.850000 815.000000 328.150000 ;
        RECT 810.000000 335.850000 815.000000 336.150000 ;
        RECT 810.000000 339.850000 815.000000 340.150000 ;
        RECT 860.000000 271.850000 865.000000 272.150000 ;
        RECT 860.000000 275.850000 865.000000 276.150000 ;
        RECT 860.000000 279.850000 865.000000 280.150000 ;
        RECT 860.000000 283.850000 865.000000 284.150000 ;
        RECT 860.000000 287.850000 865.000000 288.150000 ;
        RECT 860.000000 291.850000 865.000000 292.150000 ;
        RECT 860.000000 295.850000 865.000000 296.150000 ;
        RECT 860.000000 299.850000 865.000000 300.150000 ;
        RECT 860.000000 303.850000 865.000000 304.150000 ;
        RECT 860.000000 323.850000 865.000000 324.150000 ;
        RECT 860.000000 319.850000 865.000000 320.150000 ;
        RECT 860.000000 315.850000 865.000000 316.150000 ;
        RECT 860.000000 311.850000 865.000000 312.150000 ;
        RECT 860.000000 307.850000 865.000000 308.150000 ;
        RECT 860.000000 339.850000 865.000000 340.150000 ;
        RECT 860.000000 335.850000 865.000000 336.150000 ;
        RECT 860.000000 331.850000 865.000000 332.150000 ;
        RECT 860.000000 327.850000 865.000000 328.150000 ;
        RECT 1158.000000 47.850000 1168.000000 48.150000 ;
        RECT 1158.000000 51.850000 1168.000000 52.150000 ;
        RECT 1158.000000 63.850000 1168.000000 64.150000 ;
        RECT 1158.000000 59.850000 1168.000000 60.150000 ;
        RECT 1158.000000 55.850000 1168.000000 56.150000 ;
        RECT 1158.000000 67.850000 1168.000000 68.150000 ;
        RECT 1158.000000 71.850000 1168.000000 72.150000 ;
        RECT 1158.000000 79.850000 1168.000000 80.150000 ;
        RECT 1158.000000 75.850000 1168.000000 76.150000 ;
        RECT 1158.000000 83.850000 1168.000000 84.150000 ;
        RECT 1158.000000 87.850000 1168.000000 88.150000 ;
        RECT 1158.000000 91.850000 1168.000000 92.150000 ;
        RECT 1158.000000 99.850000 1168.000000 100.150000 ;
        RECT 1158.000000 95.850000 1168.000000 96.150000 ;
        RECT 1158.000000 103.850000 1168.000000 104.150000 ;
        RECT 1158.000000 107.850000 1168.000000 108.150000 ;
        RECT 1158.000000 119.850000 1168.000000 120.150000 ;
        RECT 1158.000000 115.850000 1168.000000 116.150000 ;
        RECT 1158.000000 111.850000 1168.000000 112.150000 ;
        RECT 1158.000000 123.850000 1168.000000 124.150000 ;
        RECT 1158.000000 127.850000 1168.000000 128.150000 ;
        RECT 1158.000000 135.850000 1168.000000 136.150000 ;
        RECT 1158.000000 131.850000 1168.000000 132.150000 ;
        RECT 1158.000000 139.850000 1168.000000 140.150000 ;
        RECT 1158.000000 143.850000 1168.000000 144.150000 ;
        RECT 1158.000000 147.850000 1168.000000 148.150000 ;
        RECT 1158.000000 155.850000 1168.000000 156.150000 ;
        RECT 1158.000000 151.850000 1168.000000 152.150000 ;
        RECT 1158.000000 159.850000 1168.000000 160.150000 ;
        RECT 1158.000000 163.850000 1168.000000 164.150000 ;
        RECT 1158.000000 175.850000 1168.000000 176.150000 ;
        RECT 1158.000000 171.850000 1168.000000 172.150000 ;
        RECT 1158.000000 167.850000 1168.000000 168.150000 ;
        RECT 1158.000000 179.850000 1168.000000 180.150000 ;
        RECT 1158.000000 183.850000 1168.000000 184.150000 ;
        RECT 1158.000000 191.850000 1168.000000 192.150000 ;
        RECT 1158.000000 187.850000 1168.000000 188.150000 ;
        RECT 960.000000 267.850000 965.000000 268.150000 ;
        RECT 960.000000 263.850000 965.000000 264.150000 ;
        RECT 960.000000 259.850000 965.000000 260.150000 ;
        RECT 910.000000 267.850000 915.000000 268.150000 ;
        RECT 910.000000 263.850000 915.000000 264.150000 ;
        RECT 910.000000 259.850000 915.000000 260.150000 ;
        RECT 1010.000000 259.850000 1015.000000 260.150000 ;
        RECT 1010.000000 263.850000 1015.000000 264.150000 ;
        RECT 1010.000000 267.850000 1015.000000 268.150000 ;
        RECT 960.000000 283.850000 965.000000 284.150000 ;
        RECT 960.000000 279.850000 965.000000 280.150000 ;
        RECT 960.000000 275.850000 965.000000 276.150000 ;
        RECT 960.000000 271.850000 965.000000 272.150000 ;
        RECT 960.000000 287.850000 965.000000 288.150000 ;
        RECT 960.000000 291.850000 965.000000 292.150000 ;
        RECT 960.000000 295.850000 965.000000 296.150000 ;
        RECT 960.000000 299.850000 965.000000 300.150000 ;
        RECT 960.000000 303.850000 965.000000 304.150000 ;
        RECT 960.000000 311.850000 965.000000 312.150000 ;
        RECT 960.000000 307.850000 965.000000 308.150000 ;
        RECT 960.000000 323.850000 965.000000 324.150000 ;
        RECT 960.000000 319.850000 965.000000 320.150000 ;
        RECT 960.000000 315.850000 965.000000 316.150000 ;
        RECT 960.000000 339.850000 965.000000 340.150000 ;
        RECT 960.000000 335.850000 965.000000 336.150000 ;
        RECT 960.000000 331.850000 965.000000 332.150000 ;
        RECT 960.000000 327.850000 965.000000 328.150000 ;
        RECT 910.000000 283.850000 915.000000 284.150000 ;
        RECT 910.000000 279.850000 915.000000 280.150000 ;
        RECT 910.000000 275.850000 915.000000 276.150000 ;
        RECT 910.000000 271.850000 915.000000 272.150000 ;
        RECT 910.000000 287.850000 915.000000 288.150000 ;
        RECT 910.000000 291.850000 915.000000 292.150000 ;
        RECT 910.000000 295.850000 915.000000 296.150000 ;
        RECT 910.000000 299.850000 915.000000 300.150000 ;
        RECT 910.000000 303.850000 915.000000 304.150000 ;
        RECT 910.000000 307.850000 915.000000 308.150000 ;
        RECT 910.000000 311.850000 915.000000 312.150000 ;
        RECT 910.000000 315.850000 915.000000 316.150000 ;
        RECT 910.000000 319.850000 915.000000 320.150000 ;
        RECT 910.000000 323.850000 915.000000 324.150000 ;
        RECT 910.000000 339.850000 915.000000 340.150000 ;
        RECT 910.000000 335.850000 915.000000 336.150000 ;
        RECT 910.000000 331.850000 915.000000 332.150000 ;
        RECT 910.000000 327.850000 915.000000 328.150000 ;
        RECT 1010.000000 275.850000 1015.000000 276.150000 ;
        RECT 1010.000000 271.850000 1015.000000 272.150000 ;
        RECT 1010.000000 283.850000 1015.000000 284.150000 ;
        RECT 1010.000000 279.850000 1015.000000 280.150000 ;
        RECT 1010.000000 287.850000 1015.000000 288.150000 ;
        RECT 1010.000000 291.850000 1015.000000 292.150000 ;
        RECT 1010.000000 295.850000 1015.000000 296.150000 ;
        RECT 1010.000000 303.850000 1015.000000 304.150000 ;
        RECT 1010.000000 299.850000 1015.000000 300.150000 ;
        RECT 1010.000000 311.850000 1015.000000 312.150000 ;
        RECT 1010.000000 307.850000 1015.000000 308.150000 ;
        RECT 1010.000000 315.850000 1015.000000 316.150000 ;
        RECT 1010.000000 319.850000 1015.000000 320.150000 ;
        RECT 1010.000000 323.850000 1015.000000 324.150000 ;
        RECT 1010.000000 331.850000 1015.000000 332.150000 ;
        RECT 1010.000000 327.850000 1015.000000 328.150000 ;
        RECT 1010.000000 335.850000 1015.000000 336.150000 ;
        RECT 1010.000000 339.850000 1015.000000 340.150000 ;
        RECT 1110.000000 267.850000 1115.000000 268.150000 ;
        RECT 1110.000000 263.850000 1115.000000 264.150000 ;
        RECT 1110.000000 259.850000 1115.000000 260.150000 ;
        RECT 1060.000000 267.850000 1065.000000 268.150000 ;
        RECT 1060.000000 263.850000 1065.000000 264.150000 ;
        RECT 1060.000000 259.850000 1065.000000 260.150000 ;
        RECT 1158.000000 203.850000 1168.000000 204.150000 ;
        RECT 1158.000000 195.850000 1168.000000 196.150000 ;
        RECT 1158.000000 199.850000 1168.000000 200.150000 ;
        RECT 1158.000000 211.850000 1168.000000 212.150000 ;
        RECT 1158.000000 207.850000 1168.000000 208.150000 ;
        RECT 1158.000000 215.850000 1168.000000 216.150000 ;
        RECT 1158.000000 219.850000 1168.000000 220.150000 ;
        RECT 1158.000000 227.850000 1168.000000 228.150000 ;
        RECT 1158.000000 223.850000 1168.000000 224.150000 ;
        RECT 1158.000000 231.850000 1168.000000 232.150000 ;
        RECT 1158.000000 235.850000 1168.000000 236.150000 ;
        RECT 1158.000000 239.850000 1168.000000 240.150000 ;
        RECT 1158.000000 247.850000 1168.000000 248.150000 ;
        RECT 1158.000000 243.850000 1168.000000 244.150000 ;
        RECT 1158.000000 251.850000 1168.000000 252.150000 ;
        RECT 1158.000000 255.850000 1168.000000 256.150000 ;
        RECT 1158.000000 267.850000 1168.000000 268.150000 ;
        RECT 1158.000000 259.850000 1168.000000 260.150000 ;
        RECT 1158.000000 263.850000 1168.000000 264.150000 ;
        RECT 1110.000000 283.850000 1115.000000 284.150000 ;
        RECT 1110.000000 279.850000 1115.000000 280.150000 ;
        RECT 1110.000000 275.850000 1115.000000 276.150000 ;
        RECT 1110.000000 271.850000 1115.000000 272.150000 ;
        RECT 1110.000000 287.850000 1115.000000 288.150000 ;
        RECT 1110.000000 291.850000 1115.000000 292.150000 ;
        RECT 1110.000000 295.850000 1115.000000 296.150000 ;
        RECT 1110.000000 299.850000 1115.000000 300.150000 ;
        RECT 1110.000000 303.850000 1115.000000 304.150000 ;
        RECT 1110.000000 311.850000 1115.000000 312.150000 ;
        RECT 1110.000000 307.850000 1115.000000 308.150000 ;
        RECT 1110.000000 323.850000 1115.000000 324.150000 ;
        RECT 1110.000000 319.850000 1115.000000 320.150000 ;
        RECT 1110.000000 315.850000 1115.000000 316.150000 ;
        RECT 1110.000000 339.850000 1115.000000 340.150000 ;
        RECT 1110.000000 335.850000 1115.000000 336.150000 ;
        RECT 1110.000000 331.850000 1115.000000 332.150000 ;
        RECT 1110.000000 327.850000 1115.000000 328.150000 ;
        RECT 1060.000000 283.850000 1065.000000 284.150000 ;
        RECT 1060.000000 279.850000 1065.000000 280.150000 ;
        RECT 1060.000000 275.850000 1065.000000 276.150000 ;
        RECT 1060.000000 271.850000 1065.000000 272.150000 ;
        RECT 1060.000000 287.850000 1065.000000 288.150000 ;
        RECT 1060.000000 291.850000 1065.000000 292.150000 ;
        RECT 1060.000000 295.850000 1065.000000 296.150000 ;
        RECT 1060.000000 299.850000 1065.000000 300.150000 ;
        RECT 1060.000000 303.850000 1065.000000 304.150000 ;
        RECT 1060.000000 307.850000 1065.000000 308.150000 ;
        RECT 1060.000000 311.850000 1065.000000 312.150000 ;
        RECT 1060.000000 315.850000 1065.000000 316.150000 ;
        RECT 1060.000000 319.850000 1065.000000 320.150000 ;
        RECT 1060.000000 323.850000 1065.000000 324.150000 ;
        RECT 1060.000000 339.850000 1065.000000 340.150000 ;
        RECT 1060.000000 335.850000 1065.000000 336.150000 ;
        RECT 1060.000000 331.850000 1065.000000 332.150000 ;
        RECT 1060.000000 327.850000 1065.000000 328.150000 ;
        RECT 1158.000000 283.850000 1168.000000 284.150000 ;
        RECT 1158.000000 279.850000 1168.000000 280.150000 ;
        RECT 1158.000000 275.850000 1168.000000 276.150000 ;
        RECT 1158.000000 271.850000 1168.000000 272.150000 ;
        RECT 1158.000000 287.850000 1168.000000 288.150000 ;
        RECT 1158.000000 291.850000 1168.000000 292.150000 ;
        RECT 1158.000000 295.850000 1168.000000 296.150000 ;
        RECT 1158.000000 299.850000 1168.000000 300.150000 ;
        RECT 1158.000000 303.850000 1168.000000 304.150000 ;
        RECT 1158.000000 307.850000 1168.000000 308.150000 ;
        RECT 1158.000000 311.850000 1168.000000 312.150000 ;
        RECT 1158.000000 315.850000 1168.000000 316.150000 ;
        RECT 1158.000000 319.850000 1168.000000 320.150000 ;
        RECT 1158.000000 323.850000 1168.000000 324.150000 ;
        RECT 1158.000000 339.850000 1168.000000 340.150000 ;
        RECT 1158.000000 335.850000 1168.000000 336.150000 ;
        RECT 1158.000000 331.850000 1168.000000 332.150000 ;
        RECT 1158.000000 327.850000 1168.000000 328.150000 ;
        RECT 60.000000 379.850000 65.000000 380.150000 ;
        RECT 18.000000 379.850000 28.000000 380.150000 ;
        RECT 18.000000 343.850000 28.000000 344.150000 ;
        RECT 18.000000 347.850000 28.000000 348.150000 ;
        RECT 18.000000 351.850000 28.000000 352.150000 ;
        RECT 18.000000 359.850000 28.000000 360.150000 ;
        RECT 18.000000 355.850000 28.000000 356.150000 ;
        RECT 18.000000 375.850000 28.000000 376.150000 ;
        RECT 18.000000 371.850000 28.000000 372.150000 ;
        RECT 18.000000 367.850000 28.000000 368.150000 ;
        RECT 18.000000 363.850000 28.000000 364.150000 ;
        RECT 60.000000 347.850000 65.000000 348.150000 ;
        RECT 60.000000 343.850000 65.000000 344.150000 ;
        RECT 60.000000 375.850000 65.000000 376.150000 ;
        RECT 60.000000 371.850000 65.000000 372.150000 ;
        RECT 60.000000 367.850000 65.000000 368.150000 ;
        RECT 60.000000 363.850000 65.000000 364.150000 ;
        RECT 18.000000 395.850000 28.000000 396.150000 ;
        RECT 18.000000 391.850000 28.000000 392.150000 ;
        RECT 18.000000 387.850000 28.000000 388.150000 ;
        RECT 18.000000 383.850000 28.000000 384.150000 ;
        RECT 18.000000 407.850000 28.000000 408.150000 ;
        RECT 18.000000 399.850000 28.000000 400.150000 ;
        RECT 18.000000 403.850000 28.000000 404.150000 ;
        RECT 18.000000 411.850000 28.000000 412.150000 ;
        RECT 18.000000 415.850000 28.000000 416.150000 ;
        RECT 60.000000 395.850000 65.000000 396.150000 ;
        RECT 60.000000 391.850000 65.000000 392.150000 ;
        RECT 60.000000 387.850000 65.000000 388.150000 ;
        RECT 60.000000 383.850000 65.000000 384.150000 ;
        RECT 60.000000 407.850000 65.000000 408.150000 ;
        RECT 60.000000 399.850000 65.000000 400.150000 ;
        RECT 60.000000 403.850000 65.000000 404.150000 ;
        RECT 60.000000 411.850000 65.000000 412.150000 ;
        RECT 60.000000 415.850000 65.000000 416.150000 ;
        RECT 110.000000 379.850000 115.000000 380.150000 ;
        RECT 110.000000 351.850000 115.000000 352.150000 ;
        RECT 110.000000 347.850000 115.000000 348.150000 ;
        RECT 110.000000 343.850000 115.000000 344.150000 ;
        RECT 110.000000 359.850000 115.000000 360.150000 ;
        RECT 110.000000 355.850000 115.000000 356.150000 ;
        RECT 110.000000 375.850000 115.000000 376.150000 ;
        RECT 110.000000 371.850000 115.000000 372.150000 ;
        RECT 110.000000 367.850000 115.000000 368.150000 ;
        RECT 110.000000 363.850000 115.000000 364.150000 ;
        RECT 110.000000 383.850000 115.000000 384.150000 ;
        RECT 110.000000 387.850000 115.000000 388.150000 ;
        RECT 110.000000 391.850000 115.000000 392.150000 ;
        RECT 110.000000 395.850000 115.000000 396.150000 ;
        RECT 110.000000 407.850000 115.000000 408.150000 ;
        RECT 110.000000 399.850000 115.000000 400.150000 ;
        RECT 110.000000 403.850000 115.000000 404.150000 ;
        RECT 110.000000 411.850000 115.000000 412.150000 ;
        RECT 110.000000 415.850000 115.000000 416.150000 ;
        RECT 18.000000 431.850000 28.000000 432.150000 ;
        RECT 18.000000 427.850000 28.000000 428.150000 ;
        RECT 18.000000 423.850000 28.000000 424.150000 ;
        RECT 18.000000 419.850000 28.000000 420.150000 ;
        RECT 18.000000 435.850000 28.000000 436.150000 ;
        RECT 18.000000 439.850000 28.000000 440.150000 ;
        RECT 18.000000 443.850000 28.000000 444.150000 ;
        RECT 18.000000 447.850000 28.000000 448.150000 ;
        RECT 18.000000 451.850000 28.000000 452.150000 ;
        RECT 60.000000 431.850000 65.000000 432.150000 ;
        RECT 60.000000 427.850000 65.000000 428.150000 ;
        RECT 60.000000 423.850000 65.000000 424.150000 ;
        RECT 60.000000 419.850000 65.000000 420.150000 ;
        RECT 60.000000 435.850000 65.000000 436.150000 ;
        RECT 60.000000 439.850000 65.000000 440.150000 ;
        RECT 60.000000 443.850000 65.000000 444.150000 ;
        RECT 60.000000 447.850000 65.000000 448.150000 ;
        RECT 60.000000 451.850000 65.000000 452.150000 ;
        RECT 18.000000 455.850000 28.000000 456.150000 ;
        RECT 18.000000 459.850000 28.000000 460.150000 ;
        RECT 18.000000 463.850000 28.000000 464.150000 ;
        RECT 18.000000 467.850000 28.000000 468.150000 ;
        RECT 18.000000 471.850000 28.000000 472.150000 ;
        RECT 18.000000 487.850000 28.000000 488.150000 ;
        RECT 18.000000 483.850000 28.000000 484.150000 ;
        RECT 18.000000 479.850000 28.000000 480.150000 ;
        RECT 18.000000 475.850000 28.000000 476.150000 ;
        RECT 60.000000 455.850000 65.000000 456.150000 ;
        RECT 60.000000 459.850000 65.000000 460.150000 ;
        RECT 60.000000 463.850000 65.000000 464.150000 ;
        RECT 60.000000 467.850000 65.000000 468.150000 ;
        RECT 60.000000 471.850000 65.000000 472.150000 ;
        RECT 60.000000 487.850000 65.000000 488.150000 ;
        RECT 60.000000 483.850000 65.000000 484.150000 ;
        RECT 60.000000 479.850000 65.000000 480.150000 ;
        RECT 60.000000 475.850000 65.000000 476.150000 ;
        RECT 110.000000 419.850000 115.000000 420.150000 ;
        RECT 110.000000 423.850000 115.000000 424.150000 ;
        RECT 110.000000 427.850000 115.000000 428.150000 ;
        RECT 110.000000 431.850000 115.000000 432.150000 ;
        RECT 110.000000 435.850000 115.000000 436.150000 ;
        RECT 110.000000 439.850000 115.000000 440.150000 ;
        RECT 110.000000 443.850000 115.000000 444.150000 ;
        RECT 110.000000 447.850000 115.000000 448.150000 ;
        RECT 110.000000 451.850000 115.000000 452.150000 ;
        RECT 110.000000 459.850000 115.000000 460.150000 ;
        RECT 110.000000 455.850000 115.000000 456.150000 ;
        RECT 110.000000 471.850000 115.000000 472.150000 ;
        RECT 110.000000 467.850000 115.000000 468.150000 ;
        RECT 110.000000 463.850000 115.000000 464.150000 ;
        RECT 110.000000 487.850000 115.000000 488.150000 ;
        RECT 110.000000 483.850000 115.000000 484.150000 ;
        RECT 110.000000 479.850000 115.000000 480.150000 ;
        RECT 110.000000 475.850000 115.000000 476.150000 ;
        RECT 160.000000 379.850000 165.000000 380.150000 ;
        RECT 210.000000 379.850000 215.000000 380.150000 ;
        RECT 160.000000 343.850000 165.000000 344.150000 ;
        RECT 160.000000 347.850000 165.000000 348.150000 ;
        RECT 160.000000 351.850000 165.000000 352.150000 ;
        RECT 160.000000 355.850000 165.000000 356.150000 ;
        RECT 160.000000 359.850000 165.000000 360.150000 ;
        RECT 160.000000 363.850000 165.000000 364.150000 ;
        RECT 160.000000 367.850000 165.000000 368.150000 ;
        RECT 160.000000 375.850000 165.000000 376.150000 ;
        RECT 160.000000 371.850000 165.000000 372.150000 ;
        RECT 210.000000 343.850000 215.000000 344.150000 ;
        RECT 210.000000 347.850000 215.000000 348.150000 ;
        RECT 210.000000 351.850000 215.000000 352.150000 ;
        RECT 210.000000 355.850000 215.000000 356.150000 ;
        RECT 210.000000 359.850000 215.000000 360.150000 ;
        RECT 210.000000 363.850000 215.000000 364.150000 ;
        RECT 210.000000 367.850000 215.000000 368.150000 ;
        RECT 210.000000 371.850000 215.000000 372.150000 ;
        RECT 210.000000 375.850000 215.000000 376.150000 ;
        RECT 160.000000 387.850000 165.000000 388.150000 ;
        RECT 160.000000 383.850000 165.000000 384.150000 ;
        RECT 160.000000 391.850000 165.000000 392.150000 ;
        RECT 160.000000 395.850000 165.000000 396.150000 ;
        RECT 160.000000 399.850000 165.000000 400.150000 ;
        RECT 210.000000 383.850000 215.000000 384.150000 ;
        RECT 210.000000 387.850000 215.000000 388.150000 ;
        RECT 210.000000 391.850000 215.000000 392.150000 ;
        RECT 210.000000 395.850000 215.000000 396.150000 ;
        RECT 210.000000 407.850000 215.000000 408.150000 ;
        RECT 210.000000 399.850000 215.000000 400.150000 ;
        RECT 210.000000 403.850000 215.000000 404.150000 ;
        RECT 210.000000 411.850000 215.000000 412.150000 ;
        RECT 210.000000 415.850000 215.000000 416.150000 ;
        RECT 260.000000 379.850000 265.000000 380.150000 ;
        RECT 260.000000 343.850000 265.000000 344.150000 ;
        RECT 260.000000 347.850000 265.000000 348.150000 ;
        RECT 260.000000 351.850000 265.000000 352.150000 ;
        RECT 260.000000 355.850000 265.000000 356.150000 ;
        RECT 260.000000 359.850000 265.000000 360.150000 ;
        RECT 260.000000 367.850000 265.000000 368.150000 ;
        RECT 260.000000 363.850000 265.000000 364.150000 ;
        RECT 260.000000 375.850000 265.000000 376.150000 ;
        RECT 260.000000 371.850000 265.000000 372.150000 ;
        RECT 260.000000 383.850000 265.000000 384.150000 ;
        RECT 260.000000 387.850000 265.000000 388.150000 ;
        RECT 260.000000 391.850000 265.000000 392.150000 ;
        RECT 260.000000 395.850000 265.000000 396.150000 ;
        RECT 260.000000 399.850000 265.000000 400.150000 ;
        RECT 210.000000 431.850000 215.000000 432.150000 ;
        RECT 210.000000 427.850000 215.000000 428.150000 ;
        RECT 210.000000 423.850000 215.000000 424.150000 ;
        RECT 210.000000 419.850000 215.000000 420.150000 ;
        RECT 210.000000 435.850000 215.000000 436.150000 ;
        RECT 210.000000 439.850000 215.000000 440.150000 ;
        RECT 210.000000 443.850000 215.000000 444.150000 ;
        RECT 210.000000 447.850000 215.000000 448.150000 ;
        RECT 210.000000 451.850000 215.000000 452.150000 ;
        RECT 160.000000 463.850000 165.000000 464.150000 ;
        RECT 160.000000 467.850000 165.000000 468.150000 ;
        RECT 160.000000 471.850000 165.000000 472.150000 ;
        RECT 160.000000 479.850000 165.000000 480.150000 ;
        RECT 160.000000 475.850000 165.000000 476.150000 ;
        RECT 160.000000 487.850000 165.000000 488.150000 ;
        RECT 160.000000 483.850000 165.000000 484.150000 ;
        RECT 210.000000 455.850000 215.000000 456.150000 ;
        RECT 210.000000 459.850000 215.000000 460.150000 ;
        RECT 210.000000 463.850000 215.000000 464.150000 ;
        RECT 210.000000 467.850000 215.000000 468.150000 ;
        RECT 210.000000 471.850000 215.000000 472.150000 ;
        RECT 210.000000 475.850000 215.000000 476.150000 ;
        RECT 210.000000 479.850000 215.000000 480.150000 ;
        RECT 210.000000 483.850000 215.000000 484.150000 ;
        RECT 210.000000 487.850000 215.000000 488.150000 ;
        RECT 260.000000 467.850000 265.000000 468.150000 ;
        RECT 260.000000 463.850000 265.000000 464.150000 ;
        RECT 260.000000 471.850000 265.000000 472.150000 ;
        RECT 260.000000 475.850000 265.000000 476.150000 ;
        RECT 260.000000 479.850000 265.000000 480.150000 ;
        RECT 260.000000 483.850000 265.000000 484.150000 ;
        RECT 260.000000 487.850000 265.000000 488.150000 ;
        RECT 18.000000 491.850000 28.000000 492.150000 ;
        RECT 18.000000 495.850000 28.000000 496.150000 ;
        RECT 18.000000 499.850000 28.000000 500.150000 ;
        RECT 18.000000 503.850000 28.000000 504.150000 ;
        RECT 18.000000 507.850000 28.000000 508.150000 ;
        RECT 18.000000 515.850000 28.000000 516.150000 ;
        RECT 18.000000 511.850000 28.000000 512.150000 ;
        RECT 60.000000 491.850000 65.000000 492.150000 ;
        RECT 60.000000 495.850000 65.000000 496.150000 ;
        RECT 60.000000 499.850000 65.000000 500.150000 ;
        RECT 60.000000 503.850000 65.000000 504.150000 ;
        RECT 60.000000 507.850000 65.000000 508.150000 ;
        RECT 60.000000 515.850000 65.000000 516.150000 ;
        RECT 60.000000 511.850000 65.000000 512.150000 ;
        RECT 110.000000 499.850000 115.000000 500.150000 ;
        RECT 110.000000 495.850000 115.000000 496.150000 ;
        RECT 110.000000 491.850000 115.000000 492.150000 ;
        RECT 110.000000 507.850000 115.000000 508.150000 ;
        RECT 110.000000 503.850000 115.000000 504.150000 ;
        RECT 110.000000 515.850000 115.000000 516.150000 ;
        RECT 110.000000 511.850000 115.000000 512.150000 ;
        RECT 160.000000 491.850000 165.000000 492.150000 ;
        RECT 160.000000 495.850000 165.000000 496.150000 ;
        RECT 160.000000 499.850000 165.000000 500.150000 ;
        RECT 160.000000 507.850000 165.000000 508.150000 ;
        RECT 160.000000 503.850000 165.000000 504.150000 ;
        RECT 160.000000 515.850000 165.000000 516.150000 ;
        RECT 160.000000 511.850000 165.000000 512.150000 ;
        RECT 210.000000 491.850000 215.000000 492.150000 ;
        RECT 210.000000 495.850000 215.000000 496.150000 ;
        RECT 210.000000 499.850000 215.000000 500.150000 ;
        RECT 210.000000 503.850000 215.000000 504.150000 ;
        RECT 210.000000 507.850000 215.000000 508.150000 ;
        RECT 210.000000 515.850000 215.000000 516.150000 ;
        RECT 210.000000 511.850000 215.000000 512.150000 ;
        RECT 260.000000 495.850000 265.000000 496.150000 ;
        RECT 260.000000 491.850000 265.000000 492.150000 ;
        RECT 260.000000 499.850000 265.000000 500.150000 ;
        RECT 260.000000 503.850000 265.000000 504.150000 ;
        RECT 260.000000 507.850000 265.000000 508.150000 ;
        RECT 260.000000 515.850000 265.000000 516.150000 ;
        RECT 260.000000 511.850000 265.000000 512.150000 ;
        RECT 360.000000 379.850000 365.000000 380.150000 ;
        RECT 310.000000 379.850000 315.000000 380.150000 ;
        RECT 310.000000 343.850000 315.000000 344.150000 ;
        RECT 310.000000 351.850000 315.000000 352.150000 ;
        RECT 310.000000 347.850000 315.000000 348.150000 ;
        RECT 310.000000 355.850000 315.000000 356.150000 ;
        RECT 310.000000 359.850000 315.000000 360.150000 ;
        RECT 310.000000 363.850000 315.000000 364.150000 ;
        RECT 310.000000 367.850000 315.000000 368.150000 ;
        RECT 310.000000 371.850000 315.000000 372.150000 ;
        RECT 310.000000 375.850000 315.000000 376.150000 ;
        RECT 360.000000 343.850000 365.000000 344.150000 ;
        RECT 360.000000 347.850000 365.000000 348.150000 ;
        RECT 360.000000 351.850000 365.000000 352.150000 ;
        RECT 360.000000 355.850000 365.000000 356.150000 ;
        RECT 360.000000 359.850000 365.000000 360.150000 ;
        RECT 360.000000 363.850000 365.000000 364.150000 ;
        RECT 360.000000 367.850000 365.000000 368.150000 ;
        RECT 360.000000 371.850000 365.000000 372.150000 ;
        RECT 360.000000 375.850000 365.000000 376.150000 ;
        RECT 310.000000 383.850000 315.000000 384.150000 ;
        RECT 310.000000 387.850000 315.000000 388.150000 ;
        RECT 310.000000 391.850000 315.000000 392.150000 ;
        RECT 310.000000 395.850000 315.000000 396.150000 ;
        RECT 310.000000 407.850000 315.000000 408.150000 ;
        RECT 310.000000 399.850000 315.000000 400.150000 ;
        RECT 310.000000 403.850000 315.000000 404.150000 ;
        RECT 310.000000 411.850000 315.000000 412.150000 ;
        RECT 310.000000 415.850000 315.000000 416.150000 ;
        RECT 360.000000 383.850000 365.000000 384.150000 ;
        RECT 360.000000 387.850000 365.000000 388.150000 ;
        RECT 360.000000 391.850000 365.000000 392.150000 ;
        RECT 360.000000 395.850000 365.000000 396.150000 ;
        RECT 360.000000 407.850000 365.000000 408.150000 ;
        RECT 360.000000 399.850000 365.000000 400.150000 ;
        RECT 360.000000 403.850000 365.000000 404.150000 ;
        RECT 360.000000 411.850000 365.000000 412.150000 ;
        RECT 360.000000 415.850000 365.000000 416.150000 ;
        RECT 410.000000 379.850000 415.000000 380.150000 ;
        RECT 410.000000 359.850000 415.000000 360.150000 ;
        RECT 410.000000 355.850000 415.000000 356.150000 ;
        RECT 410.000000 351.850000 415.000000 352.150000 ;
        RECT 410.000000 347.850000 415.000000 348.150000 ;
        RECT 410.000000 343.850000 415.000000 344.150000 ;
        RECT 410.000000 367.850000 415.000000 368.150000 ;
        RECT 410.000000 363.850000 415.000000 364.150000 ;
        RECT 410.000000 371.850000 415.000000 372.150000 ;
        RECT 410.000000 375.850000 415.000000 376.150000 ;
        RECT 410.000000 383.850000 415.000000 384.150000 ;
        RECT 410.000000 387.850000 415.000000 388.150000 ;
        RECT 410.000000 391.850000 415.000000 392.150000 ;
        RECT 410.000000 395.850000 415.000000 396.150000 ;
        RECT 410.000000 407.850000 415.000000 408.150000 ;
        RECT 410.000000 399.850000 415.000000 400.150000 ;
        RECT 410.000000 403.850000 415.000000 404.150000 ;
        RECT 410.000000 411.850000 415.000000 412.150000 ;
        RECT 410.000000 415.850000 415.000000 416.150000 ;
        RECT 361.000000 479.850000 371.000000 480.150000 ;
        RECT 361.000000 483.850000 371.000000 484.150000 ;
        RECT 361.000000 487.850000 371.000000 488.150000 ;
        RECT 310.000000 419.850000 315.000000 420.150000 ;
        RECT 310.000000 423.850000 315.000000 424.150000 ;
        RECT 310.000000 427.850000 315.000000 428.150000 ;
        RECT 310.000000 431.850000 315.000000 432.150000 ;
        RECT 310.000000 439.850000 315.000000 440.150000 ;
        RECT 310.000000 435.850000 315.000000 436.150000 ;
        RECT 310.000000 443.850000 315.000000 444.150000 ;
        RECT 310.000000 447.850000 315.000000 448.150000 ;
        RECT 310.000000 451.850000 315.000000 452.150000 ;
        RECT 360.000000 419.850000 365.000000 420.150000 ;
        RECT 360.000000 423.850000 365.000000 424.150000 ;
        RECT 360.000000 427.850000 365.000000 428.150000 ;
        RECT 360.000000 431.850000 365.000000 432.150000 ;
        RECT 360.000000 435.850000 365.000000 436.150000 ;
        RECT 360.000000 439.850000 365.000000 440.150000 ;
        RECT 360.000000 443.850000 365.000000 444.150000 ;
        RECT 360.000000 447.850000 365.000000 448.150000 ;
        RECT 360.000000 451.850000 365.000000 452.150000 ;
        RECT 310.000000 455.850000 315.000000 456.150000 ;
        RECT 310.000000 459.850000 315.000000 460.150000 ;
        RECT 310.000000 467.850000 315.000000 468.150000 ;
        RECT 310.000000 463.850000 315.000000 464.150000 ;
        RECT 310.000000 471.850000 315.000000 472.150000 ;
        RECT 310.000000 475.850000 315.000000 476.150000 ;
        RECT 310.000000 479.850000 315.000000 480.150000 ;
        RECT 310.000000 483.850000 315.000000 484.150000 ;
        RECT 310.000000 487.850000 315.000000 488.150000 ;
        RECT 360.000000 455.850000 365.000000 456.150000 ;
        RECT 360.000000 459.850000 365.000000 460.150000 ;
        RECT 360.000000 471.850000 368.500000 472.150000 ;
        RECT 360.000000 463.850000 365.000000 464.150000 ;
        RECT 360.000000 467.850000 365.000000 468.150000 ;
        RECT 363.500000 475.850000 368.500000 476.150000 ;
        RECT 410.000000 419.850000 415.000000 420.150000 ;
        RECT 410.000000 423.850000 415.000000 424.150000 ;
        RECT 410.000000 431.850000 415.000000 432.150000 ;
        RECT 410.000000 427.850000 415.000000 428.150000 ;
        RECT 410.000000 435.850000 415.000000 436.150000 ;
        RECT 410.000000 439.850000 415.000000 440.150000 ;
        RECT 410.000000 443.850000 415.000000 444.150000 ;
        RECT 410.000000 447.850000 415.000000 448.150000 ;
        RECT 410.000000 451.850000 415.000000 452.150000 ;
        RECT 410.000000 459.850000 415.000000 460.150000 ;
        RECT 410.000000 455.850000 415.000000 456.150000 ;
        RECT 410.000000 467.850000 415.000000 468.150000 ;
        RECT 410.000000 463.850000 415.000000 464.150000 ;
        RECT 410.000000 471.850000 415.000000 472.150000 ;
        RECT 410.000000 479.850000 415.000000 480.150000 ;
        RECT 410.000000 475.850000 415.000000 476.150000 ;
        RECT 410.000000 487.850000 415.000000 488.150000 ;
        RECT 410.000000 483.850000 415.000000 484.150000 ;
        RECT 460.000000 379.850000 465.000000 380.150000 ;
        RECT 510.000000 379.850000 515.000000 380.150000 ;
        RECT 460.000000 347.850000 465.000000 348.150000 ;
        RECT 460.000000 343.850000 465.000000 344.150000 ;
        RECT 460.000000 375.850000 465.000000 376.150000 ;
        RECT 460.000000 371.850000 465.000000 372.150000 ;
        RECT 510.000000 343.850000 515.000000 344.150000 ;
        RECT 510.000000 347.850000 515.000000 348.150000 ;
        RECT 510.000000 351.850000 515.000000 352.150000 ;
        RECT 510.000000 359.850000 515.000000 360.150000 ;
        RECT 510.000000 355.850000 515.000000 356.150000 ;
        RECT 510.000000 363.850000 515.000000 364.150000 ;
        RECT 510.000000 367.850000 515.000000 368.150000 ;
        RECT 510.000000 375.850000 515.000000 376.150000 ;
        RECT 510.000000 371.850000 515.000000 372.150000 ;
        RECT 460.000000 383.850000 465.000000 384.150000 ;
        RECT 460.000000 387.850000 465.000000 388.150000 ;
        RECT 460.000000 391.850000 465.000000 392.150000 ;
        RECT 460.000000 395.850000 465.000000 396.150000 ;
        RECT 510.000000 387.850000 515.000000 388.150000 ;
        RECT 510.000000 383.850000 515.000000 384.150000 ;
        RECT 510.000000 391.850000 515.000000 392.150000 ;
        RECT 510.000000 395.850000 515.000000 396.150000 ;
        RECT 510.000000 407.850000 515.000000 408.150000 ;
        RECT 510.000000 399.850000 515.000000 400.150000 ;
        RECT 510.000000 403.850000 515.000000 404.150000 ;
        RECT 510.000000 411.850000 515.000000 412.150000 ;
        RECT 510.000000 415.850000 515.000000 416.150000 ;
        RECT 560.000000 379.850000 565.000000 380.150000 ;
        RECT 560.000000 359.850000 565.000000 360.150000 ;
        RECT 560.000000 355.850000 565.000000 356.150000 ;
        RECT 560.000000 351.850000 565.000000 352.150000 ;
        RECT 560.000000 347.850000 565.000000 348.150000 ;
        RECT 560.000000 343.850000 565.000000 344.150000 ;
        RECT 560.000000 375.850000 565.000000 376.150000 ;
        RECT 560.000000 371.850000 565.000000 372.150000 ;
        RECT 560.000000 367.850000 565.000000 368.150000 ;
        RECT 560.000000 363.850000 565.000000 364.150000 ;
        RECT 560.000000 383.850000 565.000000 384.150000 ;
        RECT 560.000000 387.850000 565.000000 388.150000 ;
        RECT 560.000000 395.850000 565.000000 396.150000 ;
        RECT 560.000000 391.850000 565.000000 392.150000 ;
        RECT 560.000000 407.850000 565.000000 408.150000 ;
        RECT 560.000000 403.850000 565.000000 404.150000 ;
        RECT 560.000000 399.850000 565.000000 400.150000 ;
        RECT 560.000000 415.850000 565.000000 416.150000 ;
        RECT 560.000000 411.850000 565.000000 412.150000 ;
        RECT 460.000000 419.850000 465.000000 420.150000 ;
        RECT 460.000000 431.850000 465.000000 432.150000 ;
        RECT 460.000000 427.850000 465.000000 428.150000 ;
        RECT 460.000000 423.850000 465.000000 424.150000 ;
        RECT 460.000000 435.850000 465.000000 436.150000 ;
        RECT 460.000000 439.850000 465.000000 440.150000 ;
        RECT 460.000000 443.850000 465.000000 444.150000 ;
        RECT 460.000000 447.850000 465.000000 448.150000 ;
        RECT 460.000000 451.850000 465.000000 452.150000 ;
        RECT 510.000000 419.850000 515.000000 420.150000 ;
        RECT 510.000000 423.850000 515.000000 424.150000 ;
        RECT 510.000000 431.850000 515.000000 432.150000 ;
        RECT 510.000000 427.850000 515.000000 428.150000 ;
        RECT 510.000000 439.850000 515.000000 440.150000 ;
        RECT 510.000000 435.850000 515.000000 436.150000 ;
        RECT 510.000000 443.850000 515.000000 444.150000 ;
        RECT 510.000000 447.850000 515.000000 448.150000 ;
        RECT 510.000000 451.850000 515.000000 452.150000 ;
        RECT 460.000000 455.850000 465.000000 456.150000 ;
        RECT 460.000000 459.850000 465.000000 460.150000 ;
        RECT 460.000000 463.850000 465.000000 464.150000 ;
        RECT 460.000000 467.850000 465.000000 468.150000 ;
        RECT 460.000000 471.850000 465.000000 472.150000 ;
        RECT 460.000000 487.850000 465.000000 488.150000 ;
        RECT 460.000000 483.850000 465.000000 484.150000 ;
        RECT 460.000000 479.850000 465.000000 480.150000 ;
        RECT 460.000000 475.850000 465.000000 476.150000 ;
        RECT 510.000000 455.850000 515.000000 456.150000 ;
        RECT 510.000000 459.850000 515.000000 460.150000 ;
        RECT 510.000000 467.850000 515.000000 468.150000 ;
        RECT 510.000000 463.850000 515.000000 464.150000 ;
        RECT 510.000000 471.850000 515.000000 472.150000 ;
        RECT 510.000000 475.850000 515.000000 476.150000 ;
        RECT 510.000000 479.850000 515.000000 480.150000 ;
        RECT 510.000000 483.850000 515.000000 484.150000 ;
        RECT 510.000000 487.850000 515.000000 488.150000 ;
        RECT 560.000000 419.850000 565.000000 420.150000 ;
        RECT 560.000000 423.850000 565.000000 424.150000 ;
        RECT 560.000000 427.850000 565.000000 428.150000 ;
        RECT 560.000000 431.850000 565.000000 432.150000 ;
        RECT 560.000000 435.850000 565.000000 436.150000 ;
        RECT 560.000000 439.850000 565.000000 440.150000 ;
        RECT 560.000000 443.850000 565.000000 444.150000 ;
        RECT 560.000000 451.850000 565.000000 452.150000 ;
        RECT 560.000000 447.850000 565.000000 448.150000 ;
        RECT 560.000000 455.850000 565.000000 456.150000 ;
        RECT 560.000000 459.850000 565.000000 460.150000 ;
        RECT 560.000000 471.850000 565.000000 472.150000 ;
        RECT 560.000000 463.850000 565.000000 464.150000 ;
        RECT 560.000000 467.850000 565.000000 468.150000 ;
        RECT 560.000000 487.850000 565.000000 488.150000 ;
        RECT 560.000000 483.850000 565.000000 484.150000 ;
        RECT 560.000000 479.850000 565.000000 480.150000 ;
        RECT 560.000000 475.850000 565.000000 476.150000 ;
        RECT 360.000000 499.850000 371.000000 500.150000 ;
        RECT 360.000000 491.850000 371.000000 492.150000 ;
        RECT 360.000000 495.850000 371.000000 496.150000 ;
        RECT 360.000000 507.850000 371.000000 508.150000 ;
        RECT 360.000000 503.850000 371.000000 504.150000 ;
        RECT 360.000000 511.850000 371.000000 512.150000 ;
        RECT 360.000000 515.850000 371.000000 516.150000 ;
        RECT 360.000000 527.850000 371.000000 528.150000 ;
        RECT 360.000000 523.850000 371.000000 524.150000 ;
        RECT 360.000000 519.850000 371.000000 520.150000 ;
        RECT 360.000000 535.850000 371.000000 536.150000 ;
        RECT 360.000000 531.850000 371.000000 532.150000 ;
        RECT 360.000000 543.850000 371.000000 544.150000 ;
        RECT 360.000000 539.850000 371.000000 540.150000 ;
        RECT 360.000000 555.850000 371.000000 556.150000 ;
        RECT 360.000000 547.850000 371.000000 548.150000 ;
        RECT 360.000000 551.850000 371.000000 552.150000 ;
        RECT 360.000000 563.850000 371.000000 564.150000 ;
        RECT 360.000000 559.850000 371.000000 560.150000 ;
        RECT 310.000000 495.850000 315.000000 496.150000 ;
        RECT 310.000000 491.850000 315.000000 492.150000 ;
        RECT 310.000000 499.850000 315.000000 500.150000 ;
        RECT 310.000000 507.850000 315.000000 508.150000 ;
        RECT 310.000000 503.850000 315.000000 504.150000 ;
        RECT 310.000000 515.850000 315.000000 516.150000 ;
        RECT 310.000000 511.850000 315.000000 512.150000 ;
        RECT 410.000000 491.850000 415.000000 492.150000 ;
        RECT 410.000000 495.850000 415.000000 496.150000 ;
        RECT 410.000000 499.850000 415.000000 500.150000 ;
        RECT 410.000000 503.850000 415.000000 504.150000 ;
        RECT 360.000000 583.850000 371.000000 584.150000 ;
        RECT 360.000000 571.850000 371.000000 572.150000 ;
        RECT 360.000000 567.850000 371.000000 568.150000 ;
        RECT 360.000000 579.850000 371.000000 580.150000 ;
        RECT 360.000000 575.850000 371.000000 576.150000 ;
        RECT 360.000000 587.850000 371.000000 588.150000 ;
        RECT 360.000000 591.850000 371.000000 592.150000 ;
        RECT 360.000000 599.850000 371.000000 600.150000 ;
        RECT 360.000000 595.850000 371.000000 596.150000 ;
        RECT 360.000000 607.850000 371.000000 608.150000 ;
        RECT 360.000000 603.850000 371.000000 604.150000 ;
        RECT 360.000000 619.850000 371.000000 620.150000 ;
        RECT 360.000000 615.850000 371.000000 616.150000 ;
        RECT 360.000000 611.850000 371.000000 612.150000 ;
        RECT 360.000000 623.850000 371.000000 624.150000 ;
        RECT 360.000000 627.850000 371.000000 628.150000 ;
        RECT 360.000000 635.850000 371.000000 636.150000 ;
        RECT 360.000000 631.850000 371.000000 632.150000 ;
        RECT 460.000000 503.850000 465.000000 504.150000 ;
        RECT 460.000000 499.850000 465.000000 500.150000 ;
        RECT 460.000000 491.850000 465.000000 492.150000 ;
        RECT 460.000000 495.850000 465.000000 496.150000 ;
        RECT 510.000000 495.850000 515.000000 496.150000 ;
        RECT 510.000000 491.850000 515.000000 492.150000 ;
        RECT 510.000000 499.850000 515.000000 500.150000 ;
        RECT 510.000000 503.850000 515.000000 504.150000 ;
        RECT 560.000000 503.850000 565.000000 504.150000 ;
        RECT 560.000000 499.850000 565.000000 500.150000 ;
        RECT 560.000000 495.850000 565.000000 496.150000 ;
        RECT 560.000000 491.850000 565.000000 492.150000 ;
        RECT 360.000000 647.850000 371.000000 648.150000 ;
        RECT 360.000000 639.850000 371.000000 640.150000 ;
        RECT 360.000000 643.850000 371.000000 644.150000 ;
        RECT 360.000000 655.850000 371.000000 656.150000 ;
        RECT 360.000000 651.850000 371.000000 652.150000 ;
        RECT 360.000000 667.850000 371.000000 668.150000 ;
        RECT 360.000000 663.850000 371.000000 664.150000 ;
        RECT 360.000000 659.850000 371.000000 660.150000 ;
        RECT 360.000000 675.850000 365.000000 676.150000 ;
        RECT 360.000000 671.850000 365.000000 672.150000 ;
        RECT 310.000000 679.850000 315.000000 680.150000 ;
        RECT 310.000000 683.850000 315.000000 684.150000 ;
        RECT 360.000000 679.850000 365.000000 680.150000 ;
        RECT 360.000000 683.850000 365.000000 684.150000 ;
        RECT 410.000000 659.850000 415.000000 660.150000 ;
        RECT 410.000000 663.850000 415.000000 664.150000 ;
        RECT 410.000000 667.850000 415.000000 668.150000 ;
        RECT 410.000000 671.850000 415.000000 672.150000 ;
        RECT 410.000000 675.850000 415.000000 676.150000 ;
        RECT 410.000000 683.850000 415.000000 684.150000 ;
        RECT 410.000000 679.850000 415.000000 680.150000 ;
        RECT 460.000000 659.850000 465.000000 660.150000 ;
        RECT 460.000000 663.850000 465.000000 664.150000 ;
        RECT 460.000000 667.850000 465.000000 668.150000 ;
        RECT 460.000000 671.850000 465.000000 672.150000 ;
        RECT 460.000000 675.850000 465.000000 676.150000 ;
        RECT 510.000000 659.850000 515.000000 660.150000 ;
        RECT 510.000000 663.850000 515.000000 664.150000 ;
        RECT 510.000000 667.850000 515.000000 668.150000 ;
        RECT 510.000000 671.850000 515.000000 672.150000 ;
        RECT 510.000000 675.850000 515.000000 676.150000 ;
        RECT 460.000000 683.850000 465.000000 684.150000 ;
        RECT 460.000000 679.850000 465.000000 680.150000 ;
        RECT 510.000000 683.850000 515.000000 684.150000 ;
        RECT 510.000000 679.850000 515.000000 680.150000 ;
        RECT 560.000000 659.850000 565.000000 660.150000 ;
        RECT 560.000000 663.850000 565.000000 664.150000 ;
        RECT 560.000000 667.850000 565.000000 668.150000 ;
        RECT 560.000000 671.850000 565.000000 672.150000 ;
        RECT 560.000000 675.850000 565.000000 676.150000 ;
        RECT 560.000000 683.850000 565.000000 684.150000 ;
        RECT 560.000000 679.850000 565.000000 680.150000 ;
        RECT 610.000000 379.850000 615.000000 380.150000 ;
        RECT 660.000000 379.850000 665.000000 380.150000 ;
        RECT 610.000000 343.850000 615.000000 344.150000 ;
        RECT 610.000000 347.850000 615.000000 348.150000 ;
        RECT 610.000000 351.850000 615.000000 352.150000 ;
        RECT 610.000000 355.850000 615.000000 356.150000 ;
        RECT 610.000000 359.850000 615.000000 360.150000 ;
        RECT 610.000000 375.850000 615.000000 376.150000 ;
        RECT 610.000000 371.850000 615.000000 372.150000 ;
        RECT 610.000000 367.850000 615.000000 368.150000 ;
        RECT 610.000000 363.850000 615.000000 364.150000 ;
        RECT 660.000000 343.850000 665.000000 344.150000 ;
        RECT 660.000000 347.850000 665.000000 348.150000 ;
        RECT 660.000000 351.850000 665.000000 352.150000 ;
        RECT 660.000000 359.850000 665.000000 360.150000 ;
        RECT 660.000000 355.850000 665.000000 356.150000 ;
        RECT 660.000000 363.850000 665.000000 364.150000 ;
        RECT 660.000000 367.850000 665.000000 368.150000 ;
        RECT 660.000000 375.850000 665.000000 376.150000 ;
        RECT 660.000000 371.850000 665.000000 372.150000 ;
        RECT 610.000000 395.850000 615.000000 396.150000 ;
        RECT 610.000000 391.850000 615.000000 392.150000 ;
        RECT 610.000000 387.850000 615.000000 388.150000 ;
        RECT 610.000000 383.850000 615.000000 384.150000 ;
        RECT 610.000000 407.850000 615.000000 408.150000 ;
        RECT 610.000000 399.850000 615.000000 400.150000 ;
        RECT 610.000000 403.850000 615.000000 404.150000 ;
        RECT 610.000000 411.850000 615.000000 412.150000 ;
        RECT 610.000000 415.850000 615.000000 416.150000 ;
        RECT 660.000000 387.850000 665.000000 388.150000 ;
        RECT 660.000000 383.850000 665.000000 384.150000 ;
        RECT 660.000000 391.850000 665.000000 392.150000 ;
        RECT 660.000000 395.850000 665.000000 396.150000 ;
        RECT 660.000000 407.850000 665.000000 408.150000 ;
        RECT 660.000000 403.850000 665.000000 404.150000 ;
        RECT 660.000000 399.850000 665.000000 400.150000 ;
        RECT 660.000000 411.850000 665.000000 412.150000 ;
        RECT 660.000000 415.850000 665.000000 416.150000 ;
        RECT 710.000000 379.850000 715.000000 380.150000 ;
        RECT 710.000000 359.850000 715.000000 360.150000 ;
        RECT 710.000000 355.850000 715.000000 356.150000 ;
        RECT 710.000000 351.850000 715.000000 352.150000 ;
        RECT 710.000000 347.850000 715.000000 348.150000 ;
        RECT 710.000000 343.850000 715.000000 344.150000 ;
        RECT 710.000000 375.850000 715.000000 376.150000 ;
        RECT 710.000000 371.850000 715.000000 372.150000 ;
        RECT 710.000000 367.850000 715.000000 368.150000 ;
        RECT 710.000000 363.850000 715.000000 364.150000 ;
        RECT 710.000000 395.850000 715.000000 396.150000 ;
        RECT 710.000000 391.850000 715.000000 392.150000 ;
        RECT 710.000000 387.850000 715.000000 388.150000 ;
        RECT 710.000000 383.850000 715.000000 384.150000 ;
        RECT 710.000000 407.850000 715.000000 408.150000 ;
        RECT 710.000000 403.850000 715.000000 404.150000 ;
        RECT 710.000000 399.850000 715.000000 400.150000 ;
        RECT 710.000000 411.850000 718.500000 412.150000 ;
        RECT 713.500000 415.850000 718.500000 416.150000 ;
        RECT 610.000000 431.850000 615.000000 432.150000 ;
        RECT 610.000000 427.850000 615.000000 428.150000 ;
        RECT 610.000000 423.850000 615.000000 424.150000 ;
        RECT 610.000000 419.850000 615.000000 420.150000 ;
        RECT 610.000000 435.850000 615.000000 436.150000 ;
        RECT 610.000000 439.850000 615.000000 440.150000 ;
        RECT 610.000000 443.850000 615.000000 444.150000 ;
        RECT 610.000000 447.850000 615.000000 448.150000 ;
        RECT 610.000000 451.850000 615.000000 452.150000 ;
        RECT 660.000000 419.850000 665.000000 420.150000 ;
        RECT 660.000000 423.850000 665.000000 424.150000 ;
        RECT 660.000000 431.850000 665.000000 432.150000 ;
        RECT 660.000000 427.850000 665.000000 428.150000 ;
        RECT 660.000000 439.850000 665.000000 440.150000 ;
        RECT 660.000000 435.850000 665.000000 436.150000 ;
        RECT 660.000000 443.850000 665.000000 444.150000 ;
        RECT 660.000000 447.850000 665.000000 448.150000 ;
        RECT 660.000000 451.850000 665.000000 452.150000 ;
        RECT 610.000000 455.850000 615.000000 456.150000 ;
        RECT 610.000000 459.850000 615.000000 460.150000 ;
        RECT 610.000000 463.850000 615.000000 464.150000 ;
        RECT 610.000000 467.850000 615.000000 468.150000 ;
        RECT 610.000000 471.850000 615.000000 472.150000 ;
        RECT 610.000000 487.850000 615.000000 488.150000 ;
        RECT 610.000000 483.850000 615.000000 484.150000 ;
        RECT 610.000000 479.850000 615.000000 480.150000 ;
        RECT 610.000000 475.850000 615.000000 476.150000 ;
        RECT 660.000000 459.850000 665.000000 460.150000 ;
        RECT 660.000000 455.850000 665.000000 456.150000 ;
        RECT 660.000000 463.850000 665.000000 464.150000 ;
        RECT 660.000000 467.850000 665.000000 468.150000 ;
        RECT 660.000000 471.850000 665.000000 472.150000 ;
        RECT 660.000000 479.850000 665.000000 480.150000 ;
        RECT 660.000000 475.850000 665.000000 476.150000 ;
        RECT 660.000000 487.850000 665.000000 488.150000 ;
        RECT 660.000000 483.850000 665.000000 484.150000 ;
        RECT 711.000000 423.850000 721.000000 424.150000 ;
        RECT 711.000000 419.850000 721.000000 420.150000 ;
        RECT 710.000000 431.850000 721.000000 432.150000 ;
        RECT 711.000000 427.850000 721.000000 428.150000 ;
        RECT 710.000000 435.850000 721.000000 436.150000 ;
        RECT 710.000000 439.850000 721.000000 440.150000 ;
        RECT 710.000000 443.850000 721.000000 444.150000 ;
        RECT 710.000000 451.850000 721.000000 452.150000 ;
        RECT 710.000000 447.850000 721.000000 448.150000 ;
        RECT 710.000000 455.850000 721.000000 456.150000 ;
        RECT 710.000000 459.850000 721.000000 460.150000 ;
        RECT 710.000000 471.850000 721.000000 472.150000 ;
        RECT 710.000000 463.850000 721.000000 464.150000 ;
        RECT 710.000000 467.850000 721.000000 468.150000 ;
        RECT 710.000000 475.850000 721.000000 476.150000 ;
        RECT 710.000000 479.850000 721.000000 480.150000 ;
        RECT 710.000000 483.850000 721.000000 484.150000 ;
        RECT 710.000000 487.850000 721.000000 488.150000 ;
        RECT 810.000000 379.850000 815.000000 380.150000 ;
        RECT 760.000000 379.850000 765.000000 380.150000 ;
        RECT 760.000000 343.850000 765.000000 344.150000 ;
        RECT 760.000000 347.850000 765.000000 348.150000 ;
        RECT 760.000000 351.850000 765.000000 352.150000 ;
        RECT 760.000000 355.850000 765.000000 356.150000 ;
        RECT 760.000000 359.850000 765.000000 360.150000 ;
        RECT 760.000000 375.850000 765.000000 376.150000 ;
        RECT 760.000000 371.850000 765.000000 372.150000 ;
        RECT 760.000000 367.850000 765.000000 368.150000 ;
        RECT 760.000000 363.850000 765.000000 364.150000 ;
        RECT 810.000000 343.850000 815.000000 344.150000 ;
        RECT 810.000000 347.850000 815.000000 348.150000 ;
        RECT 810.000000 351.850000 815.000000 352.150000 ;
        RECT 810.000000 359.850000 815.000000 360.150000 ;
        RECT 810.000000 355.850000 815.000000 356.150000 ;
        RECT 810.000000 363.850000 815.000000 364.150000 ;
        RECT 810.000000 367.850000 815.000000 368.150000 ;
        RECT 810.000000 375.850000 815.000000 376.150000 ;
        RECT 810.000000 371.850000 815.000000 372.150000 ;
        RECT 760.000000 395.850000 765.000000 396.150000 ;
        RECT 760.000000 391.850000 765.000000 392.150000 ;
        RECT 760.000000 387.850000 765.000000 388.150000 ;
        RECT 760.000000 383.850000 765.000000 384.150000 ;
        RECT 760.000000 407.850000 765.000000 408.150000 ;
        RECT 760.000000 399.850000 765.000000 400.150000 ;
        RECT 760.000000 403.850000 765.000000 404.150000 ;
        RECT 760.000000 411.850000 765.000000 412.150000 ;
        RECT 760.000000 415.850000 765.000000 416.150000 ;
        RECT 810.000000 387.850000 815.000000 388.150000 ;
        RECT 810.000000 383.850000 815.000000 384.150000 ;
        RECT 810.000000 391.850000 815.000000 392.150000 ;
        RECT 810.000000 395.850000 815.000000 396.150000 ;
        RECT 810.000000 407.850000 815.000000 408.150000 ;
        RECT 810.000000 403.850000 815.000000 404.150000 ;
        RECT 810.000000 399.850000 815.000000 400.150000 ;
        RECT 810.000000 411.850000 815.000000 412.150000 ;
        RECT 810.000000 415.850000 815.000000 416.150000 ;
        RECT 860.000000 379.850000 865.000000 380.150000 ;
        RECT 860.000000 359.850000 865.000000 360.150000 ;
        RECT 860.000000 355.850000 865.000000 356.150000 ;
        RECT 860.000000 351.850000 865.000000 352.150000 ;
        RECT 860.000000 347.850000 865.000000 348.150000 ;
        RECT 860.000000 343.850000 865.000000 344.150000 ;
        RECT 860.000000 375.850000 865.000000 376.150000 ;
        RECT 860.000000 371.850000 865.000000 372.150000 ;
        RECT 860.000000 367.850000 865.000000 368.150000 ;
        RECT 860.000000 363.850000 865.000000 364.150000 ;
        RECT 860.000000 395.850000 865.000000 396.150000 ;
        RECT 860.000000 391.850000 865.000000 392.150000 ;
        RECT 860.000000 387.850000 865.000000 388.150000 ;
        RECT 860.000000 383.850000 865.000000 384.150000 ;
        RECT 860.000000 407.850000 865.000000 408.150000 ;
        RECT 860.000000 403.850000 865.000000 404.150000 ;
        RECT 860.000000 399.850000 865.000000 400.150000 ;
        RECT 860.000000 415.850000 865.000000 416.150000 ;
        RECT 860.000000 411.850000 865.000000 412.150000 ;
        RECT 760.000000 419.850000 765.000000 420.150000 ;
        RECT 760.000000 423.850000 765.000000 424.150000 ;
        RECT 760.000000 427.850000 765.000000 428.150000 ;
        RECT 760.000000 431.850000 765.000000 432.150000 ;
        RECT 760.000000 443.850000 765.000000 444.150000 ;
        RECT 760.000000 439.850000 765.000000 440.150000 ;
        RECT 760.000000 435.850000 765.000000 436.150000 ;
        RECT 810.000000 419.850000 815.000000 420.150000 ;
        RECT 810.000000 423.850000 815.000000 424.150000 ;
        RECT 810.000000 427.850000 815.000000 428.150000 ;
        RECT 810.000000 431.850000 815.000000 432.150000 ;
        RECT 810.000000 439.850000 815.000000 440.150000 ;
        RECT 810.000000 435.850000 815.000000 436.150000 ;
        RECT 810.000000 443.850000 815.000000 444.150000 ;
        RECT 860.000000 419.850000 865.000000 420.150000 ;
        RECT 860.000000 423.850000 865.000000 424.150000 ;
        RECT 860.000000 427.850000 865.000000 428.150000 ;
        RECT 860.000000 431.850000 865.000000 432.150000 ;
        RECT 860.000000 443.850000 865.000000 444.150000 ;
        RECT 860.000000 439.850000 865.000000 440.150000 ;
        RECT 860.000000 435.850000 865.000000 436.150000 ;
        RECT 610.000000 503.850000 615.000000 504.150000 ;
        RECT 610.000000 499.850000 615.000000 500.150000 ;
        RECT 610.000000 491.850000 615.000000 492.150000 ;
        RECT 610.000000 495.850000 615.000000 496.150000 ;
        RECT 660.000000 495.850000 665.000000 496.150000 ;
        RECT 660.000000 491.850000 665.000000 492.150000 ;
        RECT 660.000000 499.850000 665.000000 500.150000 ;
        RECT 660.000000 503.850000 665.000000 504.150000 ;
        RECT 710.000000 503.850000 715.000000 504.150000 ;
        RECT 710.000000 499.850000 715.000000 500.150000 ;
        RECT 710.000000 495.850000 715.000000 496.150000 ;
        RECT 710.000000 491.850000 715.000000 492.150000 ;
        RECT 960.000000 379.850000 965.000000 380.150000 ;
        RECT 960.000000 343.850000 965.000000 344.150000 ;
        RECT 960.000000 347.850000 965.000000 348.150000 ;
        RECT 960.000000 351.850000 965.000000 352.150000 ;
        RECT 960.000000 359.850000 965.000000 360.150000 ;
        RECT 960.000000 355.850000 965.000000 356.150000 ;
        RECT 960.000000 375.850000 965.000000 376.150000 ;
        RECT 960.000000 371.850000 965.000000 372.150000 ;
        RECT 960.000000 367.850000 965.000000 368.150000 ;
        RECT 960.000000 363.850000 965.000000 364.150000 ;
        RECT 960.000000 383.850000 965.000000 384.150000 ;
        RECT 960.000000 387.850000 965.000000 388.150000 ;
        RECT 960.000000 391.850000 965.000000 392.150000 ;
        RECT 960.000000 395.850000 965.000000 396.150000 ;
        RECT 960.000000 407.850000 965.000000 408.150000 ;
        RECT 960.000000 399.850000 965.000000 400.150000 ;
        RECT 960.000000 403.850000 965.000000 404.150000 ;
        RECT 960.000000 411.850000 965.000000 412.150000 ;
        RECT 960.000000 415.850000 965.000000 416.150000 ;
        RECT 910.000000 379.850000 915.000000 380.150000 ;
        RECT 910.000000 343.850000 915.000000 344.150000 ;
        RECT 910.000000 347.850000 915.000000 348.150000 ;
        RECT 910.000000 351.850000 915.000000 352.150000 ;
        RECT 910.000000 355.850000 915.000000 356.150000 ;
        RECT 910.000000 359.850000 915.000000 360.150000 ;
        RECT 910.000000 375.850000 915.000000 376.150000 ;
        RECT 910.000000 371.850000 915.000000 372.150000 ;
        RECT 910.000000 367.850000 915.000000 368.150000 ;
        RECT 910.000000 363.850000 915.000000 364.150000 ;
        RECT 910.000000 383.850000 915.000000 384.150000 ;
        RECT 910.000000 387.850000 915.000000 388.150000 ;
        RECT 910.000000 391.850000 915.000000 392.150000 ;
        RECT 910.000000 395.850000 915.000000 396.150000 ;
        RECT 910.000000 407.850000 915.000000 408.150000 ;
        RECT 910.000000 399.850000 915.000000 400.150000 ;
        RECT 910.000000 403.850000 915.000000 404.150000 ;
        RECT 910.000000 411.850000 915.000000 412.150000 ;
        RECT 910.000000 415.850000 915.000000 416.150000 ;
        RECT 1010.000000 379.850000 1015.000000 380.150000 ;
        RECT 1010.000000 343.850000 1015.000000 344.150000 ;
        RECT 1010.000000 347.850000 1015.000000 348.150000 ;
        RECT 1010.000000 351.850000 1015.000000 352.150000 ;
        RECT 1010.000000 359.850000 1015.000000 360.150000 ;
        RECT 1010.000000 355.850000 1015.000000 356.150000 ;
        RECT 1010.000000 363.850000 1015.000000 364.150000 ;
        RECT 1010.000000 367.850000 1015.000000 368.150000 ;
        RECT 1010.000000 375.850000 1015.000000 376.150000 ;
        RECT 1010.000000 371.850000 1015.000000 372.150000 ;
        RECT 1010.000000 387.850000 1015.000000 388.150000 ;
        RECT 1010.000000 383.850000 1015.000000 384.150000 ;
        RECT 1010.000000 391.850000 1015.000000 392.150000 ;
        RECT 1010.000000 395.850000 1015.000000 396.150000 ;
        RECT 1010.000000 407.850000 1015.000000 408.150000 ;
        RECT 1010.000000 403.850000 1015.000000 404.150000 ;
        RECT 1010.000000 399.850000 1015.000000 400.150000 ;
        RECT 1010.000000 411.850000 1015.000000 412.150000 ;
        RECT 1010.000000 415.850000 1015.000000 416.150000 ;
        RECT 960.000000 431.850000 965.000000 432.150000 ;
        RECT 960.000000 427.850000 965.000000 428.150000 ;
        RECT 960.000000 423.850000 965.000000 424.150000 ;
        RECT 960.000000 419.850000 965.000000 420.150000 ;
        RECT 960.000000 443.850000 965.000000 444.150000 ;
        RECT 960.000000 439.850000 965.000000 440.150000 ;
        RECT 960.000000 435.850000 965.000000 436.150000 ;
        RECT 910.000000 431.850000 915.000000 432.150000 ;
        RECT 910.000000 427.850000 915.000000 428.150000 ;
        RECT 910.000000 423.850000 915.000000 424.150000 ;
        RECT 910.000000 419.850000 915.000000 420.150000 ;
        RECT 910.000000 435.850000 915.000000 436.150000 ;
        RECT 910.000000 439.850000 915.000000 440.150000 ;
        RECT 910.000000 443.850000 915.000000 444.150000 ;
        RECT 1010.000000 419.850000 1015.000000 420.150000 ;
        RECT 1010.000000 423.850000 1015.000000 424.150000 ;
        RECT 1010.000000 427.850000 1015.000000 428.150000 ;
        RECT 1010.000000 431.850000 1015.000000 432.150000 ;
        RECT 1010.000000 435.850000 1015.000000 436.150000 ;
        RECT 1010.000000 439.850000 1015.000000 440.150000 ;
        RECT 1010.000000 443.850000 1015.000000 444.150000 ;
        RECT 1110.000000 379.850000 1115.000000 380.150000 ;
        RECT 1110.000000 343.850000 1115.000000 344.150000 ;
        RECT 1110.000000 347.850000 1115.000000 348.150000 ;
        RECT 1110.000000 351.850000 1115.000000 352.150000 ;
        RECT 1110.000000 359.850000 1115.000000 360.150000 ;
        RECT 1110.000000 355.850000 1115.000000 356.150000 ;
        RECT 1110.000000 375.850000 1115.000000 376.150000 ;
        RECT 1110.000000 371.850000 1115.000000 372.150000 ;
        RECT 1110.000000 367.850000 1115.000000 368.150000 ;
        RECT 1110.000000 363.850000 1115.000000 364.150000 ;
        RECT 1110.000000 383.850000 1115.000000 384.150000 ;
        RECT 1110.000000 387.850000 1115.000000 388.150000 ;
        RECT 1110.000000 391.850000 1115.000000 392.150000 ;
        RECT 1110.000000 395.850000 1115.000000 396.150000 ;
        RECT 1110.000000 407.850000 1115.000000 408.150000 ;
        RECT 1110.000000 399.850000 1115.000000 400.150000 ;
        RECT 1110.000000 403.850000 1115.000000 404.150000 ;
        RECT 1110.000000 411.850000 1115.000000 412.150000 ;
        RECT 1110.000000 415.850000 1115.000000 416.150000 ;
        RECT 1060.000000 379.850000 1065.000000 380.150000 ;
        RECT 1060.000000 343.850000 1065.000000 344.150000 ;
        RECT 1060.000000 347.850000 1065.000000 348.150000 ;
        RECT 1060.000000 351.850000 1065.000000 352.150000 ;
        RECT 1060.000000 355.850000 1065.000000 356.150000 ;
        RECT 1060.000000 359.850000 1065.000000 360.150000 ;
        RECT 1060.000000 375.850000 1065.000000 376.150000 ;
        RECT 1060.000000 371.850000 1065.000000 372.150000 ;
        RECT 1060.000000 367.850000 1065.000000 368.150000 ;
        RECT 1060.000000 363.850000 1065.000000 364.150000 ;
        RECT 1060.000000 383.850000 1065.000000 384.150000 ;
        RECT 1060.000000 387.850000 1065.000000 388.150000 ;
        RECT 1060.000000 391.850000 1065.000000 392.150000 ;
        RECT 1060.000000 395.850000 1065.000000 396.150000 ;
        RECT 1060.000000 407.850000 1065.000000 408.150000 ;
        RECT 1060.000000 399.850000 1065.000000 400.150000 ;
        RECT 1060.000000 403.850000 1065.000000 404.150000 ;
        RECT 1060.000000 411.850000 1065.000000 412.150000 ;
        RECT 1060.000000 415.850000 1065.000000 416.150000 ;
        RECT 1158.000000 379.850000 1168.000000 380.150000 ;
        RECT 1158.000000 343.850000 1168.000000 344.150000 ;
        RECT 1158.000000 347.850000 1168.000000 348.150000 ;
        RECT 1158.000000 351.850000 1168.000000 352.150000 ;
        RECT 1158.000000 355.850000 1168.000000 356.150000 ;
        RECT 1158.000000 359.850000 1168.000000 360.150000 ;
        RECT 1158.000000 375.850000 1168.000000 376.150000 ;
        RECT 1158.000000 371.850000 1168.000000 372.150000 ;
        RECT 1158.000000 367.850000 1168.000000 368.150000 ;
        RECT 1158.000000 363.850000 1168.000000 364.150000 ;
        RECT 1158.000000 383.850000 1168.000000 384.150000 ;
        RECT 1158.000000 387.850000 1168.000000 388.150000 ;
        RECT 1158.000000 391.850000 1168.000000 392.150000 ;
        RECT 1158.000000 395.850000 1168.000000 396.150000 ;
        RECT 1158.000000 407.850000 1168.000000 408.150000 ;
        RECT 1158.000000 399.850000 1168.000000 400.150000 ;
        RECT 1158.000000 403.850000 1168.000000 404.150000 ;
        RECT 1158.000000 411.850000 1168.000000 412.150000 ;
        RECT 1158.000000 415.850000 1168.000000 416.150000 ;
        RECT 1110.000000 431.850000 1115.000000 432.150000 ;
        RECT 1110.000000 427.850000 1115.000000 428.150000 ;
        RECT 1110.000000 423.850000 1115.000000 424.150000 ;
        RECT 1110.000000 419.850000 1115.000000 420.150000 ;
        RECT 1110.000000 443.850000 1115.000000 444.150000 ;
        RECT 1110.000000 439.850000 1115.000000 440.150000 ;
        RECT 1110.000000 435.850000 1115.000000 436.150000 ;
        RECT 1060.000000 419.850000 1065.000000 420.150000 ;
        RECT 1060.000000 423.850000 1065.000000 424.150000 ;
        RECT 1060.000000 431.850000 1065.000000 432.150000 ;
        RECT 1060.000000 427.850000 1065.000000 428.150000 ;
        RECT 1060.000000 435.850000 1065.000000 436.150000 ;
        RECT 1060.000000 439.850000 1065.000000 440.150000 ;
        RECT 1060.000000 443.850000 1065.000000 444.150000 ;
        RECT 1158.000000 427.850000 1168.000000 428.150000 ;
        RECT 1158.000000 423.850000 1168.000000 424.150000 ;
        RECT 1158.000000 419.850000 1168.000000 420.150000 ;
        RECT 1160.000000 431.850000 1165.000000 432.150000 ;
        RECT 1160.000000 435.850000 1165.000000 436.150000 ;
        RECT 1160.000000 439.850000 1165.000000 440.150000 ;
        RECT 1160.000000 443.850000 1165.000000 444.150000 ;
        RECT 1160.000000 447.850000 1165.000000 448.150000 ;
        RECT 1160.000000 451.850000 1165.000000 452.150000 ;
        RECT 1160.000000 459.850000 1165.000000 460.150000 ;
        RECT 1160.000000 455.850000 1165.000000 456.150000 ;
        RECT 1160.000000 463.850000 1165.000000 464.150000 ;
        RECT 1160.000000 467.850000 1165.000000 468.150000 ;
        RECT 1160.000000 471.850000 1165.000000 472.150000 ;
        RECT 1160.000000 479.850000 1165.000000 480.150000 ;
        RECT 1160.000000 475.850000 1165.000000 476.150000 ;
        RECT 1160.000000 487.850000 1165.000000 488.150000 ;
        RECT 1160.000000 483.850000 1165.000000 484.150000 ;
        RECT 1160.000000 491.850000 1165.000000 492.150000 ;
        RECT 1160.000000 495.850000 1165.000000 496.150000 ;
        RECT 1160.000000 499.850000 1165.000000 500.150000 ;
        RECT 1160.000000 507.850000 1165.000000 508.150000 ;
        RECT 1160.000000 503.850000 1165.000000 504.150000 ;
        RECT 1160.000000 511.850000 1165.000000 512.150000 ;
        RECT 1160.000000 515.850000 1165.000000 516.150000 ;
        RECT 1160.000000 519.850000 1165.000000 520.150000 ;
        RECT 1160.000000 523.850000 1165.000000 524.150000 ;
        RECT 1160.000000 527.850000 1165.000000 528.150000 ;
        RECT 1160.000000 535.850000 1165.000000 536.150000 ;
        RECT 1160.000000 531.850000 1165.000000 532.150000 ;
        RECT 1160.000000 539.850000 1165.000000 540.150000 ;
        RECT 1160.000000 543.850000 1165.000000 544.150000 ;
        RECT 1160.000000 555.850000 1165.000000 556.150000 ;
        RECT 1160.000000 551.850000 1165.000000 552.150000 ;
        RECT 1160.000000 547.850000 1165.000000 548.150000 ;
        RECT 1160.000000 563.850000 1165.000000 564.150000 ;
        RECT 1160.000000 559.850000 1165.000000 560.150000 ;
        RECT 1160.000000 583.850000 1165.000000 584.150000 ;
        RECT 1160.000000 567.850000 1165.000000 568.150000 ;
        RECT 1160.000000 571.850000 1165.000000 572.150000 ;
        RECT 1160.000000 579.850000 1165.000000 580.150000 ;
        RECT 1160.000000 575.850000 1165.000000 576.150000 ;
        RECT 1160.000000 591.850000 1165.000000 592.150000 ;
        RECT 1160.000000 587.850000 1165.000000 588.150000 ;
        RECT 1160.000000 595.850000 1165.000000 596.150000 ;
        RECT 1160.000000 599.850000 1165.000000 600.150000 ;
        RECT 1160.000000 607.850000 1165.000000 608.150000 ;
        RECT 1160.000000 603.850000 1165.000000 604.150000 ;
        RECT 1160.000000 611.850000 1165.000000 612.150000 ;
        RECT 1160.000000 615.850000 1165.000000 616.150000 ;
        RECT 1160.000000 619.850000 1165.000000 620.150000 ;
        RECT 1160.000000 623.850000 1165.000000 624.150000 ;
        RECT 1160.000000 627.850000 1165.000000 628.150000 ;
        RECT 1160.000000 635.850000 1165.000000 636.150000 ;
        RECT 1160.000000 631.850000 1165.000000 632.150000 ;
        RECT 610.000000 659.850000 615.000000 660.150000 ;
        RECT 610.000000 663.850000 615.000000 664.150000 ;
        RECT 610.000000 667.850000 615.000000 668.150000 ;
        RECT 610.000000 671.850000 615.000000 672.150000 ;
        RECT 610.000000 675.850000 615.000000 676.150000 ;
        RECT 660.000000 663.850000 665.000000 664.150000 ;
        RECT 660.000000 659.850000 665.000000 660.150000 ;
        RECT 660.000000 667.850000 665.000000 668.150000 ;
        RECT 660.000000 671.850000 665.000000 672.150000 ;
        RECT 660.000000 675.850000 665.000000 676.150000 ;
        RECT 610.000000 683.850000 615.000000 684.150000 ;
        RECT 610.000000 679.850000 615.000000 680.150000 ;
        RECT 660.000000 683.850000 665.000000 684.150000 ;
        RECT 660.000000 679.850000 665.000000 680.150000 ;
        RECT 1160.000000 639.850000 1165.000000 640.150000 ;
        RECT 1160.000000 643.850000 1165.000000 644.150000 ;
        RECT 1160.000000 647.850000 1165.000000 648.150000 ;
        RECT 1160.000000 655.850000 1165.000000 656.150000 ;
        RECT 1160.000000 651.850000 1165.000000 652.150000 ;
        RECT 1160.000000 663.850000 1165.000000 664.150000 ;
        RECT 1160.000000 659.850000 1165.000000 660.150000 ;
        RECT 1160.000000 667.850000 1165.000000 668.150000 ;
        RECT 1160.000000 671.850000 1165.000000 672.150000 ;
        RECT 1160.000000 675.850000 1165.000000 676.150000 ;
        RECT 1160.000000 683.850000 1165.000000 684.150000 ;
        RECT 1160.000000 679.850000 1165.000000 680.150000 ;
      LAYER M3 ;
        RECT 60.000000 3.850000 65.000000 4.150000 ;
        RECT 60.000000 7.850000 65.000000 8.150000 ;
        RECT 110.000000 7.850000 115.000000 8.150000 ;
        RECT 110.000000 3.850000 115.000000 4.150000 ;
        RECT 160.000000 7.850000 165.000000 8.150000 ;
        RECT 160.000000 3.850000 165.000000 4.150000 ;
        RECT 210.000000 7.850000 215.000000 8.150000 ;
        RECT 210.000000 3.850000 215.000000 4.150000 ;
        RECT 260.000000 7.850000 265.000000 8.150000 ;
        RECT 260.000000 3.850000 265.000000 4.150000 ;
        RECT 310.000000 7.850000 315.000000 8.150000 ;
        RECT 310.000000 3.850000 315.000000 4.150000 ;
        RECT 360.000000 7.850000 365.000000 8.150000 ;
        RECT 360.000000 3.850000 365.000000 4.150000 ;
        RECT 410.000000 7.850000 415.000000 8.150000 ;
        RECT 410.000000 3.850000 415.000000 4.150000 ;
        RECT 460.000000 7.850000 465.000000 8.150000 ;
        RECT 460.000000 3.850000 465.000000 4.150000 ;
        RECT 510.000000 7.850000 515.000000 8.150000 ;
        RECT 510.000000 3.850000 515.000000 4.150000 ;
        RECT 560.000000 3.850000 565.000000 4.150000 ;
        RECT 560.000000 7.850000 565.000000 8.150000 ;
        RECT 18.000000 259.850000 28.000000 260.150000 ;
        RECT 18.000000 263.850000 28.000000 264.150000 ;
        RECT 18.000000 267.850000 28.000000 268.150000 ;
        RECT 60.000000 267.850000 65.000000 268.150000 ;
        RECT 60.000000 263.850000 65.000000 264.150000 ;
        RECT 60.000000 259.850000 65.000000 260.150000 ;
        RECT 110.000000 267.850000 115.000000 268.150000 ;
        RECT 110.000000 259.850000 115.000000 260.150000 ;
        RECT 110.000000 263.850000 115.000000 264.150000 ;
        RECT 18.000000 283.850000 28.000000 284.150000 ;
        RECT 18.000000 279.850000 28.000000 280.150000 ;
        RECT 18.000000 275.850000 28.000000 276.150000 ;
        RECT 18.000000 271.850000 28.000000 272.150000 ;
        RECT 18.000000 287.850000 28.000000 288.150000 ;
        RECT 18.000000 291.850000 28.000000 292.150000 ;
        RECT 18.000000 295.850000 28.000000 296.150000 ;
        RECT 18.000000 299.850000 28.000000 300.150000 ;
        RECT 18.000000 303.850000 28.000000 304.150000 ;
        RECT 60.000000 283.850000 65.000000 284.150000 ;
        RECT 60.000000 279.850000 65.000000 280.150000 ;
        RECT 60.000000 275.850000 65.000000 276.150000 ;
        RECT 60.000000 271.850000 65.000000 272.150000 ;
        RECT 60.000000 287.850000 65.000000 288.150000 ;
        RECT 60.000000 291.850000 65.000000 292.150000 ;
        RECT 60.000000 295.850000 65.000000 296.150000 ;
        RECT 60.000000 299.850000 65.000000 300.150000 ;
        RECT 60.000000 303.850000 65.000000 304.150000 ;
        RECT 18.000000 307.850000 28.000000 308.150000 ;
        RECT 18.000000 311.850000 28.000000 312.150000 ;
        RECT 18.000000 315.850000 28.000000 316.150000 ;
        RECT 18.000000 319.850000 28.000000 320.150000 ;
        RECT 18.000000 323.850000 28.000000 324.150000 ;
        RECT 18.000000 339.850000 28.000000 340.150000 ;
        RECT 18.000000 335.850000 28.000000 336.150000 ;
        RECT 18.000000 331.850000 28.000000 332.150000 ;
        RECT 18.000000 327.850000 28.000000 328.150000 ;
        RECT 60.000000 307.850000 65.000000 308.150000 ;
        RECT 60.000000 311.850000 65.000000 312.150000 ;
        RECT 60.000000 315.850000 65.000000 316.150000 ;
        RECT 60.000000 319.850000 65.000000 320.150000 ;
        RECT 60.000000 323.850000 65.000000 324.150000 ;
        RECT 60.000000 339.850000 65.000000 340.150000 ;
        RECT 60.000000 335.850000 65.000000 336.150000 ;
        RECT 60.000000 331.850000 65.000000 332.150000 ;
        RECT 60.000000 327.850000 65.000000 328.150000 ;
        RECT 110.000000 271.850000 115.000000 272.150000 ;
        RECT 110.000000 275.850000 115.000000 276.150000 ;
        RECT 110.000000 279.850000 115.000000 280.150000 ;
        RECT 110.000000 283.850000 115.000000 284.150000 ;
        RECT 110.000000 287.850000 115.000000 288.150000 ;
        RECT 110.000000 291.850000 115.000000 292.150000 ;
        RECT 110.000000 295.850000 115.000000 296.150000 ;
        RECT 110.000000 299.850000 115.000000 300.150000 ;
        RECT 110.000000 303.850000 115.000000 304.150000 ;
        RECT 110.000000 311.850000 115.000000 312.150000 ;
        RECT 110.000000 307.850000 115.000000 308.150000 ;
        RECT 110.000000 323.850000 115.000000 324.150000 ;
        RECT 110.000000 319.850000 115.000000 320.150000 ;
        RECT 110.000000 315.850000 115.000000 316.150000 ;
        RECT 110.000000 339.850000 115.000000 340.150000 ;
        RECT 110.000000 335.850000 115.000000 336.150000 ;
        RECT 110.000000 331.850000 115.000000 332.150000 ;
        RECT 110.000000 327.850000 115.000000 328.150000 ;
        RECT 160.000000 259.850000 165.000000 260.150000 ;
        RECT 160.000000 263.850000 165.000000 264.150000 ;
        RECT 160.000000 267.850000 165.000000 268.150000 ;
        RECT 210.000000 267.850000 215.000000 268.150000 ;
        RECT 210.000000 263.850000 215.000000 264.150000 ;
        RECT 210.000000 259.850000 215.000000 260.150000 ;
        RECT 260.000000 267.850000 265.000000 268.150000 ;
        RECT 260.000000 259.850000 265.000000 260.150000 ;
        RECT 260.000000 263.850000 265.000000 264.150000 ;
        RECT 160.000000 275.850000 165.000000 276.150000 ;
        RECT 160.000000 271.850000 165.000000 272.150000 ;
        RECT 160.000000 283.850000 165.000000 284.150000 ;
        RECT 160.000000 279.850000 165.000000 280.150000 ;
        RECT 160.000000 287.850000 165.000000 288.150000 ;
        RECT 160.000000 291.850000 165.000000 292.150000 ;
        RECT 160.000000 295.850000 165.000000 296.150000 ;
        RECT 160.000000 303.850000 165.000000 304.150000 ;
        RECT 160.000000 299.850000 165.000000 300.150000 ;
        RECT 210.000000 271.850000 215.000000 272.150000 ;
        RECT 210.000000 275.850000 215.000000 276.150000 ;
        RECT 210.000000 279.850000 215.000000 280.150000 ;
        RECT 210.000000 283.850000 215.000000 284.150000 ;
        RECT 210.000000 287.850000 215.000000 288.150000 ;
        RECT 210.000000 291.850000 215.000000 292.150000 ;
        RECT 210.000000 295.850000 215.000000 296.150000 ;
        RECT 210.000000 299.850000 215.000000 300.150000 ;
        RECT 210.000000 303.850000 215.000000 304.150000 ;
        RECT 160.000000 311.850000 165.000000 312.150000 ;
        RECT 160.000000 307.850000 165.000000 308.150000 ;
        RECT 160.000000 315.850000 165.000000 316.150000 ;
        RECT 160.000000 319.850000 165.000000 320.150000 ;
        RECT 160.000000 323.850000 165.000000 324.150000 ;
        RECT 160.000000 331.850000 165.000000 332.150000 ;
        RECT 160.000000 327.850000 165.000000 328.150000 ;
        RECT 160.000000 335.850000 165.000000 336.150000 ;
        RECT 160.000000 339.850000 165.000000 340.150000 ;
        RECT 210.000000 307.850000 215.000000 308.150000 ;
        RECT 210.000000 311.850000 215.000000 312.150000 ;
        RECT 210.000000 315.850000 215.000000 316.150000 ;
        RECT 210.000000 319.850000 215.000000 320.150000 ;
        RECT 210.000000 323.850000 215.000000 324.150000 ;
        RECT 210.000000 327.850000 215.000000 328.150000 ;
        RECT 210.000000 331.850000 215.000000 332.150000 ;
        RECT 210.000000 335.850000 215.000000 336.150000 ;
        RECT 210.000000 339.850000 215.000000 340.150000 ;
        RECT 260.000000 271.850000 265.000000 272.150000 ;
        RECT 260.000000 275.850000 265.000000 276.150000 ;
        RECT 260.000000 279.850000 265.000000 280.150000 ;
        RECT 260.000000 283.850000 265.000000 284.150000 ;
        RECT 260.000000 295.850000 265.000000 296.150000 ;
        RECT 260.000000 291.850000 265.000000 292.150000 ;
        RECT 260.000000 287.850000 265.000000 288.150000 ;
        RECT 260.000000 303.850000 265.000000 304.150000 ;
        RECT 260.000000 299.850000 265.000000 300.150000 ;
        RECT 260.000000 323.850000 265.000000 324.150000 ;
        RECT 260.000000 319.850000 265.000000 320.150000 ;
        RECT 260.000000 315.850000 265.000000 316.150000 ;
        RECT 260.000000 311.850000 265.000000 312.150000 ;
        RECT 260.000000 307.850000 265.000000 308.150000 ;
        RECT 260.000000 327.850000 265.000000 328.150000 ;
        RECT 260.000000 331.850000 265.000000 332.150000 ;
        RECT 260.000000 335.850000 265.000000 336.150000 ;
        RECT 260.000000 339.850000 265.000000 340.150000 ;
        RECT 310.000000 263.850000 315.000000 264.150000 ;
        RECT 310.000000 259.850000 315.000000 260.150000 ;
        RECT 310.000000 267.850000 315.000000 268.150000 ;
        RECT 360.000000 259.850000 365.000000 260.150000 ;
        RECT 360.000000 263.850000 365.000000 264.150000 ;
        RECT 360.000000 267.850000 365.000000 268.150000 ;
        RECT 410.000000 259.850000 415.000000 260.150000 ;
        RECT 410.000000 263.850000 415.000000 264.150000 ;
        RECT 410.000000 267.850000 415.000000 268.150000 ;
        RECT 310.000000 275.850000 315.000000 276.150000 ;
        RECT 310.000000 271.850000 315.000000 272.150000 ;
        RECT 310.000000 279.850000 315.000000 280.150000 ;
        RECT 310.000000 283.850000 315.000000 284.150000 ;
        RECT 310.000000 287.850000 315.000000 288.150000 ;
        RECT 310.000000 291.850000 315.000000 292.150000 ;
        RECT 310.000000 295.850000 315.000000 296.150000 ;
        RECT 310.000000 303.850000 315.000000 304.150000 ;
        RECT 310.000000 299.850000 315.000000 300.150000 ;
        RECT 360.000000 283.850000 365.000000 284.150000 ;
        RECT 360.000000 279.850000 365.000000 280.150000 ;
        RECT 360.000000 275.850000 365.000000 276.150000 ;
        RECT 360.000000 271.850000 365.000000 272.150000 ;
        RECT 360.000000 287.850000 365.000000 288.150000 ;
        RECT 360.000000 291.850000 365.000000 292.150000 ;
        RECT 360.000000 295.850000 365.000000 296.150000 ;
        RECT 360.000000 299.850000 365.000000 300.150000 ;
        RECT 360.000000 303.850000 365.000000 304.150000 ;
        RECT 310.000000 311.850000 315.000000 312.150000 ;
        RECT 310.000000 307.850000 315.000000 308.150000 ;
        RECT 310.000000 315.850000 315.000000 316.150000 ;
        RECT 310.000000 319.850000 315.000000 320.150000 ;
        RECT 310.000000 323.850000 315.000000 324.150000 ;
        RECT 310.000000 327.850000 315.000000 328.150000 ;
        RECT 310.000000 331.850000 315.000000 332.150000 ;
        RECT 310.000000 335.850000 315.000000 336.150000 ;
        RECT 310.000000 339.850000 315.000000 340.150000 ;
        RECT 360.000000 307.850000 365.000000 308.150000 ;
        RECT 360.000000 311.850000 365.000000 312.150000 ;
        RECT 360.000000 315.850000 365.000000 316.150000 ;
        RECT 360.000000 319.850000 365.000000 320.150000 ;
        RECT 360.000000 323.850000 365.000000 324.150000 ;
        RECT 360.000000 327.850000 365.000000 328.150000 ;
        RECT 360.000000 331.850000 365.000000 332.150000 ;
        RECT 360.000000 335.850000 365.000000 336.150000 ;
        RECT 360.000000 339.850000 365.000000 340.150000 ;
        RECT 410.000000 271.850000 415.000000 272.150000 ;
        RECT 410.000000 275.850000 415.000000 276.150000 ;
        RECT 410.000000 283.850000 415.000000 284.150000 ;
        RECT 410.000000 279.850000 415.000000 280.150000 ;
        RECT 410.000000 295.850000 415.000000 296.150000 ;
        RECT 410.000000 291.850000 415.000000 292.150000 ;
        RECT 410.000000 287.850000 415.000000 288.150000 ;
        RECT 410.000000 299.850000 415.000000 300.150000 ;
        RECT 410.000000 303.850000 415.000000 304.150000 ;
        RECT 410.000000 323.850000 415.000000 324.150000 ;
        RECT 410.000000 319.850000 415.000000 320.150000 ;
        RECT 410.000000 315.850000 415.000000 316.150000 ;
        RECT 410.000000 311.850000 415.000000 312.150000 ;
        RECT 410.000000 307.850000 415.000000 308.150000 ;
        RECT 410.000000 327.850000 415.000000 328.150000 ;
        RECT 410.000000 331.850000 415.000000 332.150000 ;
        RECT 410.000000 335.850000 415.000000 336.150000 ;
        RECT 410.000000 339.850000 415.000000 340.150000 ;
        RECT 460.000000 259.850000 465.000000 260.150000 ;
        RECT 460.000000 263.850000 465.000000 264.150000 ;
        RECT 460.000000 267.850000 465.000000 268.150000 ;
        RECT 510.000000 259.850000 515.000000 260.150000 ;
        RECT 510.000000 263.850000 515.000000 264.150000 ;
        RECT 510.000000 267.850000 515.000000 268.150000 ;
        RECT 560.000000 263.850000 565.000000 264.150000 ;
        RECT 560.000000 259.850000 565.000000 260.150000 ;
        RECT 560.000000 267.850000 565.000000 268.150000 ;
        RECT 460.000000 283.850000 465.000000 284.150000 ;
        RECT 460.000000 279.850000 465.000000 280.150000 ;
        RECT 460.000000 275.850000 465.000000 276.150000 ;
        RECT 460.000000 271.850000 465.000000 272.150000 ;
        RECT 460.000000 287.850000 465.000000 288.150000 ;
        RECT 460.000000 291.850000 465.000000 292.150000 ;
        RECT 460.000000 295.850000 465.000000 296.150000 ;
        RECT 460.000000 301.230000 465.000000 302.230000 ;
        RECT 510.000000 275.850000 515.000000 276.150000 ;
        RECT 510.000000 271.850000 515.000000 272.150000 ;
        RECT 510.000000 283.850000 515.000000 284.150000 ;
        RECT 510.000000 279.850000 515.000000 280.150000 ;
        RECT 510.000000 291.850000 515.000000 292.150000 ;
        RECT 510.000000 287.850000 515.000000 288.150000 ;
        RECT 510.000000 295.850000 515.000000 296.150000 ;
        RECT 510.000000 303.850000 515.000000 304.150000 ;
        RECT 510.000000 299.850000 515.000000 300.150000 ;
        RECT 460.000000 319.850000 465.000000 320.150000 ;
        RECT 460.000000 323.850000 465.000000 324.150000 ;
        RECT 460.000000 339.850000 465.000000 340.150000 ;
        RECT 460.000000 335.850000 465.000000 336.150000 ;
        RECT 460.000000 331.850000 465.000000 332.150000 ;
        RECT 460.000000 327.850000 465.000000 328.150000 ;
        RECT 510.000000 311.850000 515.000000 312.150000 ;
        RECT 510.000000 307.850000 515.000000 308.150000 ;
        RECT 510.000000 315.850000 515.000000 316.150000 ;
        RECT 510.000000 319.850000 515.000000 320.150000 ;
        RECT 510.000000 323.850000 515.000000 324.150000 ;
        RECT 510.000000 331.850000 515.000000 332.150000 ;
        RECT 510.000000 327.850000 515.000000 328.150000 ;
        RECT 510.000000 335.850000 515.000000 336.150000 ;
        RECT 510.000000 339.850000 515.000000 340.150000 ;
        RECT 560.000000 271.850000 565.000000 272.150000 ;
        RECT 560.000000 275.850000 565.000000 276.150000 ;
        RECT 560.000000 279.850000 565.000000 280.150000 ;
        RECT 560.000000 283.850000 565.000000 284.150000 ;
        RECT 560.000000 291.850000 565.000000 292.150000 ;
        RECT 560.000000 287.850000 565.000000 288.150000 ;
        RECT 560.000000 295.850000 565.000000 296.150000 ;
        RECT 560.000000 303.850000 565.000000 304.150000 ;
        RECT 560.000000 299.850000 565.000000 300.150000 ;
        RECT 560.000000 323.850000 565.000000 324.150000 ;
        RECT 560.000000 319.850000 565.000000 320.150000 ;
        RECT 560.000000 315.850000 565.000000 316.150000 ;
        RECT 560.000000 311.850000 565.000000 312.150000 ;
        RECT 560.000000 307.850000 565.000000 308.150000 ;
        RECT 560.000000 339.850000 565.000000 340.150000 ;
        RECT 560.000000 335.850000 565.000000 336.150000 ;
        RECT 560.000000 331.850000 565.000000 332.150000 ;
        RECT 560.000000 327.850000 565.000000 328.150000 ;
        RECT 610.000000 3.850000 615.000000 4.150000 ;
        RECT 610.000000 7.850000 615.000000 8.150000 ;
        RECT 660.000000 7.850000 665.000000 8.150000 ;
        RECT 660.000000 3.850000 665.000000 4.150000 ;
        RECT 710.000000 7.850000 715.000000 8.150000 ;
        RECT 710.000000 3.850000 715.000000 4.150000 ;
        RECT 760.000000 7.850000 765.000000 8.150000 ;
        RECT 760.000000 3.850000 765.000000 4.150000 ;
        RECT 810.000000 7.850000 815.000000 8.150000 ;
        RECT 810.000000 3.850000 815.000000 4.150000 ;
        RECT 860.000000 7.850000 865.000000 8.150000 ;
        RECT 860.000000 3.850000 865.000000 4.150000 ;
        RECT 960.000000 7.850000 965.000000 8.150000 ;
        RECT 960.000000 3.850000 965.000000 4.150000 ;
        RECT 910.000000 7.850000 915.000000 8.150000 ;
        RECT 910.000000 3.850000 915.000000 4.150000 ;
        RECT 1010.000000 7.850000 1015.000000 8.150000 ;
        RECT 1010.000000 3.850000 1015.000000 4.150000 ;
        RECT 1110.000000 7.850000 1115.000000 8.150000 ;
        RECT 1110.000000 3.850000 1115.000000 4.150000 ;
        RECT 1060.000000 7.850000 1065.000000 8.150000 ;
        RECT 1060.000000 3.850000 1065.000000 4.150000 ;
        RECT 1160.000000 3.850000 1165.000000 4.150000 ;
        RECT 1160.000000 7.850000 1165.000000 8.150000 ;
        RECT 1158.000000 27.850000 1168.000000 28.150000 ;
        RECT 1158.000000 23.850000 1168.000000 24.150000 ;
        RECT 1158.000000 19.850000 1168.000000 20.150000 ;
        RECT 1160.000000 15.850000 1165.000000 16.150000 ;
        RECT 1160.000000 11.850000 1165.000000 12.150000 ;
        RECT 1158.000000 31.850000 1168.000000 32.150000 ;
        RECT 1158.000000 35.850000 1168.000000 36.150000 ;
        RECT 1158.000000 43.850000 1168.000000 44.150000 ;
        RECT 1158.000000 39.850000 1168.000000 40.150000 ;
        RECT 610.000000 263.850000 615.000000 264.150000 ;
        RECT 610.000000 259.850000 615.000000 260.150000 ;
        RECT 610.000000 267.850000 615.000000 268.150000 ;
        RECT 660.000000 259.850000 665.000000 260.150000 ;
        RECT 660.000000 263.850000 665.000000 264.150000 ;
        RECT 660.000000 267.850000 665.000000 268.150000 ;
        RECT 710.000000 267.850000 715.000000 268.150000 ;
        RECT 710.000000 259.850000 715.000000 260.150000 ;
        RECT 710.000000 263.850000 715.000000 264.150000 ;
        RECT 610.000000 283.850000 615.000000 284.150000 ;
        RECT 610.000000 279.850000 615.000000 280.150000 ;
        RECT 610.000000 275.850000 615.000000 276.150000 ;
        RECT 610.000000 271.850000 615.000000 272.150000 ;
        RECT 610.000000 287.850000 615.000000 288.150000 ;
        RECT 610.000000 291.850000 615.000000 292.150000 ;
        RECT 610.000000 295.850000 615.000000 296.150000 ;
        RECT 610.000000 299.850000 615.000000 300.150000 ;
        RECT 610.000000 303.850000 615.000000 304.150000 ;
        RECT 660.000000 275.850000 665.000000 276.150000 ;
        RECT 660.000000 271.850000 665.000000 272.150000 ;
        RECT 660.000000 283.850000 665.000000 284.150000 ;
        RECT 660.000000 279.850000 665.000000 280.150000 ;
        RECT 660.000000 287.850000 665.000000 288.150000 ;
        RECT 660.000000 291.850000 665.000000 292.150000 ;
        RECT 660.000000 295.850000 665.000000 296.150000 ;
        RECT 660.000000 303.850000 665.000000 304.150000 ;
        RECT 660.000000 299.850000 665.000000 300.150000 ;
        RECT 610.000000 307.850000 615.000000 308.150000 ;
        RECT 610.000000 311.850000 615.000000 312.150000 ;
        RECT 610.000000 315.850000 615.000000 316.150000 ;
        RECT 610.000000 319.850000 615.000000 320.150000 ;
        RECT 610.000000 323.850000 615.000000 324.150000 ;
        RECT 610.000000 339.850000 615.000000 340.150000 ;
        RECT 610.000000 335.850000 615.000000 336.150000 ;
        RECT 610.000000 331.850000 615.000000 332.150000 ;
        RECT 610.000000 327.850000 615.000000 328.150000 ;
        RECT 660.000000 311.850000 665.000000 312.150000 ;
        RECT 660.000000 307.850000 665.000000 308.150000 ;
        RECT 660.000000 315.850000 665.000000 316.150000 ;
        RECT 660.000000 319.850000 665.000000 320.150000 ;
        RECT 660.000000 323.850000 665.000000 324.150000 ;
        RECT 660.000000 331.850000 665.000000 332.150000 ;
        RECT 660.000000 327.850000 665.000000 328.150000 ;
        RECT 660.000000 335.850000 665.000000 336.150000 ;
        RECT 660.000000 339.850000 665.000000 340.150000 ;
        RECT 710.000000 271.850000 715.000000 272.150000 ;
        RECT 710.000000 275.850000 715.000000 276.150000 ;
        RECT 710.000000 279.850000 715.000000 280.150000 ;
        RECT 710.000000 283.850000 715.000000 284.150000 ;
        RECT 710.000000 287.850000 715.000000 288.150000 ;
        RECT 710.000000 291.850000 715.000000 292.150000 ;
        RECT 710.000000 295.850000 715.000000 296.150000 ;
        RECT 710.000000 299.850000 715.000000 300.150000 ;
        RECT 710.000000 303.850000 715.000000 304.150000 ;
        RECT 710.000000 323.850000 715.000000 324.150000 ;
        RECT 710.000000 319.850000 715.000000 320.150000 ;
        RECT 710.000000 315.850000 715.000000 316.150000 ;
        RECT 710.000000 311.850000 715.000000 312.150000 ;
        RECT 710.000000 307.850000 715.000000 308.150000 ;
        RECT 710.000000 339.850000 715.000000 340.150000 ;
        RECT 710.000000 335.850000 715.000000 336.150000 ;
        RECT 710.000000 331.850000 715.000000 332.150000 ;
        RECT 710.000000 327.850000 715.000000 328.150000 ;
        RECT 760.000000 267.850000 765.000000 268.150000 ;
        RECT 760.000000 263.850000 765.000000 264.150000 ;
        RECT 760.000000 259.850000 765.000000 260.150000 ;
        RECT 810.000000 259.850000 815.000000 260.150000 ;
        RECT 810.000000 263.850000 815.000000 264.150000 ;
        RECT 810.000000 267.850000 815.000000 268.150000 ;
        RECT 860.000000 267.850000 865.000000 268.150000 ;
        RECT 860.000000 259.850000 865.000000 260.150000 ;
        RECT 860.000000 263.850000 865.000000 264.150000 ;
        RECT 760.000000 283.850000 765.000000 284.150000 ;
        RECT 760.000000 279.850000 765.000000 280.150000 ;
        RECT 760.000000 275.850000 765.000000 276.150000 ;
        RECT 760.000000 271.850000 765.000000 272.150000 ;
        RECT 760.000000 287.850000 765.000000 288.150000 ;
        RECT 760.000000 291.850000 765.000000 292.150000 ;
        RECT 760.000000 295.850000 765.000000 296.150000 ;
        RECT 760.000000 299.850000 765.000000 300.150000 ;
        RECT 760.000000 303.850000 765.000000 304.150000 ;
        RECT 810.000000 275.850000 815.000000 276.150000 ;
        RECT 810.000000 271.850000 815.000000 272.150000 ;
        RECT 810.000000 283.850000 815.000000 284.150000 ;
        RECT 810.000000 279.850000 815.000000 280.150000 ;
        RECT 810.000000 287.850000 815.000000 288.150000 ;
        RECT 810.000000 291.850000 815.000000 292.150000 ;
        RECT 810.000000 295.850000 815.000000 296.150000 ;
        RECT 810.000000 303.850000 815.000000 304.150000 ;
        RECT 810.000000 299.850000 815.000000 300.150000 ;
        RECT 760.000000 307.850000 765.000000 308.150000 ;
        RECT 760.000000 311.850000 765.000000 312.150000 ;
        RECT 760.000000 315.850000 765.000000 316.150000 ;
        RECT 760.000000 319.850000 765.000000 320.150000 ;
        RECT 760.000000 323.850000 765.000000 324.150000 ;
        RECT 760.000000 339.850000 765.000000 340.150000 ;
        RECT 760.000000 335.850000 765.000000 336.150000 ;
        RECT 760.000000 331.850000 765.000000 332.150000 ;
        RECT 760.000000 327.850000 765.000000 328.150000 ;
        RECT 810.000000 311.850000 815.000000 312.150000 ;
        RECT 810.000000 307.850000 815.000000 308.150000 ;
        RECT 810.000000 315.850000 815.000000 316.150000 ;
        RECT 810.000000 319.850000 815.000000 320.150000 ;
        RECT 810.000000 323.850000 815.000000 324.150000 ;
        RECT 810.000000 331.850000 815.000000 332.150000 ;
        RECT 810.000000 327.850000 815.000000 328.150000 ;
        RECT 810.000000 335.850000 815.000000 336.150000 ;
        RECT 810.000000 339.850000 815.000000 340.150000 ;
        RECT 860.000000 271.850000 865.000000 272.150000 ;
        RECT 860.000000 275.850000 865.000000 276.150000 ;
        RECT 860.000000 279.850000 865.000000 280.150000 ;
        RECT 860.000000 283.850000 865.000000 284.150000 ;
        RECT 860.000000 287.850000 865.000000 288.150000 ;
        RECT 860.000000 291.850000 865.000000 292.150000 ;
        RECT 860.000000 295.850000 865.000000 296.150000 ;
        RECT 860.000000 299.850000 865.000000 300.150000 ;
        RECT 860.000000 303.850000 865.000000 304.150000 ;
        RECT 860.000000 323.850000 865.000000 324.150000 ;
        RECT 860.000000 319.850000 865.000000 320.150000 ;
        RECT 860.000000 315.850000 865.000000 316.150000 ;
        RECT 860.000000 311.850000 865.000000 312.150000 ;
        RECT 860.000000 307.850000 865.000000 308.150000 ;
        RECT 860.000000 339.850000 865.000000 340.150000 ;
        RECT 860.000000 335.850000 865.000000 336.150000 ;
        RECT 860.000000 331.850000 865.000000 332.150000 ;
        RECT 860.000000 327.850000 865.000000 328.150000 ;
        RECT 1158.000000 47.850000 1168.000000 48.150000 ;
        RECT 1158.000000 51.850000 1168.000000 52.150000 ;
        RECT 1158.000000 63.850000 1168.000000 64.150000 ;
        RECT 1158.000000 55.850000 1168.000000 56.150000 ;
        RECT 1158.000000 59.850000 1168.000000 60.150000 ;
        RECT 1158.000000 67.850000 1168.000000 68.150000 ;
        RECT 1158.000000 71.850000 1168.000000 72.150000 ;
        RECT 1158.000000 79.850000 1168.000000 80.150000 ;
        RECT 1158.000000 75.850000 1168.000000 76.150000 ;
        RECT 1158.000000 83.850000 1168.000000 84.150000 ;
        RECT 1158.000000 87.850000 1168.000000 88.150000 ;
        RECT 1158.000000 91.850000 1168.000000 92.150000 ;
        RECT 1158.000000 99.850000 1168.000000 100.150000 ;
        RECT 1158.000000 95.850000 1168.000000 96.150000 ;
        RECT 1158.000000 103.850000 1168.000000 104.150000 ;
        RECT 1158.000000 107.850000 1168.000000 108.150000 ;
        RECT 1158.000000 119.850000 1168.000000 120.150000 ;
        RECT 1158.000000 115.850000 1168.000000 116.150000 ;
        RECT 1158.000000 111.850000 1168.000000 112.150000 ;
        RECT 1158.000000 123.850000 1168.000000 124.150000 ;
        RECT 1158.000000 127.850000 1168.000000 128.150000 ;
        RECT 1158.000000 135.850000 1168.000000 136.150000 ;
        RECT 1158.000000 131.850000 1168.000000 132.150000 ;
        RECT 1158.000000 139.850000 1168.000000 140.150000 ;
        RECT 1158.000000 143.850000 1168.000000 144.150000 ;
        RECT 1158.000000 147.850000 1168.000000 148.150000 ;
        RECT 1158.000000 155.850000 1168.000000 156.150000 ;
        RECT 1158.000000 151.850000 1168.000000 152.150000 ;
        RECT 1158.000000 159.850000 1168.000000 160.150000 ;
        RECT 1158.000000 163.850000 1168.000000 164.150000 ;
        RECT 1158.000000 175.850000 1168.000000 176.150000 ;
        RECT 1158.000000 171.850000 1168.000000 172.150000 ;
        RECT 1158.000000 167.850000 1168.000000 168.150000 ;
        RECT 1158.000000 179.850000 1168.000000 180.150000 ;
        RECT 1158.000000 183.850000 1168.000000 184.150000 ;
        RECT 1158.000000 191.850000 1168.000000 192.150000 ;
        RECT 1158.000000 187.850000 1168.000000 188.150000 ;
        RECT 960.000000 267.850000 965.000000 268.150000 ;
        RECT 960.000000 263.850000 965.000000 264.150000 ;
        RECT 960.000000 259.850000 965.000000 260.150000 ;
        RECT 910.000000 267.850000 915.000000 268.150000 ;
        RECT 910.000000 263.850000 915.000000 264.150000 ;
        RECT 910.000000 259.850000 915.000000 260.150000 ;
        RECT 1010.000000 259.850000 1015.000000 260.150000 ;
        RECT 1010.000000 263.850000 1015.000000 264.150000 ;
        RECT 1010.000000 267.850000 1015.000000 268.150000 ;
        RECT 960.000000 283.850000 965.000000 284.150000 ;
        RECT 960.000000 279.850000 965.000000 280.150000 ;
        RECT 960.000000 275.850000 965.000000 276.150000 ;
        RECT 960.000000 271.850000 965.000000 272.150000 ;
        RECT 960.000000 287.850000 965.000000 288.150000 ;
        RECT 960.000000 291.850000 965.000000 292.150000 ;
        RECT 960.000000 295.850000 965.000000 296.150000 ;
        RECT 960.000000 299.850000 965.000000 300.150000 ;
        RECT 960.000000 303.850000 965.000000 304.150000 ;
        RECT 960.000000 311.850000 965.000000 312.150000 ;
        RECT 960.000000 307.850000 965.000000 308.150000 ;
        RECT 960.000000 323.850000 965.000000 324.150000 ;
        RECT 960.000000 319.850000 965.000000 320.150000 ;
        RECT 960.000000 315.850000 965.000000 316.150000 ;
        RECT 960.000000 339.850000 965.000000 340.150000 ;
        RECT 960.000000 335.850000 965.000000 336.150000 ;
        RECT 960.000000 331.850000 965.000000 332.150000 ;
        RECT 960.000000 327.850000 965.000000 328.150000 ;
        RECT 910.000000 283.850000 915.000000 284.150000 ;
        RECT 910.000000 279.850000 915.000000 280.150000 ;
        RECT 910.000000 275.850000 915.000000 276.150000 ;
        RECT 910.000000 271.850000 915.000000 272.150000 ;
        RECT 910.000000 287.850000 915.000000 288.150000 ;
        RECT 910.000000 291.850000 915.000000 292.150000 ;
        RECT 910.000000 295.850000 915.000000 296.150000 ;
        RECT 910.000000 299.850000 915.000000 300.150000 ;
        RECT 910.000000 303.850000 915.000000 304.150000 ;
        RECT 910.000000 307.850000 915.000000 308.150000 ;
        RECT 910.000000 311.850000 915.000000 312.150000 ;
        RECT 910.000000 315.850000 915.000000 316.150000 ;
        RECT 910.000000 319.850000 915.000000 320.150000 ;
        RECT 910.000000 323.850000 915.000000 324.150000 ;
        RECT 910.000000 339.850000 915.000000 340.150000 ;
        RECT 910.000000 335.850000 915.000000 336.150000 ;
        RECT 910.000000 331.850000 915.000000 332.150000 ;
        RECT 910.000000 327.850000 915.000000 328.150000 ;
        RECT 1010.000000 275.850000 1015.000000 276.150000 ;
        RECT 1010.000000 271.850000 1015.000000 272.150000 ;
        RECT 1010.000000 283.850000 1015.000000 284.150000 ;
        RECT 1010.000000 279.850000 1015.000000 280.150000 ;
        RECT 1010.000000 287.850000 1015.000000 288.150000 ;
        RECT 1010.000000 291.850000 1015.000000 292.150000 ;
        RECT 1010.000000 295.850000 1015.000000 296.150000 ;
        RECT 1010.000000 303.850000 1015.000000 304.150000 ;
        RECT 1010.000000 299.850000 1015.000000 300.150000 ;
        RECT 1010.000000 311.850000 1015.000000 312.150000 ;
        RECT 1010.000000 307.850000 1015.000000 308.150000 ;
        RECT 1010.000000 315.850000 1015.000000 316.150000 ;
        RECT 1010.000000 319.850000 1015.000000 320.150000 ;
        RECT 1010.000000 323.850000 1015.000000 324.150000 ;
        RECT 1010.000000 331.850000 1015.000000 332.150000 ;
        RECT 1010.000000 327.850000 1015.000000 328.150000 ;
        RECT 1010.000000 335.850000 1015.000000 336.150000 ;
        RECT 1010.000000 339.850000 1015.000000 340.150000 ;
        RECT 1110.000000 267.850000 1115.000000 268.150000 ;
        RECT 1110.000000 263.850000 1115.000000 264.150000 ;
        RECT 1110.000000 259.850000 1115.000000 260.150000 ;
        RECT 1060.000000 267.850000 1065.000000 268.150000 ;
        RECT 1060.000000 263.850000 1065.000000 264.150000 ;
        RECT 1060.000000 259.850000 1065.000000 260.150000 ;
        RECT 1158.000000 203.850000 1168.000000 204.150000 ;
        RECT 1158.000000 195.850000 1168.000000 196.150000 ;
        RECT 1158.000000 199.850000 1168.000000 200.150000 ;
        RECT 1158.000000 211.850000 1168.000000 212.150000 ;
        RECT 1158.000000 207.850000 1168.000000 208.150000 ;
        RECT 1158.000000 215.850000 1168.000000 216.150000 ;
        RECT 1158.000000 219.850000 1168.000000 220.150000 ;
        RECT 1158.000000 227.850000 1168.000000 228.150000 ;
        RECT 1158.000000 223.850000 1168.000000 224.150000 ;
        RECT 1158.000000 231.850000 1168.000000 232.150000 ;
        RECT 1158.000000 235.850000 1168.000000 236.150000 ;
        RECT 1158.000000 239.850000 1168.000000 240.150000 ;
        RECT 1158.000000 247.850000 1168.000000 248.150000 ;
        RECT 1158.000000 243.850000 1168.000000 244.150000 ;
        RECT 1158.000000 251.850000 1168.000000 252.150000 ;
        RECT 1158.000000 255.850000 1168.000000 256.150000 ;
        RECT 1158.000000 267.850000 1168.000000 268.150000 ;
        RECT 1158.000000 259.850000 1168.000000 260.150000 ;
        RECT 1158.000000 263.850000 1168.000000 264.150000 ;
        RECT 1110.000000 283.850000 1115.000000 284.150000 ;
        RECT 1110.000000 279.850000 1115.000000 280.150000 ;
        RECT 1110.000000 275.850000 1115.000000 276.150000 ;
        RECT 1110.000000 271.850000 1115.000000 272.150000 ;
        RECT 1110.000000 287.850000 1115.000000 288.150000 ;
        RECT 1110.000000 291.850000 1115.000000 292.150000 ;
        RECT 1110.000000 295.850000 1115.000000 296.150000 ;
        RECT 1110.000000 299.850000 1115.000000 300.150000 ;
        RECT 1110.000000 303.850000 1115.000000 304.150000 ;
        RECT 1110.000000 311.850000 1115.000000 312.150000 ;
        RECT 1110.000000 307.850000 1115.000000 308.150000 ;
        RECT 1110.000000 323.850000 1115.000000 324.150000 ;
        RECT 1110.000000 319.850000 1115.000000 320.150000 ;
        RECT 1110.000000 315.850000 1115.000000 316.150000 ;
        RECT 1110.000000 339.850000 1115.000000 340.150000 ;
        RECT 1110.000000 335.850000 1115.000000 336.150000 ;
        RECT 1110.000000 331.850000 1115.000000 332.150000 ;
        RECT 1110.000000 327.850000 1115.000000 328.150000 ;
        RECT 1060.000000 283.850000 1065.000000 284.150000 ;
        RECT 1060.000000 279.850000 1065.000000 280.150000 ;
        RECT 1060.000000 275.850000 1065.000000 276.150000 ;
        RECT 1060.000000 271.850000 1065.000000 272.150000 ;
        RECT 1060.000000 287.850000 1065.000000 288.150000 ;
        RECT 1060.000000 291.850000 1065.000000 292.150000 ;
        RECT 1060.000000 295.850000 1065.000000 296.150000 ;
        RECT 1060.000000 299.850000 1065.000000 300.150000 ;
        RECT 1060.000000 303.850000 1065.000000 304.150000 ;
        RECT 1060.000000 307.850000 1065.000000 308.150000 ;
        RECT 1060.000000 311.850000 1065.000000 312.150000 ;
        RECT 1060.000000 315.850000 1065.000000 316.150000 ;
        RECT 1060.000000 319.850000 1065.000000 320.150000 ;
        RECT 1060.000000 323.850000 1065.000000 324.150000 ;
        RECT 1060.000000 339.850000 1065.000000 340.150000 ;
        RECT 1060.000000 335.850000 1065.000000 336.150000 ;
        RECT 1060.000000 331.850000 1065.000000 332.150000 ;
        RECT 1060.000000 327.850000 1065.000000 328.150000 ;
        RECT 1158.000000 283.850000 1168.000000 284.150000 ;
        RECT 1158.000000 279.850000 1168.000000 280.150000 ;
        RECT 1158.000000 275.850000 1168.000000 276.150000 ;
        RECT 1158.000000 271.850000 1168.000000 272.150000 ;
        RECT 1158.000000 287.850000 1168.000000 288.150000 ;
        RECT 1158.000000 291.850000 1168.000000 292.150000 ;
        RECT 1158.000000 295.850000 1168.000000 296.150000 ;
        RECT 1158.000000 299.850000 1168.000000 300.150000 ;
        RECT 1158.000000 303.850000 1168.000000 304.150000 ;
        RECT 1158.000000 307.850000 1168.000000 308.150000 ;
        RECT 1158.000000 311.850000 1168.000000 312.150000 ;
        RECT 1158.000000 315.850000 1168.000000 316.150000 ;
        RECT 1158.000000 319.850000 1168.000000 320.150000 ;
        RECT 1158.000000 323.850000 1168.000000 324.150000 ;
        RECT 1158.000000 339.850000 1168.000000 340.150000 ;
        RECT 1158.000000 335.850000 1168.000000 336.150000 ;
        RECT 1158.000000 331.850000 1168.000000 332.150000 ;
        RECT 1158.000000 327.850000 1168.000000 328.150000 ;
        RECT 60.000000 379.850000 65.000000 380.150000 ;
        RECT 18.000000 379.850000 28.000000 380.150000 ;
        RECT 18.000000 343.850000 28.000000 344.150000 ;
        RECT 18.000000 347.850000 28.000000 348.150000 ;
        RECT 18.000000 351.850000 28.000000 352.150000 ;
        RECT 18.000000 359.850000 28.000000 360.150000 ;
        RECT 18.000000 355.850000 28.000000 356.150000 ;
        RECT 18.000000 375.850000 28.000000 376.150000 ;
        RECT 18.000000 371.850000 28.000000 372.150000 ;
        RECT 18.000000 367.850000 28.000000 368.150000 ;
        RECT 18.000000 363.850000 28.000000 364.150000 ;
        RECT 60.000000 347.850000 65.000000 348.150000 ;
        RECT 60.000000 343.850000 65.000000 344.150000 ;
        RECT 60.000000 352.445000 64.080000 352.745000 ;
        RECT 60.000000 375.850000 65.000000 376.150000 ;
        RECT 60.000000 371.850000 65.000000 372.150000 ;
        RECT 60.000000 367.850000 65.000000 368.150000 ;
        RECT 60.000000 363.850000 65.000000 364.150000 ;
        RECT 18.000000 395.850000 28.000000 396.150000 ;
        RECT 18.000000 391.850000 28.000000 392.150000 ;
        RECT 18.000000 387.850000 28.000000 388.150000 ;
        RECT 18.000000 383.850000 28.000000 384.150000 ;
        RECT 18.000000 407.850000 28.000000 408.150000 ;
        RECT 18.000000 399.850000 28.000000 400.150000 ;
        RECT 18.000000 403.850000 28.000000 404.150000 ;
        RECT 18.000000 411.850000 28.000000 412.150000 ;
        RECT 18.000000 415.850000 28.000000 416.150000 ;
        RECT 60.000000 395.850000 65.000000 396.150000 ;
        RECT 60.000000 391.850000 65.000000 392.150000 ;
        RECT 60.000000 387.850000 65.000000 388.150000 ;
        RECT 60.000000 383.850000 65.000000 384.150000 ;
        RECT 60.000000 407.850000 65.000000 408.150000 ;
        RECT 60.000000 399.850000 65.000000 400.150000 ;
        RECT 60.000000 403.850000 65.000000 404.150000 ;
        RECT 60.000000 411.850000 65.000000 412.150000 ;
        RECT 60.000000 415.850000 65.000000 416.150000 ;
        RECT 110.000000 379.850000 115.000000 380.150000 ;
        RECT 110.000000 351.850000 115.000000 352.150000 ;
        RECT 110.000000 347.850000 115.000000 348.150000 ;
        RECT 110.000000 343.850000 115.000000 344.150000 ;
        RECT 110.000000 359.850000 115.000000 360.150000 ;
        RECT 110.000000 355.850000 115.000000 356.150000 ;
        RECT 110.000000 375.850000 115.000000 376.150000 ;
        RECT 110.000000 371.850000 115.000000 372.150000 ;
        RECT 110.000000 367.850000 115.000000 368.150000 ;
        RECT 110.000000 363.850000 115.000000 364.150000 ;
        RECT 110.000000 383.850000 115.000000 384.150000 ;
        RECT 110.000000 387.850000 115.000000 388.150000 ;
        RECT 110.000000 391.850000 115.000000 392.150000 ;
        RECT 110.000000 395.850000 115.000000 396.150000 ;
        RECT 110.000000 407.850000 115.000000 408.150000 ;
        RECT 110.000000 399.850000 115.000000 400.150000 ;
        RECT 110.000000 403.850000 115.000000 404.150000 ;
        RECT 110.000000 411.850000 115.000000 412.150000 ;
        RECT 110.000000 415.850000 115.000000 416.150000 ;
        RECT 18.000000 431.850000 28.000000 432.150000 ;
        RECT 18.000000 427.850000 28.000000 428.150000 ;
        RECT 18.000000 423.850000 28.000000 424.150000 ;
        RECT 18.000000 419.850000 28.000000 420.150000 ;
        RECT 18.000000 435.850000 28.000000 436.150000 ;
        RECT 18.000000 439.850000 28.000000 440.150000 ;
        RECT 18.000000 443.850000 28.000000 444.150000 ;
        RECT 18.000000 447.850000 28.000000 448.150000 ;
        RECT 18.000000 451.850000 28.000000 452.150000 ;
        RECT 60.000000 431.850000 65.000000 432.150000 ;
        RECT 60.000000 427.850000 65.000000 428.150000 ;
        RECT 60.000000 423.850000 65.000000 424.150000 ;
        RECT 60.000000 419.850000 65.000000 420.150000 ;
        RECT 60.000000 435.850000 65.000000 436.150000 ;
        RECT 60.000000 439.850000 65.000000 440.150000 ;
        RECT 60.000000 443.850000 65.000000 444.150000 ;
        RECT 60.000000 447.850000 65.000000 448.150000 ;
        RECT 60.000000 451.850000 65.000000 452.150000 ;
        RECT 18.000000 455.850000 28.000000 456.150000 ;
        RECT 18.000000 459.850000 28.000000 460.150000 ;
        RECT 18.000000 463.850000 28.000000 464.150000 ;
        RECT 18.000000 467.850000 28.000000 468.150000 ;
        RECT 18.000000 471.850000 28.000000 472.150000 ;
        RECT 18.000000 487.850000 28.000000 488.150000 ;
        RECT 18.000000 483.850000 28.000000 484.150000 ;
        RECT 18.000000 479.850000 28.000000 480.150000 ;
        RECT 18.000000 475.850000 28.000000 476.150000 ;
        RECT 60.000000 455.850000 65.000000 456.150000 ;
        RECT 60.000000 459.850000 65.000000 460.150000 ;
        RECT 60.000000 463.850000 65.000000 464.150000 ;
        RECT 60.000000 467.850000 65.000000 468.150000 ;
        RECT 60.000000 471.850000 65.000000 472.150000 ;
        RECT 60.000000 487.850000 65.000000 488.150000 ;
        RECT 60.000000 483.850000 65.000000 484.150000 ;
        RECT 60.000000 479.850000 65.000000 480.150000 ;
        RECT 60.000000 475.850000 65.000000 476.150000 ;
        RECT 110.000000 419.850000 115.000000 420.150000 ;
        RECT 110.000000 423.850000 115.000000 424.150000 ;
        RECT 110.000000 427.850000 115.000000 428.150000 ;
        RECT 110.000000 431.850000 115.000000 432.150000 ;
        RECT 110.000000 435.850000 115.000000 436.150000 ;
        RECT 110.000000 439.850000 115.000000 440.150000 ;
        RECT 110.000000 443.850000 115.000000 444.150000 ;
        RECT 110.000000 447.850000 115.000000 448.150000 ;
        RECT 110.000000 451.850000 115.000000 452.150000 ;
        RECT 110.000000 459.850000 115.000000 460.150000 ;
        RECT 110.000000 455.850000 115.000000 456.150000 ;
        RECT 110.000000 471.850000 115.000000 472.150000 ;
        RECT 110.000000 467.850000 115.000000 468.150000 ;
        RECT 110.000000 463.850000 115.000000 464.150000 ;
        RECT 110.000000 487.850000 115.000000 488.150000 ;
        RECT 110.000000 483.850000 115.000000 484.150000 ;
        RECT 110.000000 479.850000 115.000000 480.150000 ;
        RECT 110.000000 475.850000 115.000000 476.150000 ;
        RECT 160.000000 379.850000 165.000000 380.150000 ;
        RECT 210.000000 379.850000 215.000000 380.150000 ;
        RECT 160.000000 343.850000 165.000000 344.150000 ;
        RECT 160.000000 347.850000 165.000000 348.150000 ;
        RECT 160.000000 351.850000 165.000000 352.150000 ;
        RECT 160.000000 355.850000 165.000000 356.150000 ;
        RECT 160.000000 359.850000 165.000000 360.150000 ;
        RECT 160.000000 363.850000 165.000000 364.150000 ;
        RECT 160.000000 367.850000 165.000000 368.150000 ;
        RECT 160.000000 375.850000 165.000000 376.150000 ;
        RECT 160.000000 371.850000 165.000000 372.150000 ;
        RECT 210.000000 343.850000 215.000000 344.150000 ;
        RECT 210.000000 347.850000 215.000000 348.150000 ;
        RECT 210.000000 351.850000 215.000000 352.150000 ;
        RECT 210.000000 355.850000 215.000000 356.150000 ;
        RECT 210.000000 359.850000 215.000000 360.150000 ;
        RECT 210.000000 363.850000 215.000000 364.150000 ;
        RECT 210.000000 367.850000 215.000000 368.150000 ;
        RECT 210.000000 371.850000 215.000000 372.150000 ;
        RECT 210.000000 375.850000 215.000000 376.150000 ;
        RECT 160.000000 387.850000 165.000000 388.150000 ;
        RECT 160.000000 383.850000 165.000000 384.150000 ;
        RECT 160.000000 391.850000 165.000000 392.150000 ;
        RECT 160.000000 395.850000 165.000000 396.150000 ;
        RECT 160.000000 399.850000 165.000000 400.150000 ;
        RECT 210.000000 383.850000 215.000000 384.150000 ;
        RECT 210.000000 387.850000 215.000000 388.150000 ;
        RECT 210.000000 391.850000 215.000000 392.150000 ;
        RECT 210.000000 395.850000 215.000000 396.150000 ;
        RECT 210.000000 407.850000 215.000000 408.150000 ;
        RECT 210.000000 399.850000 215.000000 400.150000 ;
        RECT 210.000000 403.850000 215.000000 404.150000 ;
        RECT 210.000000 411.850000 215.000000 412.150000 ;
        RECT 210.000000 415.850000 215.000000 416.150000 ;
        RECT 260.000000 379.850000 265.000000 380.150000 ;
        RECT 260.000000 343.850000 265.000000 344.150000 ;
        RECT 260.000000 347.850000 265.000000 348.150000 ;
        RECT 260.000000 351.850000 265.000000 352.150000 ;
        RECT 260.000000 355.850000 265.000000 356.150000 ;
        RECT 260.000000 359.850000 265.000000 360.150000 ;
        RECT 260.000000 367.850000 265.000000 368.150000 ;
        RECT 260.000000 363.850000 265.000000 364.150000 ;
        RECT 260.000000 375.850000 265.000000 376.150000 ;
        RECT 260.000000 371.850000 265.000000 372.150000 ;
        RECT 260.000000 383.850000 265.000000 384.150000 ;
        RECT 260.000000 387.850000 265.000000 388.150000 ;
        RECT 260.000000 391.850000 265.000000 392.150000 ;
        RECT 260.000000 395.850000 265.000000 396.150000 ;
        RECT 260.000000 399.850000 265.000000 400.150000 ;
        RECT 210.000000 431.850000 215.000000 432.150000 ;
        RECT 210.000000 427.850000 215.000000 428.150000 ;
        RECT 210.000000 423.850000 215.000000 424.150000 ;
        RECT 210.000000 419.850000 215.000000 420.150000 ;
        RECT 210.000000 435.850000 215.000000 436.150000 ;
        RECT 210.000000 439.850000 215.000000 440.150000 ;
        RECT 210.000000 443.850000 215.000000 444.150000 ;
        RECT 210.000000 447.850000 215.000000 448.150000 ;
        RECT 210.000000 451.850000 215.000000 452.150000 ;
        RECT 160.000000 463.850000 165.000000 464.150000 ;
        RECT 160.000000 467.850000 165.000000 468.150000 ;
        RECT 160.000000 471.850000 165.000000 472.150000 ;
        RECT 160.000000 479.850000 165.000000 480.150000 ;
        RECT 160.000000 475.850000 165.000000 476.150000 ;
        RECT 160.000000 487.850000 165.000000 488.150000 ;
        RECT 160.000000 483.850000 165.000000 484.150000 ;
        RECT 210.000000 455.850000 215.000000 456.150000 ;
        RECT 210.000000 459.850000 215.000000 460.150000 ;
        RECT 210.000000 463.850000 215.000000 464.150000 ;
        RECT 210.000000 467.850000 215.000000 468.150000 ;
        RECT 210.000000 471.850000 215.000000 472.150000 ;
        RECT 210.000000 475.850000 215.000000 476.150000 ;
        RECT 210.000000 479.850000 215.000000 480.150000 ;
        RECT 210.000000 483.850000 215.000000 484.150000 ;
        RECT 210.000000 487.850000 215.000000 488.150000 ;
        RECT 260.000000 467.850000 265.000000 468.150000 ;
        RECT 260.000000 463.850000 265.000000 464.150000 ;
        RECT 260.000000 471.850000 265.000000 472.150000 ;
        RECT 260.000000 475.850000 265.000000 476.150000 ;
        RECT 260.000000 479.850000 265.000000 480.150000 ;
        RECT 260.000000 483.850000 265.000000 484.150000 ;
        RECT 260.000000 487.850000 265.000000 488.150000 ;
        RECT 18.000000 491.850000 28.000000 492.150000 ;
        RECT 18.000000 495.850000 28.000000 496.150000 ;
        RECT 18.000000 499.850000 28.000000 500.150000 ;
        RECT 18.000000 503.850000 28.000000 504.150000 ;
        RECT 18.000000 507.850000 28.000000 508.150000 ;
        RECT 18.000000 515.850000 28.000000 516.150000 ;
        RECT 18.000000 511.850000 28.000000 512.150000 ;
        RECT 60.000000 491.850000 65.000000 492.150000 ;
        RECT 60.000000 495.850000 65.000000 496.150000 ;
        RECT 60.000000 499.850000 65.000000 500.150000 ;
        RECT 60.000000 503.850000 65.000000 504.150000 ;
        RECT 60.000000 507.850000 65.000000 508.150000 ;
        RECT 60.000000 515.850000 65.000000 516.150000 ;
        RECT 60.000000 511.850000 65.000000 512.150000 ;
        RECT 110.000000 499.850000 115.000000 500.150000 ;
        RECT 110.000000 495.850000 115.000000 496.150000 ;
        RECT 110.000000 491.850000 115.000000 492.150000 ;
        RECT 110.000000 507.850000 115.000000 508.150000 ;
        RECT 110.000000 503.850000 115.000000 504.150000 ;
        RECT 110.000000 515.850000 115.000000 516.150000 ;
        RECT 110.000000 511.850000 115.000000 512.150000 ;
        RECT 160.000000 491.850000 165.000000 492.150000 ;
        RECT 160.000000 495.850000 165.000000 496.150000 ;
        RECT 160.000000 499.850000 165.000000 500.150000 ;
        RECT 160.000000 507.850000 165.000000 508.150000 ;
        RECT 160.000000 503.850000 165.000000 504.150000 ;
        RECT 160.000000 515.850000 165.000000 516.150000 ;
        RECT 160.000000 511.850000 165.000000 512.150000 ;
        RECT 210.000000 491.850000 215.000000 492.150000 ;
        RECT 210.000000 495.850000 215.000000 496.150000 ;
        RECT 210.000000 499.850000 215.000000 500.150000 ;
        RECT 210.000000 503.850000 215.000000 504.150000 ;
        RECT 210.000000 507.850000 215.000000 508.150000 ;
        RECT 210.000000 515.850000 215.000000 516.150000 ;
        RECT 210.000000 511.850000 215.000000 512.150000 ;
        RECT 260.000000 495.850000 265.000000 496.150000 ;
        RECT 260.000000 491.850000 265.000000 492.150000 ;
        RECT 260.000000 499.850000 265.000000 500.150000 ;
        RECT 260.000000 503.850000 265.000000 504.150000 ;
        RECT 260.000000 507.850000 265.000000 508.150000 ;
        RECT 260.000000 515.850000 265.000000 516.150000 ;
        RECT 260.000000 511.850000 265.000000 512.150000 ;
        RECT 360.000000 379.850000 365.000000 380.150000 ;
        RECT 310.000000 379.850000 315.000000 380.150000 ;
        RECT 310.000000 343.850000 315.000000 344.150000 ;
        RECT 310.000000 351.850000 315.000000 352.150000 ;
        RECT 310.000000 347.850000 315.000000 348.150000 ;
        RECT 310.000000 355.850000 315.000000 356.150000 ;
        RECT 310.000000 359.850000 315.000000 360.150000 ;
        RECT 310.000000 363.850000 315.000000 364.150000 ;
        RECT 310.000000 367.850000 315.000000 368.150000 ;
        RECT 310.000000 371.850000 315.000000 372.150000 ;
        RECT 310.000000 375.850000 315.000000 376.150000 ;
        RECT 360.000000 343.850000 365.000000 344.150000 ;
        RECT 360.000000 347.850000 365.000000 348.150000 ;
        RECT 360.000000 351.850000 365.000000 352.150000 ;
        RECT 360.000000 355.850000 365.000000 356.150000 ;
        RECT 360.000000 359.850000 365.000000 360.150000 ;
        RECT 360.000000 363.850000 365.000000 364.150000 ;
        RECT 360.000000 367.850000 365.000000 368.150000 ;
        RECT 360.000000 371.850000 365.000000 372.150000 ;
        RECT 360.000000 375.850000 365.000000 376.150000 ;
        RECT 310.000000 383.850000 315.000000 384.150000 ;
        RECT 310.000000 387.850000 315.000000 388.150000 ;
        RECT 310.000000 391.850000 315.000000 392.150000 ;
        RECT 310.000000 395.850000 315.000000 396.150000 ;
        RECT 310.000000 407.850000 315.000000 408.150000 ;
        RECT 310.000000 399.850000 315.000000 400.150000 ;
        RECT 310.000000 403.850000 315.000000 404.150000 ;
        RECT 310.000000 411.850000 315.000000 412.150000 ;
        RECT 310.000000 415.850000 315.000000 416.150000 ;
        RECT 360.000000 383.850000 365.000000 384.150000 ;
        RECT 360.000000 387.850000 365.000000 388.150000 ;
        RECT 360.000000 391.850000 365.000000 392.150000 ;
        RECT 360.000000 395.850000 365.000000 396.150000 ;
        RECT 360.000000 407.850000 365.000000 408.150000 ;
        RECT 360.000000 399.850000 365.000000 400.150000 ;
        RECT 360.000000 403.850000 365.000000 404.150000 ;
        RECT 360.000000 411.850000 365.000000 412.150000 ;
        RECT 360.000000 415.850000 365.000000 416.150000 ;
        RECT 410.000000 379.850000 415.000000 380.150000 ;
        RECT 410.000000 359.850000 415.000000 360.150000 ;
        RECT 410.000000 355.850000 415.000000 356.150000 ;
        RECT 410.000000 351.850000 415.000000 352.150000 ;
        RECT 410.000000 347.850000 415.000000 348.150000 ;
        RECT 410.000000 343.850000 415.000000 344.150000 ;
        RECT 410.000000 367.850000 415.000000 368.150000 ;
        RECT 410.000000 363.850000 415.000000 364.150000 ;
        RECT 410.000000 371.850000 415.000000 372.150000 ;
        RECT 410.000000 375.850000 415.000000 376.150000 ;
        RECT 410.000000 383.850000 415.000000 384.150000 ;
        RECT 410.000000 387.850000 415.000000 388.150000 ;
        RECT 410.000000 391.850000 415.000000 392.150000 ;
        RECT 410.000000 395.850000 415.000000 396.150000 ;
        RECT 410.000000 407.850000 415.000000 408.150000 ;
        RECT 410.000000 399.850000 415.000000 400.150000 ;
        RECT 410.000000 403.850000 415.000000 404.150000 ;
        RECT 410.000000 411.850000 415.000000 412.150000 ;
        RECT 410.000000 415.850000 415.000000 416.150000 ;
        RECT 361.000000 479.850000 371.000000 480.150000 ;
        RECT 361.000000 483.850000 371.000000 484.150000 ;
        RECT 361.000000 487.850000 371.000000 488.150000 ;
        RECT 310.000000 419.850000 315.000000 420.150000 ;
        RECT 310.000000 423.850000 315.000000 424.150000 ;
        RECT 310.000000 427.850000 315.000000 428.150000 ;
        RECT 310.000000 431.850000 315.000000 432.150000 ;
        RECT 310.000000 439.850000 315.000000 440.150000 ;
        RECT 310.000000 435.850000 315.000000 436.150000 ;
        RECT 310.000000 443.850000 315.000000 444.150000 ;
        RECT 310.000000 447.850000 315.000000 448.150000 ;
        RECT 310.000000 451.850000 315.000000 452.150000 ;
        RECT 360.000000 419.850000 365.000000 420.150000 ;
        RECT 360.000000 423.850000 365.000000 424.150000 ;
        RECT 360.000000 427.850000 365.000000 428.150000 ;
        RECT 360.000000 431.850000 365.000000 432.150000 ;
        RECT 360.000000 435.850000 365.000000 436.150000 ;
        RECT 360.000000 439.850000 365.000000 440.150000 ;
        RECT 360.000000 443.850000 365.000000 444.150000 ;
        RECT 360.000000 447.850000 365.000000 448.150000 ;
        RECT 360.000000 451.850000 365.000000 452.150000 ;
        RECT 310.000000 455.850000 315.000000 456.150000 ;
        RECT 310.000000 459.850000 315.000000 460.150000 ;
        RECT 310.000000 467.850000 315.000000 468.150000 ;
        RECT 310.000000 463.850000 315.000000 464.150000 ;
        RECT 310.000000 471.850000 315.000000 472.150000 ;
        RECT 310.000000 475.850000 315.000000 476.150000 ;
        RECT 310.000000 479.850000 315.000000 480.150000 ;
        RECT 310.000000 483.850000 315.000000 484.150000 ;
        RECT 310.000000 487.850000 315.000000 488.150000 ;
        RECT 360.000000 455.850000 365.000000 456.150000 ;
        RECT 360.000000 459.850000 365.000000 460.150000 ;
        RECT 360.000000 471.850000 368.500000 472.150000 ;
        RECT 360.000000 463.850000 365.000000 464.150000 ;
        RECT 360.000000 467.850000 365.000000 468.150000 ;
        RECT 363.500000 475.850000 368.500000 476.150000 ;
        RECT 410.000000 419.850000 415.000000 420.150000 ;
        RECT 410.000000 423.850000 415.000000 424.150000 ;
        RECT 410.000000 431.850000 415.000000 432.150000 ;
        RECT 410.000000 427.850000 415.000000 428.150000 ;
        RECT 410.000000 435.850000 415.000000 436.150000 ;
        RECT 410.000000 439.850000 415.000000 440.150000 ;
        RECT 410.000000 443.850000 415.000000 444.150000 ;
        RECT 410.000000 447.850000 415.000000 448.150000 ;
        RECT 410.000000 451.850000 415.000000 452.150000 ;
        RECT 410.000000 459.850000 415.000000 460.150000 ;
        RECT 410.000000 455.850000 415.000000 456.150000 ;
        RECT 410.000000 471.850000 415.000000 472.150000 ;
        RECT 410.000000 467.850000 415.000000 468.150000 ;
        RECT 410.000000 463.850000 415.000000 464.150000 ;
        RECT 410.000000 479.850000 415.000000 480.150000 ;
        RECT 410.000000 475.850000 415.000000 476.150000 ;
        RECT 410.000000 487.850000 415.000000 488.150000 ;
        RECT 410.000000 483.850000 415.000000 484.150000 ;
        RECT 460.000000 379.850000 465.000000 380.150000 ;
        RECT 510.000000 379.850000 515.000000 380.150000 ;
        RECT 460.000000 347.850000 465.000000 348.150000 ;
        RECT 460.000000 343.850000 465.000000 344.150000 ;
        RECT 460.000000 351.230000 465.000000 352.230000 ;
        RECT 460.000000 375.850000 465.000000 376.150000 ;
        RECT 460.000000 371.850000 465.000000 372.150000 ;
        RECT 510.000000 343.850000 515.000000 344.150000 ;
        RECT 510.000000 347.850000 515.000000 348.150000 ;
        RECT 510.000000 351.850000 515.000000 352.150000 ;
        RECT 510.000000 359.850000 515.000000 360.150000 ;
        RECT 510.000000 355.850000 515.000000 356.150000 ;
        RECT 510.000000 363.850000 515.000000 364.150000 ;
        RECT 510.000000 367.850000 515.000000 368.150000 ;
        RECT 510.000000 375.850000 515.000000 376.150000 ;
        RECT 510.000000 371.850000 515.000000 372.150000 ;
        RECT 460.000000 383.850000 465.000000 384.150000 ;
        RECT 460.000000 387.850000 465.000000 388.150000 ;
        RECT 460.000000 391.850000 465.000000 392.150000 ;
        RECT 460.000000 395.850000 465.000000 396.150000 ;
        RECT 460.000000 401.230000 465.000000 402.230000 ;
        RECT 510.000000 387.850000 515.000000 388.150000 ;
        RECT 510.000000 383.850000 515.000000 384.150000 ;
        RECT 510.000000 391.850000 515.000000 392.150000 ;
        RECT 510.000000 395.850000 515.000000 396.150000 ;
        RECT 510.000000 407.850000 515.000000 408.150000 ;
        RECT 510.000000 399.850000 515.000000 400.150000 ;
        RECT 510.000000 403.850000 515.000000 404.150000 ;
        RECT 510.000000 411.850000 515.000000 412.150000 ;
        RECT 510.000000 415.850000 515.000000 416.150000 ;
        RECT 560.000000 379.850000 565.000000 380.150000 ;
        RECT 560.000000 359.850000 565.000000 360.150000 ;
        RECT 560.000000 355.850000 565.000000 356.150000 ;
        RECT 560.000000 351.850000 565.000000 352.150000 ;
        RECT 560.000000 347.850000 565.000000 348.150000 ;
        RECT 560.000000 343.850000 565.000000 344.150000 ;
        RECT 560.000000 375.850000 565.000000 376.150000 ;
        RECT 560.000000 371.850000 565.000000 372.150000 ;
        RECT 560.000000 367.850000 565.000000 368.150000 ;
        RECT 560.000000 363.850000 565.000000 364.150000 ;
        RECT 560.000000 383.850000 565.000000 384.150000 ;
        RECT 560.000000 387.850000 565.000000 388.150000 ;
        RECT 560.000000 395.850000 565.000000 396.150000 ;
        RECT 560.000000 391.850000 565.000000 392.150000 ;
        RECT 560.000000 407.850000 565.000000 408.150000 ;
        RECT 560.000000 403.850000 565.000000 404.150000 ;
        RECT 560.000000 399.850000 565.000000 400.150000 ;
        RECT 560.000000 415.850000 565.000000 416.150000 ;
        RECT 560.000000 411.850000 565.000000 412.150000 ;
        RECT 460.000000 419.850000 465.000000 420.150000 ;
        RECT 460.000000 431.850000 465.000000 432.150000 ;
        RECT 460.000000 427.850000 465.000000 428.150000 ;
        RECT 460.000000 423.850000 465.000000 424.150000 ;
        RECT 460.000000 435.850000 465.000000 436.150000 ;
        RECT 460.000000 439.850000 465.000000 440.150000 ;
        RECT 460.000000 443.850000 465.000000 444.150000 ;
        RECT 460.000000 447.850000 465.000000 448.150000 ;
        RECT 460.000000 451.850000 465.000000 452.150000 ;
        RECT 510.000000 419.850000 515.000000 420.150000 ;
        RECT 510.000000 423.850000 515.000000 424.150000 ;
        RECT 510.000000 431.850000 515.000000 432.150000 ;
        RECT 510.000000 427.850000 515.000000 428.150000 ;
        RECT 510.000000 439.850000 515.000000 440.150000 ;
        RECT 510.000000 435.850000 515.000000 436.150000 ;
        RECT 510.000000 443.850000 515.000000 444.150000 ;
        RECT 510.000000 447.850000 515.000000 448.150000 ;
        RECT 510.000000 451.850000 515.000000 452.150000 ;
        RECT 460.000000 455.850000 465.000000 456.150000 ;
        RECT 460.000000 459.850000 465.000000 460.150000 ;
        RECT 460.000000 463.850000 465.000000 464.150000 ;
        RECT 460.000000 467.850000 465.000000 468.150000 ;
        RECT 460.000000 471.850000 465.000000 472.150000 ;
        RECT 460.000000 487.850000 465.000000 488.150000 ;
        RECT 460.000000 483.850000 465.000000 484.150000 ;
        RECT 460.000000 479.850000 465.000000 480.150000 ;
        RECT 460.000000 475.850000 465.000000 476.150000 ;
        RECT 510.000000 455.850000 515.000000 456.150000 ;
        RECT 510.000000 459.850000 515.000000 460.150000 ;
        RECT 510.000000 467.850000 515.000000 468.150000 ;
        RECT 510.000000 463.850000 515.000000 464.150000 ;
        RECT 510.000000 471.850000 515.000000 472.150000 ;
        RECT 510.000000 475.850000 515.000000 476.150000 ;
        RECT 510.000000 479.850000 515.000000 480.150000 ;
        RECT 510.000000 483.850000 515.000000 484.150000 ;
        RECT 510.000000 487.850000 515.000000 488.150000 ;
        RECT 560.000000 419.850000 565.000000 420.150000 ;
        RECT 560.000000 423.850000 565.000000 424.150000 ;
        RECT 560.000000 427.850000 565.000000 428.150000 ;
        RECT 560.000000 431.850000 565.000000 432.150000 ;
        RECT 560.000000 435.850000 565.000000 436.150000 ;
        RECT 560.000000 439.850000 565.000000 440.150000 ;
        RECT 560.000000 443.850000 565.000000 444.150000 ;
        RECT 560.000000 451.850000 565.000000 452.150000 ;
        RECT 560.000000 447.850000 565.000000 448.150000 ;
        RECT 560.000000 455.850000 565.000000 456.150000 ;
        RECT 560.000000 459.850000 565.000000 460.150000 ;
        RECT 560.000000 463.850000 565.000000 464.150000 ;
        RECT 560.000000 467.850000 565.000000 468.150000 ;
        RECT 560.000000 471.850000 565.000000 472.150000 ;
        RECT 560.000000 487.850000 565.000000 488.150000 ;
        RECT 560.000000 483.850000 565.000000 484.150000 ;
        RECT 560.000000 479.850000 565.000000 480.150000 ;
        RECT 560.000000 475.850000 565.000000 476.150000 ;
        RECT 360.000000 499.850000 371.000000 500.150000 ;
        RECT 360.000000 491.850000 371.000000 492.150000 ;
        RECT 360.000000 495.850000 371.000000 496.150000 ;
        RECT 360.000000 507.850000 371.000000 508.150000 ;
        RECT 360.000000 503.850000 371.000000 504.150000 ;
        RECT 360.000000 511.850000 371.000000 512.150000 ;
        RECT 360.000000 515.850000 371.000000 516.150000 ;
        RECT 360.000000 527.850000 371.000000 528.150000 ;
        RECT 360.000000 523.850000 371.000000 524.150000 ;
        RECT 360.000000 519.850000 371.000000 520.150000 ;
        RECT 360.000000 535.850000 371.000000 536.150000 ;
        RECT 360.000000 531.850000 371.000000 532.150000 ;
        RECT 360.000000 543.850000 371.000000 544.150000 ;
        RECT 360.000000 539.850000 371.000000 540.150000 ;
        RECT 360.000000 555.850000 371.000000 556.150000 ;
        RECT 360.000000 547.850000 371.000000 548.150000 ;
        RECT 360.000000 551.850000 371.000000 552.150000 ;
        RECT 360.000000 563.850000 371.000000 564.150000 ;
        RECT 360.000000 559.850000 371.000000 560.150000 ;
        RECT 310.000000 495.850000 315.000000 496.150000 ;
        RECT 310.000000 491.850000 315.000000 492.150000 ;
        RECT 310.000000 499.850000 315.000000 500.150000 ;
        RECT 310.000000 507.850000 315.000000 508.150000 ;
        RECT 310.000000 503.850000 315.000000 504.150000 ;
        RECT 310.000000 515.850000 315.000000 516.150000 ;
        RECT 310.000000 511.850000 315.000000 512.150000 ;
        RECT 410.000000 491.850000 415.000000 492.150000 ;
        RECT 410.000000 495.850000 415.000000 496.150000 ;
        RECT 410.000000 499.850000 415.000000 500.150000 ;
        RECT 410.000000 503.850000 415.000000 504.150000 ;
        RECT 360.000000 583.850000 371.000000 584.150000 ;
        RECT 360.000000 571.850000 371.000000 572.150000 ;
        RECT 360.000000 567.850000 371.000000 568.150000 ;
        RECT 360.000000 579.850000 371.000000 580.150000 ;
        RECT 360.000000 575.850000 371.000000 576.150000 ;
        RECT 360.000000 587.850000 371.000000 588.150000 ;
        RECT 360.000000 591.850000 371.000000 592.150000 ;
        RECT 360.000000 599.850000 371.000000 600.150000 ;
        RECT 360.000000 595.850000 371.000000 596.150000 ;
        RECT 360.000000 607.850000 371.000000 608.150000 ;
        RECT 360.000000 603.850000 371.000000 604.150000 ;
        RECT 360.000000 619.850000 371.000000 620.150000 ;
        RECT 360.000000 615.850000 371.000000 616.150000 ;
        RECT 360.000000 611.850000 371.000000 612.150000 ;
        RECT 360.000000 623.850000 371.000000 624.150000 ;
        RECT 360.000000 627.850000 371.000000 628.150000 ;
        RECT 360.000000 635.850000 371.000000 636.150000 ;
        RECT 360.000000 631.850000 371.000000 632.150000 ;
        RECT 460.000000 503.850000 465.000000 504.150000 ;
        RECT 460.000000 499.850000 465.000000 500.150000 ;
        RECT 460.000000 491.850000 465.000000 492.150000 ;
        RECT 460.000000 495.850000 465.000000 496.150000 ;
        RECT 510.000000 495.850000 515.000000 496.150000 ;
        RECT 510.000000 491.850000 515.000000 492.150000 ;
        RECT 510.000000 499.850000 515.000000 500.150000 ;
        RECT 510.000000 503.850000 515.000000 504.150000 ;
        RECT 560.000000 503.850000 565.000000 504.150000 ;
        RECT 560.000000 499.850000 565.000000 500.150000 ;
        RECT 560.000000 495.850000 565.000000 496.150000 ;
        RECT 560.000000 491.850000 565.000000 492.150000 ;
        RECT 360.000000 639.850000 371.000000 640.150000 ;
        RECT 360.000000 643.850000 371.000000 644.150000 ;
        RECT 360.000000 647.850000 371.000000 648.150000 ;
        RECT 360.000000 655.850000 371.000000 656.150000 ;
        RECT 360.000000 651.850000 371.000000 652.150000 ;
        RECT 360.000000 667.850000 371.000000 668.150000 ;
        RECT 360.000000 663.850000 371.000000 664.150000 ;
        RECT 360.000000 659.850000 371.000000 660.150000 ;
        RECT 360.000000 675.850000 365.000000 676.150000 ;
        RECT 360.000000 671.850000 365.000000 672.150000 ;
        RECT 310.000000 679.850000 315.000000 680.150000 ;
        RECT 310.000000 683.850000 315.000000 684.150000 ;
        RECT 360.000000 679.850000 365.000000 680.150000 ;
        RECT 360.000000 683.850000 365.000000 684.150000 ;
        RECT 410.000000 659.850000 415.000000 660.150000 ;
        RECT 410.000000 663.850000 415.000000 664.150000 ;
        RECT 410.000000 667.850000 415.000000 668.150000 ;
        RECT 410.000000 671.850000 415.000000 672.150000 ;
        RECT 410.000000 675.850000 415.000000 676.150000 ;
        RECT 410.000000 683.850000 415.000000 684.150000 ;
        RECT 410.000000 679.850000 415.000000 680.150000 ;
        RECT 460.000000 659.850000 465.000000 660.150000 ;
        RECT 460.000000 663.850000 465.000000 664.150000 ;
        RECT 460.000000 667.850000 465.000000 668.150000 ;
        RECT 460.000000 671.850000 465.000000 672.150000 ;
        RECT 460.000000 675.850000 465.000000 676.150000 ;
        RECT 510.000000 659.850000 515.000000 660.150000 ;
        RECT 510.000000 663.850000 515.000000 664.150000 ;
        RECT 510.000000 667.850000 515.000000 668.150000 ;
        RECT 510.000000 671.850000 515.000000 672.150000 ;
        RECT 510.000000 675.850000 515.000000 676.150000 ;
        RECT 460.000000 683.850000 465.000000 684.150000 ;
        RECT 460.000000 679.850000 465.000000 680.150000 ;
        RECT 510.000000 683.850000 515.000000 684.150000 ;
        RECT 510.000000 679.850000 515.000000 680.150000 ;
        RECT 560.000000 659.850000 565.000000 660.150000 ;
        RECT 560.000000 663.850000 565.000000 664.150000 ;
        RECT 560.000000 667.850000 565.000000 668.150000 ;
        RECT 560.000000 671.850000 565.000000 672.150000 ;
        RECT 560.000000 675.850000 565.000000 676.150000 ;
        RECT 560.000000 683.850000 565.000000 684.150000 ;
        RECT 560.000000 679.850000 565.000000 680.150000 ;
        RECT 610.000000 379.850000 615.000000 380.150000 ;
        RECT 660.000000 379.850000 665.000000 380.150000 ;
        RECT 610.000000 343.850000 615.000000 344.150000 ;
        RECT 610.000000 347.850000 615.000000 348.150000 ;
        RECT 610.000000 351.850000 615.000000 352.150000 ;
        RECT 610.000000 355.850000 615.000000 356.150000 ;
        RECT 610.000000 359.850000 615.000000 360.150000 ;
        RECT 610.000000 375.850000 615.000000 376.150000 ;
        RECT 610.000000 371.850000 615.000000 372.150000 ;
        RECT 610.000000 367.850000 615.000000 368.150000 ;
        RECT 610.000000 363.850000 615.000000 364.150000 ;
        RECT 660.000000 343.850000 665.000000 344.150000 ;
        RECT 660.000000 347.850000 665.000000 348.150000 ;
        RECT 660.000000 351.850000 665.000000 352.150000 ;
        RECT 660.000000 359.850000 665.000000 360.150000 ;
        RECT 660.000000 355.850000 665.000000 356.150000 ;
        RECT 660.000000 363.850000 665.000000 364.150000 ;
        RECT 660.000000 367.850000 665.000000 368.150000 ;
        RECT 660.000000 375.850000 665.000000 376.150000 ;
        RECT 660.000000 371.850000 665.000000 372.150000 ;
        RECT 610.000000 395.850000 615.000000 396.150000 ;
        RECT 610.000000 391.850000 615.000000 392.150000 ;
        RECT 610.000000 387.850000 615.000000 388.150000 ;
        RECT 610.000000 383.850000 615.000000 384.150000 ;
        RECT 610.000000 407.850000 615.000000 408.150000 ;
        RECT 610.000000 399.850000 615.000000 400.150000 ;
        RECT 610.000000 403.850000 615.000000 404.150000 ;
        RECT 610.000000 411.850000 615.000000 412.150000 ;
        RECT 610.000000 415.850000 615.000000 416.150000 ;
        RECT 660.000000 387.850000 665.000000 388.150000 ;
        RECT 660.000000 383.850000 665.000000 384.150000 ;
        RECT 660.000000 391.850000 665.000000 392.150000 ;
        RECT 660.000000 395.850000 665.000000 396.150000 ;
        RECT 660.000000 407.850000 665.000000 408.150000 ;
        RECT 660.000000 403.850000 665.000000 404.150000 ;
        RECT 660.000000 399.850000 665.000000 400.150000 ;
        RECT 660.000000 411.850000 665.000000 412.150000 ;
        RECT 660.000000 415.850000 665.000000 416.150000 ;
        RECT 710.000000 379.850000 715.000000 380.150000 ;
        RECT 710.000000 359.850000 715.000000 360.150000 ;
        RECT 710.000000 355.850000 715.000000 356.150000 ;
        RECT 710.000000 351.850000 715.000000 352.150000 ;
        RECT 710.000000 347.850000 715.000000 348.150000 ;
        RECT 710.000000 343.850000 715.000000 344.150000 ;
        RECT 710.000000 375.850000 715.000000 376.150000 ;
        RECT 710.000000 371.850000 715.000000 372.150000 ;
        RECT 710.000000 367.850000 715.000000 368.150000 ;
        RECT 710.000000 363.850000 715.000000 364.150000 ;
        RECT 710.000000 395.850000 715.000000 396.150000 ;
        RECT 710.000000 391.850000 715.000000 392.150000 ;
        RECT 710.000000 387.850000 715.000000 388.150000 ;
        RECT 710.000000 383.850000 715.000000 384.150000 ;
        RECT 710.000000 407.850000 715.000000 408.150000 ;
        RECT 710.000000 403.850000 715.000000 404.150000 ;
        RECT 710.000000 399.850000 715.000000 400.150000 ;
        RECT 710.000000 411.850000 718.500000 412.150000 ;
        RECT 713.500000 415.850000 718.500000 416.150000 ;
        RECT 610.000000 431.850000 615.000000 432.150000 ;
        RECT 610.000000 427.850000 615.000000 428.150000 ;
        RECT 610.000000 423.850000 615.000000 424.150000 ;
        RECT 610.000000 419.850000 615.000000 420.150000 ;
        RECT 610.000000 435.850000 615.000000 436.150000 ;
        RECT 610.000000 439.850000 615.000000 440.150000 ;
        RECT 610.000000 443.850000 615.000000 444.150000 ;
        RECT 610.000000 447.850000 615.000000 448.150000 ;
        RECT 610.000000 451.850000 615.000000 452.150000 ;
        RECT 660.000000 419.850000 665.000000 420.150000 ;
        RECT 660.000000 423.850000 665.000000 424.150000 ;
        RECT 660.000000 431.850000 665.000000 432.150000 ;
        RECT 660.000000 427.850000 665.000000 428.150000 ;
        RECT 660.000000 439.850000 665.000000 440.150000 ;
        RECT 660.000000 435.850000 665.000000 436.150000 ;
        RECT 660.000000 443.850000 665.000000 444.150000 ;
        RECT 660.000000 447.850000 665.000000 448.150000 ;
        RECT 660.000000 451.850000 665.000000 452.150000 ;
        RECT 610.000000 455.850000 615.000000 456.150000 ;
        RECT 610.000000 459.850000 615.000000 460.150000 ;
        RECT 610.000000 463.850000 615.000000 464.150000 ;
        RECT 610.000000 467.850000 615.000000 468.150000 ;
        RECT 610.000000 471.850000 615.000000 472.150000 ;
        RECT 610.000000 487.850000 615.000000 488.150000 ;
        RECT 610.000000 483.850000 615.000000 484.150000 ;
        RECT 610.000000 479.850000 615.000000 480.150000 ;
        RECT 610.000000 475.850000 615.000000 476.150000 ;
        RECT 660.000000 459.850000 665.000000 460.150000 ;
        RECT 660.000000 455.850000 665.000000 456.150000 ;
        RECT 660.000000 463.850000 665.000000 464.150000 ;
        RECT 660.000000 467.850000 665.000000 468.150000 ;
        RECT 660.000000 471.850000 665.000000 472.150000 ;
        RECT 660.000000 479.850000 665.000000 480.150000 ;
        RECT 660.000000 475.850000 665.000000 476.150000 ;
        RECT 660.000000 487.850000 665.000000 488.150000 ;
        RECT 660.000000 483.850000 665.000000 484.150000 ;
        RECT 711.000000 423.850000 721.000000 424.150000 ;
        RECT 711.000000 419.850000 721.000000 420.150000 ;
        RECT 710.000000 431.850000 721.000000 432.150000 ;
        RECT 711.000000 427.850000 721.000000 428.150000 ;
        RECT 710.000000 435.850000 721.000000 436.150000 ;
        RECT 710.000000 439.850000 721.000000 440.150000 ;
        RECT 710.000000 443.850000 721.000000 444.150000 ;
        RECT 710.000000 451.850000 721.000000 452.150000 ;
        RECT 710.000000 447.850000 721.000000 448.150000 ;
        RECT 710.000000 455.850000 721.000000 456.150000 ;
        RECT 710.000000 459.850000 721.000000 460.150000 ;
        RECT 710.000000 471.850000 721.000000 472.150000 ;
        RECT 710.000000 463.850000 721.000000 464.150000 ;
        RECT 710.000000 467.850000 721.000000 468.150000 ;
        RECT 710.000000 475.850000 721.000000 476.150000 ;
        RECT 710.000000 479.850000 721.000000 480.150000 ;
        RECT 710.000000 483.850000 721.000000 484.150000 ;
        RECT 710.000000 487.850000 721.000000 488.150000 ;
        RECT 810.000000 379.850000 815.000000 380.150000 ;
        RECT 760.000000 379.850000 765.000000 380.150000 ;
        RECT 760.000000 343.850000 765.000000 344.150000 ;
        RECT 760.000000 347.850000 765.000000 348.150000 ;
        RECT 760.000000 351.850000 765.000000 352.150000 ;
        RECT 760.000000 355.850000 765.000000 356.150000 ;
        RECT 760.000000 359.850000 765.000000 360.150000 ;
        RECT 760.000000 375.850000 765.000000 376.150000 ;
        RECT 760.000000 371.850000 765.000000 372.150000 ;
        RECT 760.000000 367.850000 765.000000 368.150000 ;
        RECT 760.000000 363.850000 765.000000 364.150000 ;
        RECT 810.000000 343.850000 815.000000 344.150000 ;
        RECT 810.000000 347.850000 815.000000 348.150000 ;
        RECT 810.000000 351.850000 815.000000 352.150000 ;
        RECT 810.000000 359.850000 815.000000 360.150000 ;
        RECT 810.000000 355.850000 815.000000 356.150000 ;
        RECT 810.000000 363.850000 815.000000 364.150000 ;
        RECT 810.000000 367.850000 815.000000 368.150000 ;
        RECT 810.000000 375.850000 815.000000 376.150000 ;
        RECT 810.000000 371.850000 815.000000 372.150000 ;
        RECT 760.000000 395.850000 765.000000 396.150000 ;
        RECT 760.000000 391.850000 765.000000 392.150000 ;
        RECT 760.000000 387.850000 765.000000 388.150000 ;
        RECT 760.000000 383.850000 765.000000 384.150000 ;
        RECT 760.000000 407.850000 765.000000 408.150000 ;
        RECT 760.000000 399.850000 765.000000 400.150000 ;
        RECT 760.000000 403.850000 765.000000 404.150000 ;
        RECT 760.000000 411.850000 765.000000 412.150000 ;
        RECT 760.000000 415.850000 765.000000 416.150000 ;
        RECT 810.000000 387.850000 815.000000 388.150000 ;
        RECT 810.000000 383.850000 815.000000 384.150000 ;
        RECT 810.000000 391.850000 815.000000 392.150000 ;
        RECT 810.000000 395.850000 815.000000 396.150000 ;
        RECT 810.000000 407.850000 815.000000 408.150000 ;
        RECT 810.000000 403.850000 815.000000 404.150000 ;
        RECT 810.000000 399.850000 815.000000 400.150000 ;
        RECT 810.000000 411.850000 815.000000 412.150000 ;
        RECT 810.000000 415.850000 815.000000 416.150000 ;
        RECT 860.000000 379.850000 865.000000 380.150000 ;
        RECT 860.000000 359.850000 865.000000 360.150000 ;
        RECT 860.000000 355.850000 865.000000 356.150000 ;
        RECT 860.000000 351.850000 865.000000 352.150000 ;
        RECT 860.000000 347.850000 865.000000 348.150000 ;
        RECT 860.000000 343.850000 865.000000 344.150000 ;
        RECT 860.000000 375.850000 865.000000 376.150000 ;
        RECT 860.000000 371.850000 865.000000 372.150000 ;
        RECT 860.000000 367.850000 865.000000 368.150000 ;
        RECT 860.000000 363.850000 865.000000 364.150000 ;
        RECT 860.000000 395.850000 865.000000 396.150000 ;
        RECT 860.000000 391.850000 865.000000 392.150000 ;
        RECT 860.000000 387.850000 865.000000 388.150000 ;
        RECT 860.000000 383.850000 865.000000 384.150000 ;
        RECT 860.000000 407.850000 865.000000 408.150000 ;
        RECT 860.000000 403.850000 865.000000 404.150000 ;
        RECT 860.000000 399.850000 865.000000 400.150000 ;
        RECT 860.000000 415.850000 865.000000 416.150000 ;
        RECT 860.000000 411.850000 865.000000 412.150000 ;
        RECT 760.000000 419.850000 765.000000 420.150000 ;
        RECT 760.000000 423.850000 765.000000 424.150000 ;
        RECT 760.000000 427.850000 765.000000 428.150000 ;
        RECT 760.000000 431.850000 765.000000 432.150000 ;
        RECT 760.000000 443.850000 765.000000 444.150000 ;
        RECT 760.000000 439.850000 765.000000 440.150000 ;
        RECT 760.000000 435.850000 765.000000 436.150000 ;
        RECT 810.000000 419.850000 815.000000 420.150000 ;
        RECT 810.000000 423.850000 815.000000 424.150000 ;
        RECT 810.000000 427.850000 815.000000 428.150000 ;
        RECT 810.000000 431.850000 815.000000 432.150000 ;
        RECT 810.000000 439.850000 815.000000 440.150000 ;
        RECT 810.000000 435.850000 815.000000 436.150000 ;
        RECT 810.000000 443.850000 815.000000 444.150000 ;
        RECT 860.000000 419.850000 865.000000 420.150000 ;
        RECT 860.000000 423.850000 865.000000 424.150000 ;
        RECT 860.000000 427.850000 865.000000 428.150000 ;
        RECT 860.000000 431.850000 865.000000 432.150000 ;
        RECT 860.000000 443.850000 865.000000 444.150000 ;
        RECT 860.000000 439.850000 865.000000 440.150000 ;
        RECT 860.000000 435.850000 865.000000 436.150000 ;
        RECT 610.000000 503.850000 615.000000 504.150000 ;
        RECT 610.000000 499.850000 615.000000 500.150000 ;
        RECT 610.000000 491.850000 615.000000 492.150000 ;
        RECT 610.000000 495.850000 615.000000 496.150000 ;
        RECT 660.000000 495.850000 665.000000 496.150000 ;
        RECT 660.000000 491.850000 665.000000 492.150000 ;
        RECT 660.000000 499.850000 665.000000 500.150000 ;
        RECT 660.000000 503.850000 665.000000 504.150000 ;
        RECT 710.000000 503.850000 715.000000 504.150000 ;
        RECT 710.000000 499.850000 715.000000 500.150000 ;
        RECT 710.000000 495.850000 715.000000 496.150000 ;
        RECT 710.000000 491.850000 715.000000 492.150000 ;
        RECT 960.000000 379.850000 965.000000 380.150000 ;
        RECT 960.000000 343.850000 965.000000 344.150000 ;
        RECT 960.000000 347.850000 965.000000 348.150000 ;
        RECT 960.000000 351.850000 965.000000 352.150000 ;
        RECT 960.000000 355.850000 965.000000 356.150000 ;
        RECT 960.000000 359.850000 965.000000 360.150000 ;
        RECT 960.000000 375.850000 965.000000 376.150000 ;
        RECT 960.000000 371.850000 965.000000 372.150000 ;
        RECT 960.000000 367.850000 965.000000 368.150000 ;
        RECT 960.000000 363.850000 965.000000 364.150000 ;
        RECT 960.000000 383.850000 965.000000 384.150000 ;
        RECT 960.000000 387.850000 965.000000 388.150000 ;
        RECT 960.000000 391.850000 965.000000 392.150000 ;
        RECT 960.000000 395.850000 965.000000 396.150000 ;
        RECT 960.000000 407.850000 965.000000 408.150000 ;
        RECT 960.000000 399.850000 965.000000 400.150000 ;
        RECT 960.000000 403.850000 965.000000 404.150000 ;
        RECT 960.000000 411.850000 965.000000 412.150000 ;
        RECT 960.000000 415.850000 965.000000 416.150000 ;
        RECT 910.000000 379.850000 915.000000 380.150000 ;
        RECT 910.000000 343.850000 915.000000 344.150000 ;
        RECT 910.000000 347.850000 915.000000 348.150000 ;
        RECT 910.000000 351.850000 915.000000 352.150000 ;
        RECT 910.000000 355.850000 915.000000 356.150000 ;
        RECT 910.000000 359.850000 915.000000 360.150000 ;
        RECT 910.000000 375.850000 915.000000 376.150000 ;
        RECT 910.000000 371.850000 915.000000 372.150000 ;
        RECT 910.000000 367.850000 915.000000 368.150000 ;
        RECT 910.000000 363.850000 915.000000 364.150000 ;
        RECT 910.000000 383.850000 915.000000 384.150000 ;
        RECT 910.000000 387.850000 915.000000 388.150000 ;
        RECT 910.000000 391.850000 915.000000 392.150000 ;
        RECT 910.000000 395.850000 915.000000 396.150000 ;
        RECT 910.000000 407.850000 915.000000 408.150000 ;
        RECT 910.000000 399.850000 915.000000 400.150000 ;
        RECT 910.000000 403.850000 915.000000 404.150000 ;
        RECT 910.000000 411.850000 915.000000 412.150000 ;
        RECT 910.000000 415.850000 915.000000 416.150000 ;
        RECT 1010.000000 379.850000 1015.000000 380.150000 ;
        RECT 1010.000000 343.850000 1015.000000 344.150000 ;
        RECT 1010.000000 347.850000 1015.000000 348.150000 ;
        RECT 1010.000000 351.850000 1015.000000 352.150000 ;
        RECT 1010.000000 359.850000 1015.000000 360.150000 ;
        RECT 1010.000000 355.850000 1015.000000 356.150000 ;
        RECT 1010.000000 363.850000 1015.000000 364.150000 ;
        RECT 1010.000000 367.850000 1015.000000 368.150000 ;
        RECT 1010.000000 375.850000 1015.000000 376.150000 ;
        RECT 1010.000000 371.850000 1015.000000 372.150000 ;
        RECT 1010.000000 387.850000 1015.000000 388.150000 ;
        RECT 1010.000000 383.850000 1015.000000 384.150000 ;
        RECT 1010.000000 391.850000 1015.000000 392.150000 ;
        RECT 1010.000000 395.850000 1015.000000 396.150000 ;
        RECT 1010.000000 407.850000 1015.000000 408.150000 ;
        RECT 1010.000000 403.850000 1015.000000 404.150000 ;
        RECT 1010.000000 399.850000 1015.000000 400.150000 ;
        RECT 1010.000000 411.850000 1015.000000 412.150000 ;
        RECT 1010.000000 415.850000 1015.000000 416.150000 ;
        RECT 960.000000 431.850000 965.000000 432.150000 ;
        RECT 960.000000 427.850000 965.000000 428.150000 ;
        RECT 960.000000 423.850000 965.000000 424.150000 ;
        RECT 960.000000 419.850000 965.000000 420.150000 ;
        RECT 960.000000 443.850000 965.000000 444.150000 ;
        RECT 960.000000 439.850000 965.000000 440.150000 ;
        RECT 960.000000 435.850000 965.000000 436.150000 ;
        RECT 910.000000 431.850000 915.000000 432.150000 ;
        RECT 910.000000 427.850000 915.000000 428.150000 ;
        RECT 910.000000 423.850000 915.000000 424.150000 ;
        RECT 910.000000 419.850000 915.000000 420.150000 ;
        RECT 910.000000 435.850000 915.000000 436.150000 ;
        RECT 910.000000 439.850000 915.000000 440.150000 ;
        RECT 910.000000 443.850000 915.000000 444.150000 ;
        RECT 1010.000000 419.850000 1015.000000 420.150000 ;
        RECT 1010.000000 423.850000 1015.000000 424.150000 ;
        RECT 1010.000000 427.850000 1015.000000 428.150000 ;
        RECT 1010.000000 431.850000 1015.000000 432.150000 ;
        RECT 1010.000000 435.850000 1015.000000 436.150000 ;
        RECT 1010.000000 439.850000 1015.000000 440.150000 ;
        RECT 1010.000000 443.850000 1015.000000 444.150000 ;
        RECT 1110.000000 379.850000 1115.000000 380.150000 ;
        RECT 1110.000000 343.850000 1115.000000 344.150000 ;
        RECT 1110.000000 347.850000 1115.000000 348.150000 ;
        RECT 1110.000000 351.850000 1115.000000 352.150000 ;
        RECT 1110.000000 355.850000 1115.000000 356.150000 ;
        RECT 1110.000000 359.850000 1115.000000 360.150000 ;
        RECT 1110.000000 375.850000 1115.000000 376.150000 ;
        RECT 1110.000000 371.850000 1115.000000 372.150000 ;
        RECT 1110.000000 367.850000 1115.000000 368.150000 ;
        RECT 1110.000000 363.850000 1115.000000 364.150000 ;
        RECT 1110.000000 383.850000 1115.000000 384.150000 ;
        RECT 1110.000000 387.850000 1115.000000 388.150000 ;
        RECT 1110.000000 391.850000 1115.000000 392.150000 ;
        RECT 1110.000000 395.850000 1115.000000 396.150000 ;
        RECT 1110.000000 407.850000 1115.000000 408.150000 ;
        RECT 1110.000000 399.850000 1115.000000 400.150000 ;
        RECT 1110.000000 403.850000 1115.000000 404.150000 ;
        RECT 1110.000000 411.850000 1115.000000 412.150000 ;
        RECT 1110.000000 415.850000 1115.000000 416.150000 ;
        RECT 1060.000000 379.850000 1065.000000 380.150000 ;
        RECT 1060.000000 343.850000 1065.000000 344.150000 ;
        RECT 1060.000000 347.850000 1065.000000 348.150000 ;
        RECT 1060.000000 351.850000 1065.000000 352.150000 ;
        RECT 1060.000000 355.850000 1065.000000 356.150000 ;
        RECT 1060.000000 359.850000 1065.000000 360.150000 ;
        RECT 1060.000000 375.850000 1065.000000 376.150000 ;
        RECT 1060.000000 371.850000 1065.000000 372.150000 ;
        RECT 1060.000000 367.850000 1065.000000 368.150000 ;
        RECT 1060.000000 363.850000 1065.000000 364.150000 ;
        RECT 1060.000000 383.850000 1065.000000 384.150000 ;
        RECT 1060.000000 387.850000 1065.000000 388.150000 ;
        RECT 1060.000000 391.850000 1065.000000 392.150000 ;
        RECT 1060.000000 395.850000 1065.000000 396.150000 ;
        RECT 1060.000000 407.850000 1065.000000 408.150000 ;
        RECT 1060.000000 399.850000 1065.000000 400.150000 ;
        RECT 1060.000000 403.850000 1065.000000 404.150000 ;
        RECT 1060.000000 411.850000 1065.000000 412.150000 ;
        RECT 1060.000000 415.850000 1065.000000 416.150000 ;
        RECT 1158.000000 379.850000 1168.000000 380.150000 ;
        RECT 1158.000000 343.850000 1168.000000 344.150000 ;
        RECT 1158.000000 347.850000 1168.000000 348.150000 ;
        RECT 1158.000000 351.850000 1168.000000 352.150000 ;
        RECT 1158.000000 355.850000 1168.000000 356.150000 ;
        RECT 1158.000000 359.850000 1168.000000 360.150000 ;
        RECT 1158.000000 375.850000 1168.000000 376.150000 ;
        RECT 1158.000000 371.850000 1168.000000 372.150000 ;
        RECT 1158.000000 367.850000 1168.000000 368.150000 ;
        RECT 1158.000000 363.850000 1168.000000 364.150000 ;
        RECT 1158.000000 383.850000 1168.000000 384.150000 ;
        RECT 1158.000000 387.850000 1168.000000 388.150000 ;
        RECT 1158.000000 391.850000 1168.000000 392.150000 ;
        RECT 1158.000000 395.850000 1168.000000 396.150000 ;
        RECT 1158.000000 407.850000 1168.000000 408.150000 ;
        RECT 1158.000000 399.850000 1168.000000 400.150000 ;
        RECT 1158.000000 403.850000 1168.000000 404.150000 ;
        RECT 1158.000000 411.850000 1168.000000 412.150000 ;
        RECT 1158.000000 415.850000 1168.000000 416.150000 ;
        RECT 1110.000000 431.850000 1115.000000 432.150000 ;
        RECT 1110.000000 427.850000 1115.000000 428.150000 ;
        RECT 1110.000000 423.850000 1115.000000 424.150000 ;
        RECT 1110.000000 419.850000 1115.000000 420.150000 ;
        RECT 1110.000000 443.850000 1115.000000 444.150000 ;
        RECT 1110.000000 439.850000 1115.000000 440.150000 ;
        RECT 1110.000000 435.850000 1115.000000 436.150000 ;
        RECT 1060.000000 419.850000 1065.000000 420.150000 ;
        RECT 1060.000000 423.850000 1065.000000 424.150000 ;
        RECT 1060.000000 431.850000 1065.000000 432.150000 ;
        RECT 1060.000000 427.850000 1065.000000 428.150000 ;
        RECT 1060.000000 435.850000 1065.000000 436.150000 ;
        RECT 1060.000000 439.850000 1065.000000 440.150000 ;
        RECT 1060.000000 443.850000 1065.000000 444.150000 ;
        RECT 1158.000000 427.850000 1168.000000 428.150000 ;
        RECT 1158.000000 423.850000 1168.000000 424.150000 ;
        RECT 1158.000000 419.850000 1168.000000 420.150000 ;
        RECT 1160.000000 431.850000 1165.000000 432.150000 ;
        RECT 1160.000000 435.850000 1165.000000 436.150000 ;
        RECT 1160.000000 439.850000 1165.000000 440.150000 ;
        RECT 1160.000000 443.850000 1165.000000 444.150000 ;
        RECT 1160.000000 447.850000 1165.000000 448.150000 ;
        RECT 1160.000000 451.850000 1165.000000 452.150000 ;
        RECT 1160.000000 459.850000 1165.000000 460.150000 ;
        RECT 1160.000000 455.850000 1165.000000 456.150000 ;
        RECT 1160.000000 463.850000 1165.000000 464.150000 ;
        RECT 1160.000000 467.850000 1165.000000 468.150000 ;
        RECT 1160.000000 471.850000 1165.000000 472.150000 ;
        RECT 1160.000000 479.850000 1165.000000 480.150000 ;
        RECT 1160.000000 475.850000 1165.000000 476.150000 ;
        RECT 1160.000000 487.850000 1165.000000 488.150000 ;
        RECT 1160.000000 483.850000 1165.000000 484.150000 ;
        RECT 1160.000000 491.850000 1165.000000 492.150000 ;
        RECT 1160.000000 495.850000 1165.000000 496.150000 ;
        RECT 1160.000000 499.850000 1165.000000 500.150000 ;
        RECT 1160.000000 507.850000 1165.000000 508.150000 ;
        RECT 1160.000000 503.850000 1165.000000 504.150000 ;
        RECT 1160.000000 511.850000 1165.000000 512.150000 ;
        RECT 1160.000000 515.850000 1165.000000 516.150000 ;
        RECT 1160.000000 519.850000 1165.000000 520.150000 ;
        RECT 1160.000000 523.850000 1165.000000 524.150000 ;
        RECT 1160.000000 527.850000 1165.000000 528.150000 ;
        RECT 1160.000000 535.850000 1165.000000 536.150000 ;
        RECT 1160.000000 531.850000 1165.000000 532.150000 ;
        RECT 1160.000000 539.850000 1165.000000 540.150000 ;
        RECT 1160.000000 543.850000 1165.000000 544.150000 ;
        RECT 1160.000000 555.850000 1165.000000 556.150000 ;
        RECT 1160.000000 551.850000 1165.000000 552.150000 ;
        RECT 1160.000000 547.850000 1165.000000 548.150000 ;
        RECT 1160.000000 563.850000 1165.000000 564.150000 ;
        RECT 1160.000000 559.850000 1165.000000 560.150000 ;
        RECT 1160.000000 583.850000 1165.000000 584.150000 ;
        RECT 1160.000000 567.850000 1165.000000 568.150000 ;
        RECT 1160.000000 571.850000 1165.000000 572.150000 ;
        RECT 1160.000000 579.850000 1165.000000 580.150000 ;
        RECT 1160.000000 575.850000 1165.000000 576.150000 ;
        RECT 1160.000000 591.850000 1165.000000 592.150000 ;
        RECT 1160.000000 587.850000 1165.000000 588.150000 ;
        RECT 1160.000000 595.850000 1165.000000 596.150000 ;
        RECT 1160.000000 599.850000 1165.000000 600.150000 ;
        RECT 1160.000000 607.850000 1165.000000 608.150000 ;
        RECT 1160.000000 603.850000 1165.000000 604.150000 ;
        RECT 1160.000000 611.850000 1165.000000 612.150000 ;
        RECT 1160.000000 615.850000 1165.000000 616.150000 ;
        RECT 1160.000000 619.850000 1165.000000 620.150000 ;
        RECT 1160.000000 623.850000 1165.000000 624.150000 ;
        RECT 1160.000000 627.850000 1165.000000 628.150000 ;
        RECT 1160.000000 635.850000 1165.000000 636.150000 ;
        RECT 1160.000000 631.850000 1165.000000 632.150000 ;
        RECT 610.000000 659.850000 615.000000 660.150000 ;
        RECT 610.000000 663.850000 615.000000 664.150000 ;
        RECT 610.000000 667.850000 615.000000 668.150000 ;
        RECT 610.000000 671.850000 615.000000 672.150000 ;
        RECT 610.000000 675.850000 615.000000 676.150000 ;
        RECT 660.000000 663.850000 665.000000 664.150000 ;
        RECT 660.000000 659.850000 665.000000 660.150000 ;
        RECT 660.000000 667.850000 665.000000 668.150000 ;
        RECT 660.000000 671.850000 665.000000 672.150000 ;
        RECT 660.000000 675.850000 665.000000 676.150000 ;
        RECT 610.000000 683.850000 615.000000 684.150000 ;
        RECT 610.000000 679.850000 615.000000 680.150000 ;
        RECT 660.000000 683.850000 665.000000 684.150000 ;
        RECT 660.000000 679.850000 665.000000 680.150000 ;
        RECT 1160.000000 639.850000 1165.000000 640.150000 ;
        RECT 1160.000000 643.850000 1165.000000 644.150000 ;
        RECT 1160.000000 647.850000 1165.000000 648.150000 ;
        RECT 1160.000000 655.850000 1165.000000 656.150000 ;
        RECT 1160.000000 651.850000 1165.000000 652.150000 ;
        RECT 1160.000000 663.850000 1165.000000 664.150000 ;
        RECT 1160.000000 659.850000 1165.000000 660.150000 ;
        RECT 1160.000000 667.850000 1165.000000 668.150000 ;
        RECT 1160.000000 671.850000 1165.000000 672.150000 ;
        RECT 1160.000000 675.850000 1165.000000 676.150000 ;
        RECT 1160.000000 683.850000 1165.000000 684.150000 ;
        RECT 1160.000000 679.850000 1165.000000 680.150000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  OBS
    LAYER OVERLAP ;
      RECT 0.000000 656.000000 670.000000 686.000000 ;
      RECT 0.000000 506.000000 389.000000 656.000000 ;
      RECT 1139.000000 446.000000 1186.000000 686.000000 ;
      RECT 0.000000 446.000000 739.000000 506.000000 ;
      RECT 0.000000 0.000000 1186.000000 446.000000 ;
    LAYER M1 ;
      RECT 0.000000 656.000000 670.000000 686.000000 ;
      RECT 0.000000 506.000000 389.000000 656.000000 ;
      RECT 1139.000000 446.000000 1186.000000 686.000000 ;
      RECT 0.000000 446.000000 739.000000 506.000000 ;
      RECT 0.000000 0.000000 1186.000000 446.000000 ;
    LAYER M2 ;
      RECT 1139.000000 685.650000 1186.000000 686.000000 ;
      RECT 647.765000 685.650000 670.000000 686.000000 ;
      RECT 561.965000 685.650000 624.430000 686.000000 ;
      RECT 556.285000 685.650000 558.865000 686.000000 ;
      RECT 476.165000 685.650000 538.630000 686.000000 ;
      RECT 455.930000 685.650000 463.425000 686.000000 ;
      RECT 390.365000 685.650000 452.830000 686.000000 ;
      RECT 304.565000 685.650000 367.030000 686.000000 ;
      RECT 647.765000 683.980000 658.500000 685.650000 ;
      RECT 642.085000 683.980000 644.665000 686.000000 ;
      RECT 638.125000 683.980000 638.985000 686.000000 ;
      RECT 627.530000 683.980000 635.025000 686.000000 ;
      RECT 616.500000 683.980000 624.430000 685.650000 ;
      RECT 556.285000 683.980000 558.500000 685.650000 ;
      RECT 552.325000 683.980000 553.185000 686.000000 ;
      RECT 541.730000 683.980000 549.225000 686.000000 ;
      RECT 516.500000 683.980000 538.630000 685.650000 ;
      RECT 476.165000 683.980000 508.500000 685.650000 ;
      RECT 470.485000 683.980000 473.065000 686.000000 ;
      RECT 466.525000 683.980000 467.385000 686.000000 ;
      RECT 455.930000 683.980000 458.500000 685.650000 ;
      RECT 416.500000 683.980000 452.830000 685.650000 ;
      RECT 390.365000 683.980000 408.500000 685.650000 ;
      RECT 384.685000 683.980000 387.265000 686.000000 ;
      RECT 380.725000 683.980000 381.585000 686.000000 ;
      RECT 370.130000 683.980000 377.625000 686.000000 ;
      RECT 366.500000 683.980000 367.030000 685.650000 ;
      RECT 304.565000 683.980000 308.500000 685.650000 ;
      RECT 298.885000 683.980000 301.465000 686.000000 ;
      RECT 294.925000 683.980000 295.785000 686.000000 ;
      RECT 284.330000 683.980000 291.825000 686.000000 ;
      RECT 218.765000 683.980000 281.230000 686.000000 ;
      RECT 213.085000 683.980000 215.665000 686.000000 ;
      RECT 209.125000 683.980000 209.985000 686.000000 ;
      RECT 198.530000 683.980000 206.025000 686.000000 ;
      RECT 132.965000 683.980000 195.430000 686.000000 ;
      RECT 127.285000 683.980000 129.865000 686.000000 ;
      RECT 123.325000 683.980000 124.185000 686.000000 ;
      RECT 112.730000 683.980000 120.225000 686.000000 ;
      RECT 47.165000 683.980000 109.630000 686.000000 ;
      RECT 41.485000 683.980000 44.065000 686.000000 ;
      RECT 37.525000 683.980000 38.385000 686.000000 ;
      RECT 26.930000 683.980000 34.425000 686.000000 ;
      RECT 0.000000 683.980000 23.830000 686.000000 ;
      RECT 1139.000000 683.650000 1158.500000 685.650000 ;
      RECT 616.500000 683.650000 658.500000 683.980000 ;
      RECT 566.500000 683.650000 608.500000 685.650000 ;
      RECT 516.500000 683.650000 558.500000 683.980000 ;
      RECT 466.500000 683.650000 508.500000 683.980000 ;
      RECT 416.500000 683.650000 458.500000 683.980000 ;
      RECT 366.500000 683.650000 408.500000 683.980000 ;
      RECT 316.500000 683.650000 358.500000 685.650000 ;
      RECT 0.000000 683.650000 308.500000 683.980000 ;
      RECT 1166.500000 682.350000 1186.000000 685.650000 ;
      RECT 1157.500000 682.350000 1158.500000 683.650000 ;
      RECT 666.500000 682.350000 670.000000 685.650000 ;
      RECT 657.500000 682.350000 658.500000 683.650000 ;
      RECT 616.500000 682.350000 649.500000 683.650000 ;
      RECT 607.500000 682.350000 608.500000 683.650000 ;
      RECT 566.500000 682.350000 599.500000 683.650000 ;
      RECT 557.500000 682.350000 558.500000 683.650000 ;
      RECT 516.500000 682.350000 549.500000 683.650000 ;
      RECT 507.500000 682.350000 508.500000 683.650000 ;
      RECT 466.500000 682.350000 499.500000 683.650000 ;
      RECT 457.500000 682.350000 458.500000 683.650000 ;
      RECT 416.500000 682.350000 449.500000 683.650000 ;
      RECT 407.500000 682.350000 408.500000 683.650000 ;
      RECT 366.500000 682.350000 373.500000 683.650000 ;
      RECT 357.500000 682.350000 358.500000 683.650000 ;
      RECT 316.500000 682.350000 349.500000 683.650000 ;
      RECT 307.500000 682.350000 308.500000 683.650000 ;
      RECT 1157.500000 681.650000 1186.000000 682.350000 ;
      RECT 657.500000 681.650000 670.000000 682.350000 ;
      RECT 607.500000 681.650000 649.500000 682.350000 ;
      RECT 557.500000 681.650000 599.500000 682.350000 ;
      RECT 507.500000 681.650000 549.500000 682.350000 ;
      RECT 457.500000 681.650000 499.500000 682.350000 ;
      RECT 407.500000 681.650000 449.500000 682.350000 ;
      RECT 357.500000 681.650000 373.500000 682.350000 ;
      RECT 307.500000 681.650000 349.500000 682.350000 ;
      RECT 1157.500000 680.350000 1158.500000 681.650000 ;
      RECT 1139.000000 680.350000 1149.500000 683.650000 ;
      RECT 657.500000 680.350000 658.500000 681.650000 ;
      RECT 616.500000 680.350000 649.500000 681.650000 ;
      RECT 607.500000 680.350000 608.500000 681.650000 ;
      RECT 566.500000 680.350000 599.500000 681.650000 ;
      RECT 557.500000 680.350000 558.500000 681.650000 ;
      RECT 516.500000 680.350000 549.500000 681.650000 ;
      RECT 507.500000 680.350000 508.500000 681.650000 ;
      RECT 466.500000 680.350000 499.500000 681.650000 ;
      RECT 457.500000 680.350000 458.500000 681.650000 ;
      RECT 416.500000 680.350000 449.500000 681.650000 ;
      RECT 407.500000 680.350000 408.500000 681.650000 ;
      RECT 386.500000 680.350000 399.500000 683.650000 ;
      RECT 366.500000 680.350000 373.500000 681.650000 ;
      RECT 357.500000 680.350000 358.500000 681.650000 ;
      RECT 316.500000 680.350000 349.500000 681.650000 ;
      RECT 307.500000 680.350000 308.500000 681.650000 ;
      RECT 0.000000 680.350000 299.500000 683.650000 ;
      RECT 1139.000000 679.650000 1158.500000 680.350000 ;
      RECT 616.500000 679.650000 658.500000 680.350000 ;
      RECT 566.500000 679.650000 608.500000 680.350000 ;
      RECT 516.500000 679.650000 558.500000 680.350000 ;
      RECT 466.500000 679.650000 508.500000 680.350000 ;
      RECT 416.500000 679.650000 458.500000 680.350000 ;
      RECT 366.500000 679.650000 408.500000 680.350000 ;
      RECT 316.500000 679.650000 358.500000 680.350000 ;
      RECT 0.000000 679.650000 308.500000 680.350000 ;
      RECT 1166.500000 678.350000 1186.000000 681.650000 ;
      RECT 1157.500000 678.350000 1158.500000 679.650000 ;
      RECT 666.500000 678.350000 670.000000 681.650000 ;
      RECT 657.500000 678.350000 658.500000 679.650000 ;
      RECT 616.500000 678.350000 649.500000 679.650000 ;
      RECT 607.500000 678.350000 608.500000 679.650000 ;
      RECT 566.500000 678.350000 599.500000 679.650000 ;
      RECT 557.500000 678.350000 558.500000 679.650000 ;
      RECT 516.500000 678.350000 549.500000 679.650000 ;
      RECT 507.500000 678.350000 508.500000 679.650000 ;
      RECT 466.500000 678.350000 499.500000 679.650000 ;
      RECT 457.500000 678.350000 458.500000 679.650000 ;
      RECT 416.500000 678.350000 449.500000 679.650000 ;
      RECT 407.500000 678.350000 408.500000 679.650000 ;
      RECT 366.500000 678.350000 373.500000 679.650000 ;
      RECT 357.500000 678.350000 358.500000 679.650000 ;
      RECT 316.500000 678.350000 349.500000 679.650000 ;
      RECT 307.500000 678.350000 308.500000 679.650000 ;
      RECT 1157.500000 677.650000 1186.000000 678.350000 ;
      RECT 657.500000 677.650000 670.000000 678.350000 ;
      RECT 607.500000 677.650000 649.500000 678.350000 ;
      RECT 557.500000 677.650000 599.500000 678.350000 ;
      RECT 507.500000 677.650000 549.500000 678.350000 ;
      RECT 457.500000 677.650000 499.500000 678.350000 ;
      RECT 407.500000 677.650000 449.500000 678.350000 ;
      RECT 357.500000 677.650000 373.500000 678.350000 ;
      RECT 1157.500000 676.350000 1158.500000 677.650000 ;
      RECT 1139.000000 676.350000 1149.500000 679.650000 ;
      RECT 657.500000 676.350000 658.500000 677.650000 ;
      RECT 616.500000 676.350000 649.500000 677.650000 ;
      RECT 607.500000 676.350000 608.500000 677.650000 ;
      RECT 566.500000 676.350000 599.500000 677.650000 ;
      RECT 557.500000 676.350000 558.500000 677.650000 ;
      RECT 516.500000 676.350000 549.500000 677.650000 ;
      RECT 507.500000 676.350000 508.500000 677.650000 ;
      RECT 466.500000 676.350000 499.500000 677.650000 ;
      RECT 457.500000 676.350000 458.500000 677.650000 ;
      RECT 416.500000 676.350000 449.500000 677.650000 ;
      RECT 407.500000 676.350000 408.500000 677.650000 ;
      RECT 386.500000 676.350000 399.500000 679.650000 ;
      RECT 366.500000 676.350000 373.500000 677.650000 ;
      RECT 357.500000 676.350000 358.500000 677.650000 ;
      RECT 307.500000 676.350000 349.500000 678.350000 ;
      RECT 0.000000 676.350000 299.500000 679.650000 ;
      RECT 1139.000000 675.650000 1158.500000 676.350000 ;
      RECT 616.500000 675.650000 658.500000 676.350000 ;
      RECT 566.500000 675.650000 608.500000 676.350000 ;
      RECT 516.500000 675.650000 558.500000 676.350000 ;
      RECT 466.500000 675.650000 508.500000 676.350000 ;
      RECT 416.500000 675.650000 458.500000 676.350000 ;
      RECT 366.500000 675.650000 408.500000 676.350000 ;
      RECT 0.000000 675.650000 358.500000 676.350000 ;
      RECT 1166.500000 674.350000 1186.000000 677.650000 ;
      RECT 1157.500000 674.350000 1158.500000 675.650000 ;
      RECT 666.500000 674.350000 670.000000 677.650000 ;
      RECT 657.500000 674.350000 658.500000 675.650000 ;
      RECT 616.500000 674.350000 649.500000 675.650000 ;
      RECT 607.500000 674.350000 608.500000 675.650000 ;
      RECT 566.500000 674.350000 599.500000 675.650000 ;
      RECT 557.500000 674.350000 558.500000 675.650000 ;
      RECT 516.500000 674.350000 549.500000 675.650000 ;
      RECT 507.500000 674.350000 508.500000 675.650000 ;
      RECT 466.500000 674.350000 499.500000 675.650000 ;
      RECT 457.500000 674.350000 458.500000 675.650000 ;
      RECT 416.500000 674.350000 449.500000 675.650000 ;
      RECT 407.500000 674.350000 408.500000 675.650000 ;
      RECT 366.500000 674.350000 373.500000 675.650000 ;
      RECT 357.500000 674.350000 358.500000 675.650000 ;
      RECT 1157.500000 673.650000 1186.000000 674.350000 ;
      RECT 657.500000 673.650000 670.000000 674.350000 ;
      RECT 607.500000 673.650000 649.500000 674.350000 ;
      RECT 557.500000 673.650000 599.500000 674.350000 ;
      RECT 507.500000 673.650000 549.500000 674.350000 ;
      RECT 457.500000 673.650000 499.500000 674.350000 ;
      RECT 407.500000 673.650000 449.500000 674.350000 ;
      RECT 357.500000 673.650000 373.500000 674.350000 ;
      RECT 1157.500000 672.350000 1158.500000 673.650000 ;
      RECT 1139.000000 672.350000 1149.500000 675.650000 ;
      RECT 657.500000 672.350000 658.500000 673.650000 ;
      RECT 616.500000 672.350000 649.500000 673.650000 ;
      RECT 607.500000 672.350000 608.500000 673.650000 ;
      RECT 566.500000 672.350000 599.500000 673.650000 ;
      RECT 557.500000 672.350000 558.500000 673.650000 ;
      RECT 516.500000 672.350000 549.500000 673.650000 ;
      RECT 507.500000 672.350000 508.500000 673.650000 ;
      RECT 466.500000 672.350000 499.500000 673.650000 ;
      RECT 457.500000 672.350000 458.500000 673.650000 ;
      RECT 416.500000 672.350000 449.500000 673.650000 ;
      RECT 407.500000 672.350000 408.500000 673.650000 ;
      RECT 386.500000 672.350000 399.500000 675.650000 ;
      RECT 366.500000 672.350000 373.500000 673.650000 ;
      RECT 357.500000 672.350000 358.500000 673.650000 ;
      RECT 0.000000 672.350000 349.500000 675.650000 ;
      RECT 1139.000000 671.650000 1158.500000 672.350000 ;
      RECT 616.500000 671.650000 658.500000 672.350000 ;
      RECT 566.500000 671.650000 608.500000 672.350000 ;
      RECT 516.500000 671.650000 558.500000 672.350000 ;
      RECT 466.500000 671.650000 508.500000 672.350000 ;
      RECT 416.500000 671.650000 458.500000 672.350000 ;
      RECT 366.500000 671.650000 408.500000 672.350000 ;
      RECT 0.000000 671.650000 358.500000 672.350000 ;
      RECT 1166.500000 670.350000 1186.000000 673.650000 ;
      RECT 1157.500000 670.350000 1158.500000 671.650000 ;
      RECT 666.500000 670.350000 670.000000 673.650000 ;
      RECT 657.500000 670.350000 658.500000 671.650000 ;
      RECT 616.500000 670.350000 649.500000 671.650000 ;
      RECT 607.500000 670.350000 608.500000 671.650000 ;
      RECT 566.500000 670.350000 599.500000 671.650000 ;
      RECT 557.500000 670.350000 558.500000 671.650000 ;
      RECT 516.500000 670.350000 549.500000 671.650000 ;
      RECT 507.500000 670.350000 508.500000 671.650000 ;
      RECT 466.500000 670.350000 499.500000 671.650000 ;
      RECT 457.500000 670.350000 458.500000 671.650000 ;
      RECT 416.500000 670.350000 449.500000 671.650000 ;
      RECT 407.500000 670.350000 408.500000 671.650000 ;
      RECT 366.500000 670.350000 373.500000 671.650000 ;
      RECT 357.500000 670.350000 358.500000 671.650000 ;
      RECT 1157.500000 669.650000 1186.000000 670.350000 ;
      RECT 657.500000 669.650000 670.000000 670.350000 ;
      RECT 607.500000 669.650000 649.500000 670.350000 ;
      RECT 557.500000 669.650000 599.500000 670.350000 ;
      RECT 507.500000 669.650000 549.500000 670.350000 ;
      RECT 457.500000 669.650000 499.500000 670.350000 ;
      RECT 407.500000 669.650000 449.500000 670.350000 ;
      RECT 357.500000 669.650000 373.500000 670.350000 ;
      RECT 1157.500000 668.350000 1158.500000 669.650000 ;
      RECT 1139.000000 668.350000 1149.500000 671.650000 ;
      RECT 657.500000 668.350000 658.500000 669.650000 ;
      RECT 616.500000 668.350000 649.500000 669.650000 ;
      RECT 607.500000 668.350000 608.500000 669.650000 ;
      RECT 566.500000 668.350000 599.500000 669.650000 ;
      RECT 557.500000 668.350000 558.500000 669.650000 ;
      RECT 516.500000 668.350000 549.500000 669.650000 ;
      RECT 507.500000 668.350000 508.500000 669.650000 ;
      RECT 466.500000 668.350000 499.500000 669.650000 ;
      RECT 457.500000 668.350000 458.500000 669.650000 ;
      RECT 416.500000 668.350000 449.500000 669.650000 ;
      RECT 407.500000 668.350000 408.500000 669.650000 ;
      RECT 386.500000 668.350000 399.500000 671.650000 ;
      RECT 372.500000 668.350000 373.500000 669.650000 ;
      RECT 357.500000 668.350000 358.500000 669.650000 ;
      RECT 0.000000 668.350000 349.500000 671.650000 ;
      RECT 1139.000000 667.650000 1158.500000 668.350000 ;
      RECT 616.500000 667.650000 658.500000 668.350000 ;
      RECT 566.500000 667.650000 608.500000 668.350000 ;
      RECT 516.500000 667.650000 558.500000 668.350000 ;
      RECT 466.500000 667.650000 508.500000 668.350000 ;
      RECT 416.500000 667.650000 458.500000 668.350000 ;
      RECT 372.500000 667.650000 408.500000 668.350000 ;
      RECT 0.000000 667.650000 358.500000 668.350000 ;
      RECT 1166.500000 666.350000 1186.000000 669.650000 ;
      RECT 1157.500000 666.350000 1158.500000 667.650000 ;
      RECT 666.500000 666.350000 670.000000 669.650000 ;
      RECT 657.500000 666.350000 658.500000 667.650000 ;
      RECT 616.500000 666.350000 649.500000 667.650000 ;
      RECT 607.500000 666.350000 608.500000 667.650000 ;
      RECT 566.500000 666.350000 599.500000 667.650000 ;
      RECT 557.500000 666.350000 558.500000 667.650000 ;
      RECT 516.500000 666.350000 549.500000 667.650000 ;
      RECT 507.500000 666.350000 508.500000 667.650000 ;
      RECT 466.500000 666.350000 499.500000 667.650000 ;
      RECT 457.500000 666.350000 458.500000 667.650000 ;
      RECT 416.500000 666.350000 449.500000 667.650000 ;
      RECT 407.500000 666.350000 408.500000 667.650000 ;
      RECT 372.500000 666.350000 373.500000 667.650000 ;
      RECT 357.500000 666.350000 358.500000 667.650000 ;
      RECT 1157.500000 665.650000 1186.000000 666.350000 ;
      RECT 657.500000 665.650000 670.000000 666.350000 ;
      RECT 607.500000 665.650000 649.500000 666.350000 ;
      RECT 557.500000 665.650000 599.500000 666.350000 ;
      RECT 507.500000 665.650000 549.500000 666.350000 ;
      RECT 457.500000 665.650000 499.500000 666.350000 ;
      RECT 407.500000 665.650000 449.500000 666.350000 ;
      RECT 357.500000 665.650000 373.500000 666.350000 ;
      RECT 1157.500000 664.350000 1158.500000 665.650000 ;
      RECT 1139.000000 664.350000 1149.500000 667.650000 ;
      RECT 657.500000 664.350000 658.500000 665.650000 ;
      RECT 616.500000 664.350000 649.500000 665.650000 ;
      RECT 607.500000 664.350000 608.500000 665.650000 ;
      RECT 566.500000 664.350000 599.500000 665.650000 ;
      RECT 557.500000 664.350000 558.500000 665.650000 ;
      RECT 516.500000 664.350000 549.500000 665.650000 ;
      RECT 507.500000 664.350000 508.500000 665.650000 ;
      RECT 466.500000 664.350000 499.500000 665.650000 ;
      RECT 457.500000 664.350000 458.500000 665.650000 ;
      RECT 416.500000 664.350000 449.500000 665.650000 ;
      RECT 407.500000 664.350000 408.500000 665.650000 ;
      RECT 386.500000 664.350000 399.500000 667.650000 ;
      RECT 372.500000 664.350000 373.500000 665.650000 ;
      RECT 357.500000 664.350000 358.500000 665.650000 ;
      RECT 0.000000 664.350000 349.500000 667.650000 ;
      RECT 1139.000000 663.650000 1158.500000 664.350000 ;
      RECT 616.500000 663.650000 658.500000 664.350000 ;
      RECT 566.500000 663.650000 608.500000 664.350000 ;
      RECT 516.500000 663.650000 558.500000 664.350000 ;
      RECT 466.500000 663.650000 508.500000 664.350000 ;
      RECT 416.500000 663.650000 458.500000 664.350000 ;
      RECT 372.500000 663.650000 408.500000 664.350000 ;
      RECT 0.000000 663.650000 358.500000 664.350000 ;
      RECT 0.000000 663.170000 349.500000 663.650000 ;
      RECT 1166.500000 663.165000 1186.000000 665.650000 ;
      RECT 1166.500000 662.350000 1183.980000 663.165000 ;
      RECT 1157.500000 662.350000 1158.500000 663.650000 ;
      RECT 666.500000 662.350000 670.000000 665.650000 ;
      RECT 657.500000 662.350000 658.500000 663.650000 ;
      RECT 616.500000 662.350000 649.500000 663.650000 ;
      RECT 607.500000 662.350000 608.500000 663.650000 ;
      RECT 566.500000 662.350000 599.500000 663.650000 ;
      RECT 557.500000 662.350000 558.500000 663.650000 ;
      RECT 516.500000 662.350000 549.500000 663.650000 ;
      RECT 507.500000 662.350000 508.500000 663.650000 ;
      RECT 466.500000 662.350000 499.500000 663.650000 ;
      RECT 457.500000 662.350000 458.500000 663.650000 ;
      RECT 416.500000 662.350000 449.500000 663.650000 ;
      RECT 407.500000 662.350000 408.500000 663.650000 ;
      RECT 372.500000 662.350000 373.500000 663.650000 ;
      RECT 357.500000 662.350000 358.500000 663.650000 ;
      RECT 1157.500000 661.650000 1183.980000 662.350000 ;
      RECT 657.500000 661.650000 670.000000 662.350000 ;
      RECT 607.500000 661.650000 649.500000 662.350000 ;
      RECT 557.500000 661.650000 599.500000 662.350000 ;
      RECT 507.500000 661.650000 549.500000 662.350000 ;
      RECT 457.500000 661.650000 499.500000 662.350000 ;
      RECT 407.500000 661.650000 449.500000 662.350000 ;
      RECT 357.500000 661.650000 373.500000 662.350000 ;
      RECT 1157.500000 660.350000 1158.500000 661.650000 ;
      RECT 1139.000000 660.350000 1149.500000 663.650000 ;
      RECT 657.500000 660.350000 658.500000 661.650000 ;
      RECT 616.500000 660.350000 649.500000 661.650000 ;
      RECT 607.500000 660.350000 608.500000 661.650000 ;
      RECT 566.500000 660.350000 599.500000 661.650000 ;
      RECT 557.500000 660.350000 558.500000 661.650000 ;
      RECT 516.500000 660.350000 549.500000 661.650000 ;
      RECT 507.500000 660.350000 508.500000 661.650000 ;
      RECT 466.500000 660.350000 499.500000 661.650000 ;
      RECT 457.500000 660.350000 458.500000 661.650000 ;
      RECT 416.500000 660.350000 449.500000 661.650000 ;
      RECT 407.500000 660.350000 408.500000 661.650000 ;
      RECT 386.500000 660.350000 399.500000 663.650000 ;
      RECT 372.500000 660.350000 373.500000 661.650000 ;
      RECT 357.500000 660.350000 358.500000 661.650000 ;
      RECT 2.020000 660.350000 349.500000 663.170000 ;
      RECT 2.020000 660.070000 358.500000 660.350000 ;
      RECT 1166.500000 660.065000 1183.980000 661.650000 ;
      RECT 1139.000000 659.650000 1158.500000 660.350000 ;
      RECT 616.500000 659.650000 658.500000 660.350000 ;
      RECT 566.500000 659.650000 608.500000 660.350000 ;
      RECT 516.500000 659.650000 558.500000 660.350000 ;
      RECT 466.500000 659.650000 508.500000 660.350000 ;
      RECT 416.500000 659.650000 458.500000 660.350000 ;
      RECT 372.500000 659.650000 408.500000 660.350000 ;
      RECT 0.000000 659.650000 358.500000 660.070000 ;
      RECT 1166.500000 658.350000 1186.000000 660.065000 ;
      RECT 1157.500000 658.350000 1158.500000 659.650000 ;
      RECT 666.500000 658.350000 670.000000 661.650000 ;
      RECT 657.500000 658.350000 658.500000 659.650000 ;
      RECT 616.500000 658.350000 649.500000 659.650000 ;
      RECT 607.500000 658.350000 608.500000 659.650000 ;
      RECT 566.500000 658.350000 599.500000 659.650000 ;
      RECT 557.500000 658.350000 558.500000 659.650000 ;
      RECT 516.500000 658.350000 549.500000 659.650000 ;
      RECT 507.500000 658.350000 508.500000 659.650000 ;
      RECT 466.500000 658.350000 499.500000 659.650000 ;
      RECT 457.500000 658.350000 458.500000 659.650000 ;
      RECT 416.500000 658.350000 449.500000 659.650000 ;
      RECT 407.500000 658.350000 408.500000 659.650000 ;
      RECT 372.500000 658.350000 373.500000 659.650000 ;
      RECT 357.500000 658.350000 358.500000 659.650000 ;
      RECT 1157.500000 657.650000 1186.000000 658.350000 ;
      RECT 357.500000 657.650000 373.500000 658.350000 ;
      RECT 1166.500000 657.485000 1186.000000 657.650000 ;
      RECT 1157.500000 656.350000 1158.500000 657.650000 ;
      RECT 1139.000000 656.350000 1149.500000 659.650000 ;
      RECT 657.500000 656.350000 670.000000 658.350000 ;
      RECT 607.500000 656.350000 649.500000 658.350000 ;
      RECT 557.500000 656.350000 599.500000 658.350000 ;
      RECT 507.500000 656.350000 549.500000 658.350000 ;
      RECT 457.500000 656.350000 499.500000 658.350000 ;
      RECT 407.500000 656.350000 449.500000 658.350000 ;
      RECT 386.500000 656.350000 399.500000 659.650000 ;
      RECT 372.500000 656.350000 373.500000 657.650000 ;
      RECT 357.500000 656.350000 358.500000 657.650000 ;
      RECT 0.000000 656.350000 349.500000 659.650000 ;
      RECT 372.500000 656.000000 670.000000 656.350000 ;
      RECT 1139.000000 655.650000 1158.500000 656.350000 ;
      RECT 372.500000 655.650000 389.000000 656.000000 ;
      RECT 0.000000 655.650000 358.500000 656.350000 ;
      RECT 1166.500000 654.385000 1183.980000 657.485000 ;
      RECT 1166.500000 654.350000 1186.000000 654.385000 ;
      RECT 1157.500000 654.350000 1158.500000 655.650000 ;
      RECT 372.500000 654.350000 373.500000 655.650000 ;
      RECT 357.500000 654.350000 358.500000 655.650000 ;
      RECT 1157.500000 653.650000 1186.000000 654.350000 ;
      RECT 357.500000 653.650000 373.500000 654.350000 ;
      RECT 1166.500000 653.525000 1186.000000 653.650000 ;
      RECT 0.000000 652.575000 349.500000 655.650000 ;
      RECT 1157.500000 652.350000 1158.500000 653.650000 ;
      RECT 1139.000000 652.350000 1149.500000 655.650000 ;
      RECT 386.500000 652.350000 389.000000 655.650000 ;
      RECT 372.500000 652.350000 373.500000 653.650000 ;
      RECT 357.500000 652.350000 358.500000 653.650000 ;
      RECT 2.020000 652.350000 349.500000 652.575000 ;
      RECT 1139.000000 651.650000 1158.500000 652.350000 ;
      RECT 372.500000 651.650000 389.000000 652.350000 ;
      RECT 2.020000 651.650000 358.500000 652.350000 ;
      RECT 1166.500000 650.425000 1183.980000 653.525000 ;
      RECT 1166.500000 650.350000 1186.000000 650.425000 ;
      RECT 1157.500000 650.350000 1158.500000 651.650000 ;
      RECT 372.500000 650.350000 373.500000 651.650000 ;
      RECT 357.500000 650.350000 358.500000 651.650000 ;
      RECT 1157.500000 649.650000 1186.000000 650.350000 ;
      RECT 357.500000 649.650000 373.500000 650.350000 ;
      RECT 2.020000 649.475000 349.500000 651.650000 ;
      RECT 0.000000 648.615000 349.500000 649.475000 ;
      RECT 1157.500000 648.350000 1158.500000 649.650000 ;
      RECT 1139.000000 648.350000 1149.500000 651.650000 ;
      RECT 386.500000 648.350000 389.000000 651.650000 ;
      RECT 372.500000 648.350000 373.500000 649.650000 ;
      RECT 357.500000 648.350000 358.500000 649.650000 ;
      RECT 2.020000 648.350000 349.500000 648.615000 ;
      RECT 1139.000000 647.650000 1158.500000 648.350000 ;
      RECT 372.500000 647.650000 389.000000 648.350000 ;
      RECT 2.020000 647.650000 358.500000 648.350000 ;
      RECT 1166.500000 646.350000 1186.000000 649.650000 ;
      RECT 1157.500000 646.350000 1158.500000 647.650000 ;
      RECT 372.500000 646.350000 373.500000 647.650000 ;
      RECT 357.500000 646.350000 358.500000 647.650000 ;
      RECT 1157.500000 645.650000 1186.000000 646.350000 ;
      RECT 357.500000 645.650000 373.500000 646.350000 ;
      RECT 2.020000 645.515000 349.500000 647.650000 ;
      RECT 1157.500000 644.350000 1158.500000 645.650000 ;
      RECT 1139.000000 644.350000 1149.500000 647.650000 ;
      RECT 386.500000 644.350000 389.000000 647.650000 ;
      RECT 372.500000 644.350000 373.500000 645.650000 ;
      RECT 357.500000 644.350000 358.500000 645.650000 ;
      RECT 0.000000 644.350000 349.500000 645.515000 ;
      RECT 1139.000000 643.650000 1158.500000 644.350000 ;
      RECT 372.500000 643.650000 389.000000 644.350000 ;
      RECT 0.000000 643.650000 358.500000 644.350000 ;
      RECT 0.000000 642.935000 349.500000 643.650000 ;
      RECT 1166.500000 642.930000 1186.000000 645.650000 ;
      RECT 1166.500000 642.350000 1183.980000 642.930000 ;
      RECT 1157.500000 642.350000 1158.500000 643.650000 ;
      RECT 372.500000 642.350000 373.500000 643.650000 ;
      RECT 357.500000 642.350000 358.500000 643.650000 ;
      RECT 1157.500000 641.650000 1183.980000 642.350000 ;
      RECT 357.500000 641.650000 373.500000 642.350000 ;
      RECT 1157.500000 640.350000 1158.500000 641.650000 ;
      RECT 1139.000000 640.350000 1149.500000 643.650000 ;
      RECT 386.500000 640.350000 389.000000 643.650000 ;
      RECT 372.500000 640.350000 373.500000 641.650000 ;
      RECT 357.500000 640.350000 358.500000 641.650000 ;
      RECT 2.020000 640.350000 349.500000 642.935000 ;
      RECT 2.020000 639.835000 358.500000 640.350000 ;
      RECT 1166.500000 639.830000 1183.980000 641.650000 ;
      RECT 1139.000000 639.650000 1158.500000 640.350000 ;
      RECT 372.500000 639.650000 389.000000 640.350000 ;
      RECT 0.000000 639.650000 358.500000 639.835000 ;
      RECT 1166.500000 638.350000 1186.000000 639.830000 ;
      RECT 1157.500000 638.350000 1158.500000 639.650000 ;
      RECT 372.500000 638.350000 373.500000 639.650000 ;
      RECT 357.500000 638.350000 358.500000 639.650000 ;
      RECT 1157.500000 637.650000 1186.000000 638.350000 ;
      RECT 357.500000 637.650000 373.500000 638.350000 ;
      RECT 1157.500000 636.350000 1158.500000 637.650000 ;
      RECT 1139.000000 636.350000 1149.500000 639.650000 ;
      RECT 386.500000 636.350000 389.000000 639.650000 ;
      RECT 372.500000 636.350000 373.500000 637.650000 ;
      RECT 357.500000 636.350000 358.500000 637.650000 ;
      RECT 0.000000 636.350000 349.500000 639.650000 ;
      RECT 1139.000000 635.650000 1158.500000 636.350000 ;
      RECT 372.500000 635.650000 389.000000 636.350000 ;
      RECT 0.000000 635.650000 358.500000 636.350000 ;
      RECT 1166.500000 634.350000 1186.000000 637.650000 ;
      RECT 1157.500000 634.350000 1158.500000 635.650000 ;
      RECT 372.500000 634.350000 373.500000 635.650000 ;
      RECT 357.500000 634.350000 358.500000 635.650000 ;
      RECT 1157.500000 633.650000 1186.000000 634.350000 ;
      RECT 357.500000 633.650000 373.500000 634.350000 ;
      RECT 1157.500000 632.350000 1158.500000 633.650000 ;
      RECT 1139.000000 632.350000 1149.500000 635.650000 ;
      RECT 386.500000 632.350000 389.000000 635.650000 ;
      RECT 372.500000 632.350000 373.500000 633.650000 ;
      RECT 357.500000 632.350000 358.500000 633.650000 ;
      RECT 0.000000 632.350000 349.500000 635.650000 ;
      RECT 1139.000000 631.650000 1158.500000 632.350000 ;
      RECT 372.500000 631.650000 389.000000 632.350000 ;
      RECT 0.000000 631.650000 358.500000 632.350000 ;
      RECT 1166.500000 630.350000 1186.000000 633.650000 ;
      RECT 1157.500000 630.350000 1158.500000 631.650000 ;
      RECT 372.500000 630.350000 373.500000 631.650000 ;
      RECT 357.500000 630.350000 358.500000 631.650000 ;
      RECT 1157.500000 629.650000 1186.000000 630.350000 ;
      RECT 357.500000 629.650000 373.500000 630.350000 ;
      RECT 1157.500000 628.350000 1158.500000 629.650000 ;
      RECT 1139.000000 628.350000 1149.500000 631.650000 ;
      RECT 386.500000 628.350000 389.000000 631.650000 ;
      RECT 372.500000 628.350000 373.500000 629.650000 ;
      RECT 357.500000 628.350000 358.500000 629.650000 ;
      RECT 0.000000 628.350000 349.500000 631.650000 ;
      RECT 1139.000000 627.650000 1158.500000 628.350000 ;
      RECT 372.500000 627.650000 389.000000 628.350000 ;
      RECT 0.000000 627.650000 358.500000 628.350000 ;
      RECT 1166.500000 626.350000 1186.000000 629.650000 ;
      RECT 1157.500000 626.350000 1158.500000 627.650000 ;
      RECT 372.500000 626.350000 373.500000 627.650000 ;
      RECT 357.500000 626.350000 358.500000 627.650000 ;
      RECT 1157.500000 625.650000 1186.000000 626.350000 ;
      RECT 357.500000 625.650000 373.500000 626.350000 ;
      RECT 1157.500000 624.350000 1158.500000 625.650000 ;
      RECT 1139.000000 624.350000 1149.500000 627.650000 ;
      RECT 386.500000 624.350000 389.000000 627.650000 ;
      RECT 372.500000 624.350000 373.500000 625.650000 ;
      RECT 357.500000 624.350000 358.500000 625.650000 ;
      RECT 0.000000 624.350000 349.500000 627.650000 ;
      RECT 1139.000000 623.650000 1158.500000 624.350000 ;
      RECT 372.500000 623.650000 389.000000 624.350000 ;
      RECT 0.000000 623.650000 358.500000 624.350000 ;
      RECT 1166.500000 622.350000 1186.000000 625.650000 ;
      RECT 1157.500000 622.350000 1158.500000 623.650000 ;
      RECT 372.500000 622.350000 373.500000 623.650000 ;
      RECT 357.500000 622.350000 358.500000 623.650000 ;
      RECT 1157.500000 621.650000 1186.000000 622.350000 ;
      RECT 357.500000 621.650000 373.500000 622.350000 ;
      RECT 1157.500000 620.350000 1158.500000 621.650000 ;
      RECT 1139.000000 620.350000 1149.500000 623.650000 ;
      RECT 386.500000 620.350000 389.000000 623.650000 ;
      RECT 372.500000 620.350000 373.500000 621.650000 ;
      RECT 357.500000 620.350000 358.500000 621.650000 ;
      RECT 0.000000 620.350000 349.500000 623.650000 ;
      RECT 1139.000000 619.650000 1158.500000 620.350000 ;
      RECT 372.500000 619.650000 389.000000 620.350000 ;
      RECT 0.000000 619.650000 358.500000 620.350000 ;
      RECT 1166.500000 618.350000 1186.000000 621.650000 ;
      RECT 1157.500000 618.350000 1158.500000 619.650000 ;
      RECT 372.500000 618.350000 373.500000 619.650000 ;
      RECT 357.500000 618.350000 358.500000 619.650000 ;
      RECT 1157.500000 617.650000 1186.000000 618.350000 ;
      RECT 357.500000 617.650000 373.500000 618.350000 ;
      RECT 1157.500000 616.350000 1158.500000 617.650000 ;
      RECT 1139.000000 616.350000 1149.500000 619.650000 ;
      RECT 386.500000 616.350000 389.000000 619.650000 ;
      RECT 372.500000 616.350000 373.500000 617.650000 ;
      RECT 357.500000 616.350000 358.500000 617.650000 ;
      RECT 0.000000 616.350000 349.500000 619.650000 ;
      RECT 372.500000 616.115000 389.000000 616.350000 ;
      RECT 1139.000000 615.695000 1158.500000 616.350000 ;
      RECT 1141.020000 615.650000 1158.500000 615.695000 ;
      RECT 372.500000 615.650000 386.980000 616.115000 ;
      RECT 0.000000 615.650000 358.500000 616.350000 ;
      RECT 1166.500000 614.350000 1186.000000 617.650000 ;
      RECT 1157.500000 614.350000 1158.500000 615.650000 ;
      RECT 372.500000 614.350000 373.500000 615.650000 ;
      RECT 357.500000 614.350000 358.500000 615.650000 ;
      RECT 1157.500000 613.650000 1186.000000 614.350000 ;
      RECT 357.500000 613.650000 373.500000 614.350000 ;
      RECT 1157.500000 612.350000 1158.500000 613.650000 ;
      RECT 1141.020000 612.350000 1149.500000 615.650000 ;
      RECT 386.500000 612.350000 386.980000 615.650000 ;
      RECT 372.500000 612.350000 373.500000 613.650000 ;
      RECT 357.500000 612.350000 358.500000 613.650000 ;
      RECT 0.000000 612.350000 349.500000 615.650000 ;
      RECT 1141.020000 611.650000 1158.500000 612.350000 ;
      RECT 372.500000 611.650000 386.980000 612.350000 ;
      RECT 0.000000 611.650000 358.500000 612.350000 ;
      RECT 1166.500000 610.350000 1186.000000 613.650000 ;
      RECT 1157.500000 610.350000 1158.500000 611.650000 ;
      RECT 372.500000 610.350000 373.500000 611.650000 ;
      RECT 357.500000 610.350000 358.500000 611.650000 ;
      RECT 1157.500000 609.650000 1186.000000 610.350000 ;
      RECT 357.500000 609.650000 373.500000 610.350000 ;
      RECT 1157.500000 608.350000 1158.500000 609.650000 ;
      RECT 1141.020000 608.350000 1149.500000 611.650000 ;
      RECT 386.500000 608.350000 386.980000 611.650000 ;
      RECT 372.500000 608.350000 373.500000 609.650000 ;
      RECT 357.500000 608.350000 358.500000 609.650000 ;
      RECT 0.000000 608.350000 349.500000 611.650000 ;
      RECT 1141.020000 607.650000 1158.500000 608.350000 ;
      RECT 372.500000 607.650000 386.980000 608.350000 ;
      RECT 0.000000 607.650000 358.500000 608.350000 ;
      RECT 1166.500000 606.350000 1186.000000 609.650000 ;
      RECT 1157.500000 606.350000 1158.500000 607.650000 ;
      RECT 372.500000 606.350000 373.500000 607.650000 ;
      RECT 357.500000 606.350000 358.500000 607.650000 ;
      RECT 1157.500000 605.650000 1186.000000 606.350000 ;
      RECT 357.500000 605.650000 373.500000 606.350000 ;
      RECT 1157.500000 604.350000 1158.500000 605.650000 ;
      RECT 1141.020000 604.350000 1149.500000 607.650000 ;
      RECT 386.500000 604.350000 386.980000 607.650000 ;
      RECT 372.500000 604.350000 373.500000 605.650000 ;
      RECT 357.500000 604.350000 358.500000 605.650000 ;
      RECT 0.000000 604.350000 349.500000 607.650000 ;
      RECT 1141.020000 603.650000 1158.500000 604.350000 ;
      RECT 372.500000 603.650000 386.980000 604.350000 ;
      RECT 0.000000 603.650000 358.500000 604.350000 ;
      RECT 1166.500000 602.350000 1186.000000 605.650000 ;
      RECT 1157.500000 602.350000 1158.500000 603.650000 ;
      RECT 372.500000 602.350000 373.500000 603.650000 ;
      RECT 357.500000 602.350000 358.500000 603.650000 ;
      RECT 1157.500000 601.650000 1186.000000 602.350000 ;
      RECT 357.500000 601.650000 373.500000 602.350000 ;
      RECT 1157.500000 600.350000 1158.500000 601.650000 ;
      RECT 1141.020000 600.350000 1149.500000 603.650000 ;
      RECT 386.500000 600.350000 386.980000 603.650000 ;
      RECT 372.500000 600.350000 373.500000 601.650000 ;
      RECT 357.500000 600.350000 358.500000 601.650000 ;
      RECT 0.000000 600.350000 349.500000 603.650000 ;
      RECT 1141.020000 599.650000 1158.500000 600.350000 ;
      RECT 372.500000 599.650000 386.980000 600.350000 ;
      RECT 0.000000 599.650000 358.500000 600.350000 ;
      RECT 1166.500000 598.350000 1186.000000 601.650000 ;
      RECT 1157.500000 598.350000 1158.500000 599.650000 ;
      RECT 372.500000 598.350000 373.500000 599.650000 ;
      RECT 357.500000 598.350000 358.500000 599.650000 ;
      RECT 1141.020000 597.880000 1149.500000 599.650000 ;
      RECT 1157.500000 597.650000 1186.000000 598.350000 ;
      RECT 357.500000 597.650000 373.500000 598.350000 ;
      RECT 1157.500000 596.350000 1158.500000 597.650000 ;
      RECT 1139.000000 596.350000 1149.500000 597.880000 ;
      RECT 386.500000 596.350000 386.980000 599.650000 ;
      RECT 372.500000 596.350000 373.500000 597.650000 ;
      RECT 357.500000 596.350000 358.500000 597.650000 ;
      RECT 0.000000 596.350000 349.500000 599.650000 ;
      RECT 1139.000000 595.650000 1158.500000 596.350000 ;
      RECT 372.500000 595.650000 386.980000 596.350000 ;
      RECT 0.000000 595.650000 358.500000 596.350000 ;
      RECT 1166.500000 594.350000 1186.000000 597.650000 ;
      RECT 1157.500000 594.350000 1158.500000 595.650000 ;
      RECT 372.500000 594.350000 373.500000 595.650000 ;
      RECT 357.500000 594.350000 358.500000 595.650000 ;
      RECT 1157.500000 593.650000 1186.000000 594.350000 ;
      RECT 357.500000 593.650000 373.500000 594.350000 ;
      RECT 1157.500000 592.350000 1158.500000 593.650000 ;
      RECT 1139.000000 592.350000 1149.500000 595.650000 ;
      RECT 386.500000 592.350000 386.980000 595.650000 ;
      RECT 372.500000 592.350000 373.500000 593.650000 ;
      RECT 357.500000 592.350000 358.500000 593.650000 ;
      RECT 0.000000 592.350000 349.500000 595.650000 ;
      RECT 1139.000000 591.650000 1158.500000 592.350000 ;
      RECT 372.500000 591.650000 386.980000 592.350000 ;
      RECT 0.000000 591.650000 358.500000 592.350000 ;
      RECT 1166.500000 590.350000 1186.000000 593.650000 ;
      RECT 1157.500000 590.350000 1158.500000 591.650000 ;
      RECT 372.500000 590.350000 373.500000 591.650000 ;
      RECT 357.500000 590.350000 358.500000 591.650000 ;
      RECT 1157.500000 589.650000 1186.000000 590.350000 ;
      RECT 357.500000 589.650000 373.500000 590.350000 ;
      RECT 1157.500000 588.350000 1158.500000 589.650000 ;
      RECT 1139.000000 588.350000 1149.500000 591.650000 ;
      RECT 386.500000 588.350000 386.980000 591.650000 ;
      RECT 372.500000 588.350000 373.500000 589.650000 ;
      RECT 357.500000 588.350000 358.500000 589.650000 ;
      RECT 0.000000 588.350000 349.500000 591.650000 ;
      RECT 1139.000000 587.650000 1158.500000 588.350000 ;
      RECT 372.500000 587.650000 386.980000 588.350000 ;
      RECT 0.000000 587.650000 358.500000 588.350000 ;
      RECT 1166.500000 586.350000 1186.000000 589.650000 ;
      RECT 1157.500000 586.350000 1158.500000 587.650000 ;
      RECT 372.500000 586.350000 373.500000 587.650000 ;
      RECT 357.500000 586.350000 358.500000 587.650000 ;
      RECT 1157.500000 585.650000 1186.000000 586.350000 ;
      RECT 357.500000 585.650000 373.500000 586.350000 ;
      RECT 1157.500000 584.350000 1158.500000 585.650000 ;
      RECT 1139.000000 584.350000 1149.500000 587.650000 ;
      RECT 386.500000 584.350000 386.980000 587.650000 ;
      RECT 372.500000 584.350000 373.500000 585.650000 ;
      RECT 357.500000 584.350000 358.500000 585.650000 ;
      RECT 0.000000 584.350000 349.500000 587.650000 ;
      RECT 1139.000000 583.650000 1158.500000 584.350000 ;
      RECT 372.500000 583.650000 386.980000 584.350000 ;
      RECT 0.000000 583.650000 358.500000 584.350000 ;
      RECT 1166.500000 582.350000 1186.000000 585.650000 ;
      RECT 1157.500000 582.350000 1158.500000 583.650000 ;
      RECT 372.500000 582.350000 373.500000 583.650000 ;
      RECT 357.500000 582.350000 358.500000 583.650000 ;
      RECT 1157.500000 581.650000 1186.000000 582.350000 ;
      RECT 357.500000 581.650000 373.500000 582.350000 ;
      RECT 1157.500000 580.350000 1158.500000 581.650000 ;
      RECT 1139.000000 580.350000 1149.500000 583.650000 ;
      RECT 386.500000 580.350000 386.980000 583.650000 ;
      RECT 372.500000 580.350000 373.500000 581.650000 ;
      RECT 357.500000 580.350000 358.500000 581.650000 ;
      RECT 0.000000 580.350000 349.500000 583.650000 ;
      RECT 1139.000000 579.650000 1158.500000 580.350000 ;
      RECT 372.500000 579.650000 386.980000 580.350000 ;
      RECT 0.000000 579.650000 358.500000 580.350000 ;
      RECT 1166.500000 578.350000 1186.000000 581.650000 ;
      RECT 1157.500000 578.350000 1158.500000 579.650000 ;
      RECT 372.500000 578.350000 373.500000 579.650000 ;
      RECT 357.500000 578.350000 358.500000 579.650000 ;
      RECT 1157.500000 577.650000 1186.000000 578.350000 ;
      RECT 357.500000 577.650000 373.500000 578.350000 ;
      RECT 386.500000 577.590000 386.980000 579.650000 ;
      RECT 1157.500000 576.350000 1158.500000 577.650000 ;
      RECT 1139.000000 576.350000 1149.500000 579.650000 ;
      RECT 386.500000 576.350000 389.000000 577.590000 ;
      RECT 372.500000 576.350000 373.500000 577.650000 ;
      RECT 357.500000 576.350000 358.500000 577.650000 ;
      RECT 0.000000 576.350000 349.500000 579.650000 ;
      RECT 1139.000000 575.650000 1158.500000 576.350000 ;
      RECT 372.500000 575.650000 389.000000 576.350000 ;
      RECT 0.000000 575.650000 358.500000 576.350000 ;
      RECT 0.000000 575.170000 349.500000 575.650000 ;
      RECT 1166.500000 575.165000 1186.000000 577.650000 ;
      RECT 1166.500000 574.350000 1183.980000 575.165000 ;
      RECT 1157.500000 574.350000 1158.500000 575.650000 ;
      RECT 372.500000 574.350000 373.500000 575.650000 ;
      RECT 357.500000 574.350000 358.500000 575.650000 ;
      RECT 1157.500000 573.650000 1183.980000 574.350000 ;
      RECT 357.500000 573.650000 373.500000 574.350000 ;
      RECT 1157.500000 572.350000 1158.500000 573.650000 ;
      RECT 1139.000000 572.350000 1149.500000 575.650000 ;
      RECT 386.500000 572.350000 389.000000 575.650000 ;
      RECT 372.500000 572.350000 373.500000 573.650000 ;
      RECT 357.500000 572.350000 358.500000 573.650000 ;
      RECT 2.020000 572.350000 349.500000 575.170000 ;
      RECT 2.020000 572.070000 358.500000 572.350000 ;
      RECT 1166.500000 572.065000 1183.980000 573.650000 ;
      RECT 1139.000000 571.650000 1158.500000 572.350000 ;
      RECT 372.500000 571.650000 389.000000 572.350000 ;
      RECT 0.000000 571.650000 358.500000 572.070000 ;
      RECT 1166.500000 570.350000 1186.000000 572.065000 ;
      RECT 1157.500000 570.350000 1158.500000 571.650000 ;
      RECT 372.500000 570.350000 373.500000 571.650000 ;
      RECT 357.500000 570.350000 358.500000 571.650000 ;
      RECT 1157.500000 569.650000 1186.000000 570.350000 ;
      RECT 357.500000 569.650000 373.500000 570.350000 ;
      RECT 1166.500000 569.485000 1186.000000 569.650000 ;
      RECT 1157.500000 568.350000 1158.500000 569.650000 ;
      RECT 1139.000000 568.350000 1149.500000 571.650000 ;
      RECT 386.500000 568.350000 389.000000 571.650000 ;
      RECT 372.500000 568.350000 373.500000 569.650000 ;
      RECT 357.500000 568.350000 358.500000 569.650000 ;
      RECT 0.000000 568.350000 349.500000 571.650000 ;
      RECT 1139.000000 567.650000 1158.500000 568.350000 ;
      RECT 372.500000 567.650000 389.000000 568.350000 ;
      RECT 0.000000 567.650000 358.500000 568.350000 ;
      RECT 1166.500000 566.385000 1183.980000 569.485000 ;
      RECT 1166.500000 566.350000 1186.000000 566.385000 ;
      RECT 1157.500000 566.350000 1158.500000 567.650000 ;
      RECT 372.500000 566.350000 373.500000 567.650000 ;
      RECT 357.500000 566.350000 358.500000 567.650000 ;
      RECT 1157.500000 565.650000 1186.000000 566.350000 ;
      RECT 357.500000 565.650000 373.500000 566.350000 ;
      RECT 1166.500000 565.525000 1186.000000 565.650000 ;
      RECT 0.000000 564.575000 349.500000 567.650000 ;
      RECT 1157.500000 564.350000 1158.500000 565.650000 ;
      RECT 1139.000000 564.350000 1149.500000 567.650000 ;
      RECT 386.500000 564.350000 389.000000 567.650000 ;
      RECT 372.500000 564.350000 373.500000 565.650000 ;
      RECT 357.500000 564.350000 358.500000 565.650000 ;
      RECT 2.020000 564.350000 349.500000 564.575000 ;
      RECT 1139.000000 563.650000 1158.500000 564.350000 ;
      RECT 372.500000 563.650000 389.000000 564.350000 ;
      RECT 2.020000 563.650000 358.500000 564.350000 ;
      RECT 1166.500000 562.425000 1183.980000 565.525000 ;
      RECT 1166.500000 562.350000 1186.000000 562.425000 ;
      RECT 1157.500000 562.350000 1158.500000 563.650000 ;
      RECT 372.500000 562.350000 373.500000 563.650000 ;
      RECT 357.500000 562.350000 358.500000 563.650000 ;
      RECT 1157.500000 561.650000 1186.000000 562.350000 ;
      RECT 357.500000 561.650000 373.500000 562.350000 ;
      RECT 2.020000 561.475000 349.500000 563.650000 ;
      RECT 0.000000 560.615000 349.500000 561.475000 ;
      RECT 1157.500000 560.350000 1158.500000 561.650000 ;
      RECT 1139.000000 560.350000 1149.500000 563.650000 ;
      RECT 386.500000 560.350000 389.000000 563.650000 ;
      RECT 372.500000 560.350000 373.500000 561.650000 ;
      RECT 357.500000 560.350000 358.500000 561.650000 ;
      RECT 2.020000 560.350000 349.500000 560.615000 ;
      RECT 1139.000000 559.650000 1158.500000 560.350000 ;
      RECT 372.500000 559.650000 389.000000 560.350000 ;
      RECT 2.020000 559.650000 358.500000 560.350000 ;
      RECT 1166.500000 558.350000 1186.000000 561.650000 ;
      RECT 1157.500000 558.350000 1158.500000 559.650000 ;
      RECT 372.500000 558.350000 373.500000 559.650000 ;
      RECT 357.500000 558.350000 358.500000 559.650000 ;
      RECT 1157.500000 557.650000 1186.000000 558.350000 ;
      RECT 357.500000 557.650000 373.500000 558.350000 ;
      RECT 2.020000 557.515000 349.500000 559.650000 ;
      RECT 1157.500000 556.350000 1158.500000 557.650000 ;
      RECT 1139.000000 556.350000 1149.500000 559.650000 ;
      RECT 386.500000 556.350000 389.000000 559.650000 ;
      RECT 372.500000 556.350000 373.500000 557.650000 ;
      RECT 357.500000 556.350000 358.500000 557.650000 ;
      RECT 0.000000 556.350000 349.500000 557.515000 ;
      RECT 1139.000000 555.650000 1158.500000 556.350000 ;
      RECT 372.500000 555.650000 389.000000 556.350000 ;
      RECT 0.000000 555.650000 358.500000 556.350000 ;
      RECT 0.000000 554.935000 349.500000 555.650000 ;
      RECT 1166.500000 554.930000 1186.000000 557.650000 ;
      RECT 1166.500000 554.350000 1183.980000 554.930000 ;
      RECT 1157.500000 554.350000 1158.500000 555.650000 ;
      RECT 372.500000 554.350000 373.500000 555.650000 ;
      RECT 357.500000 554.350000 358.500000 555.650000 ;
      RECT 1157.500000 553.650000 1183.980000 554.350000 ;
      RECT 357.500000 553.650000 373.500000 554.350000 ;
      RECT 1157.500000 552.350000 1158.500000 553.650000 ;
      RECT 1139.000000 552.350000 1149.500000 555.650000 ;
      RECT 386.500000 552.350000 389.000000 555.650000 ;
      RECT 372.500000 552.350000 373.500000 553.650000 ;
      RECT 357.500000 552.350000 358.500000 553.650000 ;
      RECT 2.020000 552.350000 349.500000 554.935000 ;
      RECT 2.020000 551.835000 358.500000 552.350000 ;
      RECT 1166.500000 551.830000 1183.980000 553.650000 ;
      RECT 1139.000000 551.650000 1158.500000 552.350000 ;
      RECT 372.500000 551.650000 389.000000 552.350000 ;
      RECT 0.000000 551.650000 358.500000 551.835000 ;
      RECT 1166.500000 550.350000 1186.000000 551.830000 ;
      RECT 1157.500000 550.350000 1158.500000 551.650000 ;
      RECT 372.500000 550.350000 373.500000 551.650000 ;
      RECT 357.500000 550.350000 358.500000 551.650000 ;
      RECT 1157.500000 549.650000 1186.000000 550.350000 ;
      RECT 357.500000 549.650000 373.500000 550.350000 ;
      RECT 1157.500000 548.350000 1158.500000 549.650000 ;
      RECT 1139.000000 548.350000 1149.500000 551.650000 ;
      RECT 386.500000 548.350000 389.000000 551.650000 ;
      RECT 372.500000 548.350000 373.500000 549.650000 ;
      RECT 357.500000 548.350000 358.500000 549.650000 ;
      RECT 0.000000 548.350000 349.500000 551.650000 ;
      RECT 1139.000000 547.650000 1158.500000 548.350000 ;
      RECT 372.500000 547.650000 389.000000 548.350000 ;
      RECT 0.000000 547.650000 358.500000 548.350000 ;
      RECT 1166.500000 546.350000 1186.000000 549.650000 ;
      RECT 1157.500000 546.350000 1158.500000 547.650000 ;
      RECT 372.500000 546.350000 373.500000 547.650000 ;
      RECT 357.500000 546.350000 358.500000 547.650000 ;
      RECT 1157.500000 545.650000 1186.000000 546.350000 ;
      RECT 357.500000 545.650000 373.500000 546.350000 ;
      RECT 1157.500000 544.350000 1158.500000 545.650000 ;
      RECT 1139.000000 544.350000 1149.500000 547.650000 ;
      RECT 386.500000 544.350000 389.000000 547.650000 ;
      RECT 372.500000 544.350000 373.500000 545.650000 ;
      RECT 357.500000 544.350000 358.500000 545.650000 ;
      RECT 0.000000 544.350000 349.500000 547.650000 ;
      RECT 1139.000000 543.650000 1158.500000 544.350000 ;
      RECT 372.500000 543.650000 389.000000 544.350000 ;
      RECT 0.000000 543.650000 358.500000 544.350000 ;
      RECT 1166.500000 542.350000 1186.000000 545.650000 ;
      RECT 1157.500000 542.350000 1158.500000 543.650000 ;
      RECT 372.500000 542.350000 373.500000 543.650000 ;
      RECT 357.500000 542.350000 358.500000 543.650000 ;
      RECT 1157.500000 541.650000 1186.000000 542.350000 ;
      RECT 357.500000 541.650000 373.500000 542.350000 ;
      RECT 1157.500000 540.350000 1158.500000 541.650000 ;
      RECT 1139.000000 540.350000 1149.500000 543.650000 ;
      RECT 386.500000 540.350000 389.000000 543.650000 ;
      RECT 372.500000 540.350000 373.500000 541.650000 ;
      RECT 357.500000 540.350000 358.500000 541.650000 ;
      RECT 0.000000 540.350000 349.500000 543.650000 ;
      RECT 1139.000000 539.650000 1158.500000 540.350000 ;
      RECT 372.500000 539.650000 389.000000 540.350000 ;
      RECT 0.000000 539.650000 358.500000 540.350000 ;
      RECT 1166.500000 538.350000 1186.000000 541.650000 ;
      RECT 1157.500000 538.350000 1158.500000 539.650000 ;
      RECT 372.500000 538.350000 373.500000 539.650000 ;
      RECT 357.500000 538.350000 358.500000 539.650000 ;
      RECT 1157.500000 537.650000 1186.000000 538.350000 ;
      RECT 357.500000 537.650000 373.500000 538.350000 ;
      RECT 1157.500000 536.350000 1158.500000 537.650000 ;
      RECT 1139.000000 536.350000 1149.500000 539.650000 ;
      RECT 386.500000 536.350000 389.000000 539.650000 ;
      RECT 372.500000 536.350000 373.500000 537.650000 ;
      RECT 357.500000 536.350000 358.500000 537.650000 ;
      RECT 0.000000 536.350000 349.500000 539.650000 ;
      RECT 1139.000000 535.650000 1158.500000 536.350000 ;
      RECT 372.500000 535.650000 389.000000 536.350000 ;
      RECT 0.000000 535.650000 358.500000 536.350000 ;
      RECT 1166.500000 534.350000 1186.000000 537.650000 ;
      RECT 1157.500000 534.350000 1158.500000 535.650000 ;
      RECT 372.500000 534.350000 373.500000 535.650000 ;
      RECT 357.500000 534.350000 358.500000 535.650000 ;
      RECT 1157.500000 533.650000 1186.000000 534.350000 ;
      RECT 357.500000 533.650000 373.500000 534.350000 ;
      RECT 1157.500000 532.350000 1158.500000 533.650000 ;
      RECT 1139.000000 532.350000 1149.500000 535.650000 ;
      RECT 386.500000 532.350000 389.000000 535.650000 ;
      RECT 372.500000 532.350000 373.500000 533.650000 ;
      RECT 357.500000 532.350000 358.500000 533.650000 ;
      RECT 0.000000 532.350000 349.500000 535.650000 ;
      RECT 1139.000000 531.650000 1158.500000 532.350000 ;
      RECT 372.500000 531.650000 389.000000 532.350000 ;
      RECT 0.000000 531.650000 358.500000 532.350000 ;
      RECT 1166.500000 530.350000 1186.000000 533.650000 ;
      RECT 1157.500000 530.350000 1158.500000 531.650000 ;
      RECT 372.500000 530.350000 373.500000 531.650000 ;
      RECT 357.500000 530.350000 358.500000 531.650000 ;
      RECT 1157.500000 529.650000 1186.000000 530.350000 ;
      RECT 357.500000 529.650000 373.500000 530.350000 ;
      RECT 1157.500000 528.350000 1158.500000 529.650000 ;
      RECT 1139.000000 528.350000 1149.500000 531.650000 ;
      RECT 386.500000 528.350000 389.000000 531.650000 ;
      RECT 372.500000 528.350000 373.500000 529.650000 ;
      RECT 357.500000 528.350000 358.500000 529.650000 ;
      RECT 0.000000 528.350000 349.500000 531.650000 ;
      RECT 1139.000000 527.650000 1158.500000 528.350000 ;
      RECT 372.500000 527.650000 389.000000 528.350000 ;
      RECT 0.000000 527.650000 358.500000 528.350000 ;
      RECT 1166.500000 526.350000 1186.000000 529.650000 ;
      RECT 1157.500000 526.350000 1158.500000 527.650000 ;
      RECT 372.500000 526.350000 373.500000 527.650000 ;
      RECT 357.500000 526.350000 358.500000 527.650000 ;
      RECT 1157.500000 525.650000 1186.000000 526.350000 ;
      RECT 357.500000 525.650000 373.500000 526.350000 ;
      RECT 1157.500000 524.350000 1158.500000 525.650000 ;
      RECT 1139.000000 524.350000 1149.500000 527.650000 ;
      RECT 386.500000 524.350000 389.000000 527.650000 ;
      RECT 372.500000 524.350000 373.500000 525.650000 ;
      RECT 357.500000 524.350000 358.500000 525.650000 ;
      RECT 0.000000 524.350000 349.500000 527.650000 ;
      RECT 1139.000000 523.650000 1158.500000 524.350000 ;
      RECT 372.500000 523.650000 389.000000 524.350000 ;
      RECT 0.000000 523.650000 358.500000 524.350000 ;
      RECT 1166.500000 522.350000 1186.000000 525.650000 ;
      RECT 1157.500000 522.350000 1158.500000 523.650000 ;
      RECT 372.500000 522.350000 373.500000 523.650000 ;
      RECT 357.500000 522.350000 358.500000 523.650000 ;
      RECT 1157.500000 521.650000 1186.000000 522.350000 ;
      RECT 357.500000 521.650000 373.500000 522.350000 ;
      RECT 1157.500000 520.350000 1158.500000 521.650000 ;
      RECT 1139.000000 520.350000 1149.500000 523.650000 ;
      RECT 386.500000 520.350000 389.000000 523.650000 ;
      RECT 372.500000 520.350000 373.500000 521.650000 ;
      RECT 357.500000 520.350000 358.500000 521.650000 ;
      RECT 0.000000 520.350000 349.500000 523.650000 ;
      RECT 1139.000000 519.650000 1158.500000 520.350000 ;
      RECT 372.500000 519.650000 389.000000 520.350000 ;
      RECT 0.000000 519.650000 358.500000 520.350000 ;
      RECT 1166.500000 518.350000 1186.000000 521.650000 ;
      RECT 1157.500000 518.350000 1158.500000 519.650000 ;
      RECT 372.500000 518.350000 373.500000 519.650000 ;
      RECT 357.500000 518.350000 358.500000 519.650000 ;
      RECT 1157.500000 517.650000 1186.000000 518.350000 ;
      RECT 357.500000 517.650000 373.500000 518.350000 ;
      RECT 307.500000 517.650000 349.500000 519.650000 ;
      RECT 0.000000 517.650000 299.500000 519.650000 ;
      RECT 1157.500000 516.350000 1158.500000 517.650000 ;
      RECT 1139.000000 516.350000 1149.500000 519.650000 ;
      RECT 386.500000 516.350000 389.000000 519.650000 ;
      RECT 372.500000 516.350000 373.500000 517.650000 ;
      RECT 357.500000 516.350000 358.500000 517.650000 ;
      RECT 316.500000 516.350000 349.500000 517.650000 ;
      RECT 307.500000 516.350000 308.500000 517.650000 ;
      RECT 266.500000 516.350000 299.500000 517.650000 ;
      RECT 1139.000000 515.650000 1158.500000 516.350000 ;
      RECT 372.500000 515.650000 389.000000 516.350000 ;
      RECT 316.500000 515.650000 358.500000 516.350000 ;
      RECT 266.500000 515.650000 308.500000 516.350000 ;
      RECT 216.500000 515.650000 258.500000 517.650000 ;
      RECT 166.500000 515.650000 208.500000 517.650000 ;
      RECT 116.500000 515.650000 158.500000 517.650000 ;
      RECT 66.500000 515.650000 108.500000 517.650000 ;
      RECT 29.500000 515.650000 58.500000 517.650000 ;
      RECT 0.000000 515.650000 16.500000 517.650000 ;
      RECT 1166.500000 514.350000 1186.000000 517.650000 ;
      RECT 1157.500000 514.350000 1158.500000 515.650000 ;
      RECT 372.500000 514.350000 373.500000 515.650000 ;
      RECT 357.500000 514.350000 358.500000 515.650000 ;
      RECT 316.500000 514.350000 349.500000 515.650000 ;
      RECT 307.500000 514.350000 308.500000 515.650000 ;
      RECT 266.500000 514.350000 299.500000 515.650000 ;
      RECT 257.500000 514.350000 258.500000 515.650000 ;
      RECT 216.500000 514.350000 249.500000 515.650000 ;
      RECT 207.500000 514.350000 208.500000 515.650000 ;
      RECT 166.500000 514.350000 199.500000 515.650000 ;
      RECT 157.500000 514.350000 158.500000 515.650000 ;
      RECT 116.500000 514.350000 149.500000 515.650000 ;
      RECT 107.500000 514.350000 108.500000 515.650000 ;
      RECT 66.500000 514.350000 99.500000 515.650000 ;
      RECT 57.500000 514.350000 58.500000 515.650000 ;
      RECT 29.500000 514.350000 49.500000 515.650000 ;
      RECT 15.500000 514.350000 16.500000 515.650000 ;
      RECT 1157.500000 513.650000 1186.000000 514.350000 ;
      RECT 357.500000 513.650000 373.500000 514.350000 ;
      RECT 307.500000 513.650000 349.500000 514.350000 ;
      RECT 257.500000 513.650000 299.500000 514.350000 ;
      RECT 207.500000 513.650000 249.500000 514.350000 ;
      RECT 157.500000 513.650000 199.500000 514.350000 ;
      RECT 107.500000 513.650000 149.500000 514.350000 ;
      RECT 57.500000 513.650000 99.500000 514.350000 ;
      RECT 15.500000 513.650000 49.500000 514.350000 ;
      RECT 1157.500000 512.350000 1158.500000 513.650000 ;
      RECT 1139.000000 512.350000 1149.500000 515.650000 ;
      RECT 386.500000 512.350000 389.000000 515.650000 ;
      RECT 372.500000 512.350000 373.500000 513.650000 ;
      RECT 357.500000 512.350000 358.500000 513.650000 ;
      RECT 316.500000 512.350000 349.500000 513.650000 ;
      RECT 307.500000 512.350000 308.500000 513.650000 ;
      RECT 266.500000 512.350000 299.500000 513.650000 ;
      RECT 257.500000 512.350000 258.500000 513.650000 ;
      RECT 216.500000 512.350000 249.500000 513.650000 ;
      RECT 207.500000 512.350000 208.500000 513.650000 ;
      RECT 166.500000 512.350000 199.500000 513.650000 ;
      RECT 157.500000 512.350000 158.500000 513.650000 ;
      RECT 116.500000 512.350000 149.500000 513.650000 ;
      RECT 107.500000 512.350000 108.500000 513.650000 ;
      RECT 66.500000 512.350000 99.500000 513.650000 ;
      RECT 57.500000 512.350000 58.500000 513.650000 ;
      RECT 29.500000 512.350000 49.500000 513.650000 ;
      RECT 15.500000 512.350000 16.500000 513.650000 ;
      RECT 0.000000 512.350000 2.500000 515.650000 ;
      RECT 1139.000000 511.650000 1158.500000 512.350000 ;
      RECT 372.500000 511.650000 389.000000 512.350000 ;
      RECT 316.500000 511.650000 358.500000 512.350000 ;
      RECT 266.500000 511.650000 308.500000 512.350000 ;
      RECT 216.500000 511.650000 258.500000 512.350000 ;
      RECT 166.500000 511.650000 208.500000 512.350000 ;
      RECT 116.500000 511.650000 158.500000 512.350000 ;
      RECT 66.500000 511.650000 108.500000 512.350000 ;
      RECT 29.500000 511.650000 58.500000 512.350000 ;
      RECT 0.000000 511.650000 16.500000 512.350000 ;
      RECT 1166.500000 510.350000 1186.000000 513.650000 ;
      RECT 1157.500000 510.350000 1158.500000 511.650000 ;
      RECT 372.500000 510.350000 373.500000 511.650000 ;
      RECT 357.500000 510.350000 358.500000 511.650000 ;
      RECT 316.500000 510.350000 349.500000 511.650000 ;
      RECT 307.500000 510.350000 308.500000 511.650000 ;
      RECT 266.500000 510.350000 299.500000 511.650000 ;
      RECT 257.500000 510.350000 258.500000 511.650000 ;
      RECT 216.500000 510.350000 249.500000 511.650000 ;
      RECT 207.500000 510.350000 208.500000 511.650000 ;
      RECT 166.500000 510.350000 199.500000 511.650000 ;
      RECT 157.500000 510.350000 158.500000 511.650000 ;
      RECT 116.500000 510.350000 149.500000 511.650000 ;
      RECT 107.500000 510.350000 108.500000 511.650000 ;
      RECT 66.500000 510.350000 99.500000 511.650000 ;
      RECT 57.500000 510.350000 58.500000 511.650000 ;
      RECT 29.500000 510.350000 49.500000 511.650000 ;
      RECT 15.500000 510.350000 16.500000 511.650000 ;
      RECT 1157.500000 509.650000 1186.000000 510.350000 ;
      RECT 357.500000 509.650000 373.500000 510.350000 ;
      RECT 307.500000 509.650000 349.500000 510.350000 ;
      RECT 257.500000 509.650000 299.500000 510.350000 ;
      RECT 207.500000 509.650000 249.500000 510.350000 ;
      RECT 157.500000 509.650000 199.500000 510.350000 ;
      RECT 107.500000 509.650000 149.500000 510.350000 ;
      RECT 57.500000 509.650000 99.500000 510.350000 ;
      RECT 15.500000 509.650000 49.500000 510.350000 ;
      RECT 1157.500000 508.350000 1158.500000 509.650000 ;
      RECT 1139.000000 508.350000 1149.500000 511.650000 ;
      RECT 386.500000 508.350000 389.000000 511.650000 ;
      RECT 372.500000 508.350000 373.500000 509.650000 ;
      RECT 357.500000 508.350000 358.500000 509.650000 ;
      RECT 316.500000 508.350000 349.500000 509.650000 ;
      RECT 307.500000 508.350000 308.500000 509.650000 ;
      RECT 266.500000 508.350000 299.500000 509.650000 ;
      RECT 257.500000 508.350000 258.500000 509.650000 ;
      RECT 216.500000 508.350000 249.500000 509.650000 ;
      RECT 207.500000 508.350000 208.500000 509.650000 ;
      RECT 166.500000 508.350000 199.500000 509.650000 ;
      RECT 157.500000 508.350000 158.500000 509.650000 ;
      RECT 116.500000 508.350000 149.500000 509.650000 ;
      RECT 107.500000 508.350000 108.500000 509.650000 ;
      RECT 66.500000 508.350000 99.500000 509.650000 ;
      RECT 57.500000 508.350000 58.500000 509.650000 ;
      RECT 29.500000 508.350000 49.500000 509.650000 ;
      RECT 15.500000 508.350000 16.500000 509.650000 ;
      RECT 0.000000 508.350000 2.500000 511.650000 ;
      RECT 1139.000000 507.650000 1158.500000 508.350000 ;
      RECT 372.500000 507.650000 389.000000 508.350000 ;
      RECT 316.500000 507.650000 358.500000 508.350000 ;
      RECT 266.500000 507.650000 308.500000 508.350000 ;
      RECT 216.500000 507.650000 258.500000 508.350000 ;
      RECT 166.500000 507.650000 208.500000 508.350000 ;
      RECT 116.500000 507.650000 158.500000 508.350000 ;
      RECT 66.500000 507.650000 108.500000 508.350000 ;
      RECT 29.500000 507.650000 58.500000 508.350000 ;
      RECT 0.000000 507.650000 16.500000 508.350000 ;
      RECT 1166.500000 506.350000 1186.000000 509.650000 ;
      RECT 1157.500000 506.350000 1158.500000 507.650000 ;
      RECT 372.500000 506.350000 373.500000 507.650000 ;
      RECT 357.500000 506.350000 358.500000 507.650000 ;
      RECT 316.500000 506.350000 349.500000 507.650000 ;
      RECT 307.500000 506.350000 308.500000 507.650000 ;
      RECT 266.500000 506.350000 299.500000 507.650000 ;
      RECT 257.500000 506.350000 258.500000 507.650000 ;
      RECT 216.500000 506.350000 249.500000 507.650000 ;
      RECT 207.500000 506.350000 208.500000 507.650000 ;
      RECT 166.500000 506.350000 199.500000 507.650000 ;
      RECT 157.500000 506.350000 158.500000 507.650000 ;
      RECT 116.500000 506.350000 149.500000 507.650000 ;
      RECT 107.500000 506.350000 108.500000 507.650000 ;
      RECT 66.500000 506.350000 99.500000 507.650000 ;
      RECT 57.500000 506.350000 58.500000 507.650000 ;
      RECT 29.500000 506.350000 49.500000 507.650000 ;
      RECT 15.500000 506.350000 16.500000 507.650000 ;
      RECT 386.500000 506.000000 389.000000 507.650000 ;
      RECT 1157.500000 505.650000 1186.000000 506.350000 ;
      RECT 386.500000 505.650000 739.000000 506.000000 ;
      RECT 357.500000 505.650000 373.500000 506.350000 ;
      RECT 307.500000 505.650000 349.500000 506.350000 ;
      RECT 257.500000 505.650000 299.500000 506.350000 ;
      RECT 207.500000 505.650000 249.500000 506.350000 ;
      RECT 157.500000 505.650000 199.500000 506.350000 ;
      RECT 107.500000 505.650000 149.500000 506.350000 ;
      RECT 57.500000 505.650000 99.500000 506.350000 ;
      RECT 15.500000 505.650000 49.500000 506.350000 ;
      RECT 1157.500000 504.350000 1158.500000 505.650000 ;
      RECT 1139.000000 504.350000 1149.500000 507.650000 ;
      RECT 386.500000 504.350000 408.500000 505.650000 ;
      RECT 372.500000 504.350000 373.500000 505.650000 ;
      RECT 357.500000 504.350000 358.500000 505.650000 ;
      RECT 316.500000 504.350000 349.500000 505.650000 ;
      RECT 307.500000 504.350000 308.500000 505.650000 ;
      RECT 266.500000 504.350000 299.500000 505.650000 ;
      RECT 257.500000 504.350000 258.500000 505.650000 ;
      RECT 216.500000 504.350000 249.500000 505.650000 ;
      RECT 207.500000 504.350000 208.500000 505.650000 ;
      RECT 166.500000 504.350000 199.500000 505.650000 ;
      RECT 157.500000 504.350000 158.500000 505.650000 ;
      RECT 116.500000 504.350000 149.500000 505.650000 ;
      RECT 107.500000 504.350000 108.500000 505.650000 ;
      RECT 66.500000 504.350000 99.500000 505.650000 ;
      RECT 57.500000 504.350000 58.500000 505.650000 ;
      RECT 29.500000 504.350000 49.500000 505.650000 ;
      RECT 15.500000 504.350000 16.500000 505.650000 ;
      RECT 0.000000 504.350000 2.500000 507.650000 ;
      RECT 1139.000000 503.650000 1158.500000 504.350000 ;
      RECT 716.500000 503.650000 739.000000 505.650000 ;
      RECT 666.500000 503.650000 708.500000 505.650000 ;
      RECT 616.500000 503.650000 658.500000 505.650000 ;
      RECT 566.500000 503.650000 608.500000 505.650000 ;
      RECT 516.500000 503.650000 558.500000 505.650000 ;
      RECT 466.500000 503.650000 508.500000 505.650000 ;
      RECT 416.500000 503.650000 458.500000 505.650000 ;
      RECT 372.500000 503.650000 408.500000 504.350000 ;
      RECT 316.500000 503.650000 358.500000 504.350000 ;
      RECT 266.500000 503.650000 308.500000 504.350000 ;
      RECT 216.500000 503.650000 258.500000 504.350000 ;
      RECT 166.500000 503.650000 208.500000 504.350000 ;
      RECT 116.500000 503.650000 158.500000 504.350000 ;
      RECT 66.500000 503.650000 108.500000 504.350000 ;
      RECT 29.500000 503.650000 58.500000 504.350000 ;
      RECT 0.000000 503.650000 16.500000 504.350000 ;
      RECT 1166.500000 502.350000 1186.000000 505.650000 ;
      RECT 1157.500000 502.350000 1158.500000 503.650000 ;
      RECT 716.500000 502.350000 723.500000 503.650000 ;
      RECT 707.500000 502.350000 708.500000 503.650000 ;
      RECT 666.500000 502.350000 699.500000 503.650000 ;
      RECT 657.500000 502.350000 658.500000 503.650000 ;
      RECT 616.500000 502.350000 649.500000 503.650000 ;
      RECT 607.500000 502.350000 608.500000 503.650000 ;
      RECT 566.500000 502.350000 599.500000 503.650000 ;
      RECT 557.500000 502.350000 558.500000 503.650000 ;
      RECT 516.500000 502.350000 549.500000 503.650000 ;
      RECT 507.500000 502.350000 508.500000 503.650000 ;
      RECT 466.500000 502.350000 499.500000 503.650000 ;
      RECT 457.500000 502.350000 458.500000 503.650000 ;
      RECT 416.500000 502.350000 449.500000 503.650000 ;
      RECT 407.500000 502.350000 408.500000 503.650000 ;
      RECT 372.500000 502.350000 373.500000 503.650000 ;
      RECT 357.500000 502.350000 358.500000 503.650000 ;
      RECT 316.500000 502.350000 349.500000 503.650000 ;
      RECT 307.500000 502.350000 308.500000 503.650000 ;
      RECT 266.500000 502.350000 299.500000 503.650000 ;
      RECT 257.500000 502.350000 258.500000 503.650000 ;
      RECT 216.500000 502.350000 249.500000 503.650000 ;
      RECT 207.500000 502.350000 208.500000 503.650000 ;
      RECT 166.500000 502.350000 199.500000 503.650000 ;
      RECT 157.500000 502.350000 158.500000 503.650000 ;
      RECT 116.500000 502.350000 149.500000 503.650000 ;
      RECT 107.500000 502.350000 108.500000 503.650000 ;
      RECT 66.500000 502.350000 99.500000 503.650000 ;
      RECT 57.500000 502.350000 58.500000 503.650000 ;
      RECT 29.500000 502.350000 49.500000 503.650000 ;
      RECT 15.500000 502.350000 16.500000 503.650000 ;
      RECT 1157.500000 501.650000 1186.000000 502.350000 ;
      RECT 707.500000 501.650000 723.500000 502.350000 ;
      RECT 657.500000 501.650000 699.500000 502.350000 ;
      RECT 607.500000 501.650000 649.500000 502.350000 ;
      RECT 557.500000 501.650000 599.500000 502.350000 ;
      RECT 507.500000 501.650000 549.500000 502.350000 ;
      RECT 457.500000 501.650000 499.500000 502.350000 ;
      RECT 407.500000 501.650000 449.500000 502.350000 ;
      RECT 357.500000 501.650000 373.500000 502.350000 ;
      RECT 307.500000 501.650000 349.500000 502.350000 ;
      RECT 257.500000 501.650000 299.500000 502.350000 ;
      RECT 207.500000 501.650000 249.500000 502.350000 ;
      RECT 157.500000 501.650000 199.500000 502.350000 ;
      RECT 107.500000 501.650000 149.500000 502.350000 ;
      RECT 57.500000 501.650000 99.500000 502.350000 ;
      RECT 15.500000 501.650000 49.500000 502.350000 ;
      RECT 1157.500000 500.350000 1158.500000 501.650000 ;
      RECT 1139.000000 500.350000 1149.500000 503.650000 ;
      RECT 736.500000 500.350000 739.000000 503.650000 ;
      RECT 716.500000 500.350000 723.500000 501.650000 ;
      RECT 707.500000 500.350000 708.500000 501.650000 ;
      RECT 666.500000 500.350000 699.500000 501.650000 ;
      RECT 657.500000 500.350000 658.500000 501.650000 ;
      RECT 616.500000 500.350000 649.500000 501.650000 ;
      RECT 607.500000 500.350000 608.500000 501.650000 ;
      RECT 566.500000 500.350000 599.500000 501.650000 ;
      RECT 557.500000 500.350000 558.500000 501.650000 ;
      RECT 516.500000 500.350000 549.500000 501.650000 ;
      RECT 507.500000 500.350000 508.500000 501.650000 ;
      RECT 466.500000 500.350000 499.500000 501.650000 ;
      RECT 457.500000 500.350000 458.500000 501.650000 ;
      RECT 416.500000 500.350000 449.500000 501.650000 ;
      RECT 407.500000 500.350000 408.500000 501.650000 ;
      RECT 386.500000 500.350000 399.500000 503.650000 ;
      RECT 372.500000 500.350000 373.500000 501.650000 ;
      RECT 357.500000 500.350000 358.500000 501.650000 ;
      RECT 316.500000 500.350000 349.500000 501.650000 ;
      RECT 307.500000 500.350000 308.500000 501.650000 ;
      RECT 266.500000 500.350000 299.500000 501.650000 ;
      RECT 257.500000 500.350000 258.500000 501.650000 ;
      RECT 216.500000 500.350000 249.500000 501.650000 ;
      RECT 207.500000 500.350000 208.500000 501.650000 ;
      RECT 166.500000 500.350000 199.500000 501.650000 ;
      RECT 157.500000 500.350000 158.500000 501.650000 ;
      RECT 116.500000 500.350000 149.500000 501.650000 ;
      RECT 107.500000 500.350000 108.500000 501.650000 ;
      RECT 66.500000 500.350000 99.500000 501.650000 ;
      RECT 57.500000 500.350000 58.500000 501.650000 ;
      RECT 29.500000 500.350000 49.500000 501.650000 ;
      RECT 15.500000 500.350000 16.500000 501.650000 ;
      RECT 0.000000 500.350000 2.500000 503.650000 ;
      RECT 1139.000000 499.650000 1158.500000 500.350000 ;
      RECT 716.500000 499.650000 739.000000 500.350000 ;
      RECT 666.500000 499.650000 708.500000 500.350000 ;
      RECT 616.500000 499.650000 658.500000 500.350000 ;
      RECT 566.500000 499.650000 608.500000 500.350000 ;
      RECT 516.500000 499.650000 558.500000 500.350000 ;
      RECT 466.500000 499.650000 508.500000 500.350000 ;
      RECT 416.500000 499.650000 458.500000 500.350000 ;
      RECT 372.500000 499.650000 408.500000 500.350000 ;
      RECT 316.500000 499.650000 358.500000 500.350000 ;
      RECT 266.500000 499.650000 308.500000 500.350000 ;
      RECT 216.500000 499.650000 258.500000 500.350000 ;
      RECT 166.500000 499.650000 208.500000 500.350000 ;
      RECT 116.500000 499.650000 158.500000 500.350000 ;
      RECT 66.500000 499.650000 108.500000 500.350000 ;
      RECT 29.500000 499.650000 58.500000 500.350000 ;
      RECT 0.000000 499.650000 16.500000 500.350000 ;
      RECT 1166.500000 498.350000 1186.000000 501.650000 ;
      RECT 1157.500000 498.350000 1158.500000 499.650000 ;
      RECT 716.500000 498.350000 723.500000 499.650000 ;
      RECT 707.500000 498.350000 708.500000 499.650000 ;
      RECT 666.500000 498.350000 699.500000 499.650000 ;
      RECT 657.500000 498.350000 658.500000 499.650000 ;
      RECT 616.500000 498.350000 649.500000 499.650000 ;
      RECT 607.500000 498.350000 608.500000 499.650000 ;
      RECT 566.500000 498.350000 599.500000 499.650000 ;
      RECT 557.500000 498.350000 558.500000 499.650000 ;
      RECT 516.500000 498.350000 549.500000 499.650000 ;
      RECT 507.500000 498.350000 508.500000 499.650000 ;
      RECT 466.500000 498.350000 499.500000 499.650000 ;
      RECT 457.500000 498.350000 458.500000 499.650000 ;
      RECT 416.500000 498.350000 449.500000 499.650000 ;
      RECT 407.500000 498.350000 408.500000 499.650000 ;
      RECT 372.500000 498.350000 373.500000 499.650000 ;
      RECT 357.500000 498.350000 358.500000 499.650000 ;
      RECT 316.500000 498.350000 349.500000 499.650000 ;
      RECT 307.500000 498.350000 308.500000 499.650000 ;
      RECT 266.500000 498.350000 299.500000 499.650000 ;
      RECT 257.500000 498.350000 258.500000 499.650000 ;
      RECT 216.500000 498.350000 249.500000 499.650000 ;
      RECT 207.500000 498.350000 208.500000 499.650000 ;
      RECT 166.500000 498.350000 199.500000 499.650000 ;
      RECT 157.500000 498.350000 158.500000 499.650000 ;
      RECT 116.500000 498.350000 149.500000 499.650000 ;
      RECT 107.500000 498.350000 108.500000 499.650000 ;
      RECT 66.500000 498.350000 99.500000 499.650000 ;
      RECT 57.500000 498.350000 58.500000 499.650000 ;
      RECT 29.500000 498.350000 49.500000 499.650000 ;
      RECT 15.500000 498.350000 16.500000 499.650000 ;
      RECT 1157.500000 497.650000 1186.000000 498.350000 ;
      RECT 707.500000 497.650000 723.500000 498.350000 ;
      RECT 657.500000 497.650000 699.500000 498.350000 ;
      RECT 607.500000 497.650000 649.500000 498.350000 ;
      RECT 557.500000 497.650000 599.500000 498.350000 ;
      RECT 507.500000 497.650000 549.500000 498.350000 ;
      RECT 457.500000 497.650000 499.500000 498.350000 ;
      RECT 407.500000 497.650000 449.500000 498.350000 ;
      RECT 357.500000 497.650000 373.500000 498.350000 ;
      RECT 307.500000 497.650000 349.500000 498.350000 ;
      RECT 257.500000 497.650000 299.500000 498.350000 ;
      RECT 207.500000 497.650000 249.500000 498.350000 ;
      RECT 157.500000 497.650000 199.500000 498.350000 ;
      RECT 107.500000 497.650000 149.500000 498.350000 ;
      RECT 57.500000 497.650000 99.500000 498.350000 ;
      RECT 15.500000 497.650000 49.500000 498.350000 ;
      RECT 1157.500000 496.350000 1158.500000 497.650000 ;
      RECT 1139.000000 496.350000 1149.500000 499.650000 ;
      RECT 736.500000 496.350000 739.000000 499.650000 ;
      RECT 716.500000 496.350000 723.500000 497.650000 ;
      RECT 707.500000 496.350000 708.500000 497.650000 ;
      RECT 666.500000 496.350000 699.500000 497.650000 ;
      RECT 657.500000 496.350000 658.500000 497.650000 ;
      RECT 616.500000 496.350000 649.500000 497.650000 ;
      RECT 607.500000 496.350000 608.500000 497.650000 ;
      RECT 566.500000 496.350000 599.500000 497.650000 ;
      RECT 557.500000 496.350000 558.500000 497.650000 ;
      RECT 516.500000 496.350000 549.500000 497.650000 ;
      RECT 507.500000 496.350000 508.500000 497.650000 ;
      RECT 466.500000 496.350000 499.500000 497.650000 ;
      RECT 457.500000 496.350000 458.500000 497.650000 ;
      RECT 416.500000 496.350000 449.500000 497.650000 ;
      RECT 407.500000 496.350000 408.500000 497.650000 ;
      RECT 386.500000 496.350000 399.500000 499.650000 ;
      RECT 372.500000 496.350000 373.500000 497.650000 ;
      RECT 357.500000 496.350000 358.500000 497.650000 ;
      RECT 316.500000 496.350000 349.500000 497.650000 ;
      RECT 307.500000 496.350000 308.500000 497.650000 ;
      RECT 266.500000 496.350000 299.500000 497.650000 ;
      RECT 257.500000 496.350000 258.500000 497.650000 ;
      RECT 216.500000 496.350000 249.500000 497.650000 ;
      RECT 207.500000 496.350000 208.500000 497.650000 ;
      RECT 166.500000 496.350000 199.500000 497.650000 ;
      RECT 157.500000 496.350000 158.500000 497.650000 ;
      RECT 116.500000 496.350000 149.500000 497.650000 ;
      RECT 107.500000 496.350000 108.500000 497.650000 ;
      RECT 66.500000 496.350000 99.500000 497.650000 ;
      RECT 57.500000 496.350000 58.500000 497.650000 ;
      RECT 29.500000 496.350000 49.500000 497.650000 ;
      RECT 15.500000 496.350000 16.500000 497.650000 ;
      RECT 0.000000 496.350000 2.500000 499.650000 ;
      RECT 1139.000000 495.650000 1158.500000 496.350000 ;
      RECT 716.500000 495.650000 739.000000 496.350000 ;
      RECT 666.500000 495.650000 708.500000 496.350000 ;
      RECT 616.500000 495.650000 658.500000 496.350000 ;
      RECT 566.500000 495.650000 608.500000 496.350000 ;
      RECT 516.500000 495.650000 558.500000 496.350000 ;
      RECT 466.500000 495.650000 508.500000 496.350000 ;
      RECT 416.500000 495.650000 458.500000 496.350000 ;
      RECT 372.500000 495.650000 408.500000 496.350000 ;
      RECT 316.500000 495.650000 358.500000 496.350000 ;
      RECT 266.500000 495.650000 308.500000 496.350000 ;
      RECT 216.500000 495.650000 258.500000 496.350000 ;
      RECT 166.500000 495.650000 208.500000 496.350000 ;
      RECT 116.500000 495.650000 158.500000 496.350000 ;
      RECT 66.500000 495.650000 108.500000 496.350000 ;
      RECT 29.500000 495.650000 58.500000 496.350000 ;
      RECT 0.000000 495.650000 16.500000 496.350000 ;
      RECT 1166.500000 494.350000 1186.000000 497.650000 ;
      RECT 1157.500000 494.350000 1158.500000 495.650000 ;
      RECT 716.500000 494.350000 723.500000 495.650000 ;
      RECT 707.500000 494.350000 708.500000 495.650000 ;
      RECT 666.500000 494.350000 699.500000 495.650000 ;
      RECT 657.500000 494.350000 658.500000 495.650000 ;
      RECT 616.500000 494.350000 649.500000 495.650000 ;
      RECT 607.500000 494.350000 608.500000 495.650000 ;
      RECT 566.500000 494.350000 599.500000 495.650000 ;
      RECT 557.500000 494.350000 558.500000 495.650000 ;
      RECT 516.500000 494.350000 549.500000 495.650000 ;
      RECT 507.500000 494.350000 508.500000 495.650000 ;
      RECT 466.500000 494.350000 499.500000 495.650000 ;
      RECT 457.500000 494.350000 458.500000 495.650000 ;
      RECT 416.500000 494.350000 449.500000 495.650000 ;
      RECT 407.500000 494.350000 408.500000 495.650000 ;
      RECT 372.500000 494.350000 373.500000 495.650000 ;
      RECT 357.500000 494.350000 358.500000 495.650000 ;
      RECT 316.500000 494.350000 349.500000 495.650000 ;
      RECT 307.500000 494.350000 308.500000 495.650000 ;
      RECT 266.500000 494.350000 299.500000 495.650000 ;
      RECT 257.500000 494.350000 258.500000 495.650000 ;
      RECT 216.500000 494.350000 249.500000 495.650000 ;
      RECT 207.500000 494.350000 208.500000 495.650000 ;
      RECT 166.500000 494.350000 199.500000 495.650000 ;
      RECT 157.500000 494.350000 158.500000 495.650000 ;
      RECT 116.500000 494.350000 149.500000 495.650000 ;
      RECT 107.500000 494.350000 108.500000 495.650000 ;
      RECT 66.500000 494.350000 99.500000 495.650000 ;
      RECT 57.500000 494.350000 58.500000 495.650000 ;
      RECT 29.500000 494.350000 49.500000 495.650000 ;
      RECT 15.500000 494.350000 16.500000 495.650000 ;
      RECT 1157.500000 493.650000 1186.000000 494.350000 ;
      RECT 707.500000 493.650000 723.500000 494.350000 ;
      RECT 657.500000 493.650000 699.500000 494.350000 ;
      RECT 607.500000 493.650000 649.500000 494.350000 ;
      RECT 557.500000 493.650000 599.500000 494.350000 ;
      RECT 507.500000 493.650000 549.500000 494.350000 ;
      RECT 457.500000 493.650000 499.500000 494.350000 ;
      RECT 407.500000 493.650000 449.500000 494.350000 ;
      RECT 357.500000 493.650000 373.500000 494.350000 ;
      RECT 307.500000 493.650000 349.500000 494.350000 ;
      RECT 257.500000 493.650000 299.500000 494.350000 ;
      RECT 207.500000 493.650000 249.500000 494.350000 ;
      RECT 157.500000 493.650000 199.500000 494.350000 ;
      RECT 107.500000 493.650000 149.500000 494.350000 ;
      RECT 57.500000 493.650000 99.500000 494.350000 ;
      RECT 15.500000 493.650000 49.500000 494.350000 ;
      RECT 1157.500000 492.350000 1158.500000 493.650000 ;
      RECT 1139.000000 492.350000 1149.500000 495.650000 ;
      RECT 736.500000 492.350000 739.000000 495.650000 ;
      RECT 716.500000 492.350000 723.500000 493.650000 ;
      RECT 707.500000 492.350000 708.500000 493.650000 ;
      RECT 666.500000 492.350000 699.500000 493.650000 ;
      RECT 657.500000 492.350000 658.500000 493.650000 ;
      RECT 616.500000 492.350000 649.500000 493.650000 ;
      RECT 607.500000 492.350000 608.500000 493.650000 ;
      RECT 566.500000 492.350000 599.500000 493.650000 ;
      RECT 557.500000 492.350000 558.500000 493.650000 ;
      RECT 516.500000 492.350000 549.500000 493.650000 ;
      RECT 507.500000 492.350000 508.500000 493.650000 ;
      RECT 466.500000 492.350000 499.500000 493.650000 ;
      RECT 457.500000 492.350000 458.500000 493.650000 ;
      RECT 416.500000 492.350000 449.500000 493.650000 ;
      RECT 407.500000 492.350000 408.500000 493.650000 ;
      RECT 386.500000 492.350000 399.500000 495.650000 ;
      RECT 372.500000 492.350000 373.500000 493.650000 ;
      RECT 357.500000 492.350000 358.500000 493.650000 ;
      RECT 316.500000 492.350000 349.500000 493.650000 ;
      RECT 307.500000 492.350000 308.500000 493.650000 ;
      RECT 266.500000 492.350000 299.500000 493.650000 ;
      RECT 257.500000 492.350000 258.500000 493.650000 ;
      RECT 216.500000 492.350000 249.500000 493.650000 ;
      RECT 207.500000 492.350000 208.500000 493.650000 ;
      RECT 166.500000 492.350000 199.500000 493.650000 ;
      RECT 157.500000 492.350000 158.500000 493.650000 ;
      RECT 116.500000 492.350000 149.500000 493.650000 ;
      RECT 107.500000 492.350000 108.500000 493.650000 ;
      RECT 66.500000 492.350000 99.500000 493.650000 ;
      RECT 57.500000 492.350000 58.500000 493.650000 ;
      RECT 29.500000 492.350000 49.500000 493.650000 ;
      RECT 15.500000 492.350000 16.500000 493.650000 ;
      RECT 0.000000 492.350000 2.500000 495.650000 ;
      RECT 1139.000000 491.650000 1158.500000 492.350000 ;
      RECT 716.500000 491.650000 739.000000 492.350000 ;
      RECT 666.500000 491.650000 708.500000 492.350000 ;
      RECT 616.500000 491.650000 658.500000 492.350000 ;
      RECT 566.500000 491.650000 608.500000 492.350000 ;
      RECT 516.500000 491.650000 558.500000 492.350000 ;
      RECT 466.500000 491.650000 508.500000 492.350000 ;
      RECT 416.500000 491.650000 458.500000 492.350000 ;
      RECT 372.500000 491.650000 408.500000 492.350000 ;
      RECT 316.500000 491.650000 358.500000 492.350000 ;
      RECT 266.500000 491.650000 308.500000 492.350000 ;
      RECT 216.500000 491.650000 258.500000 492.350000 ;
      RECT 166.500000 491.650000 208.500000 492.350000 ;
      RECT 116.500000 491.650000 158.500000 492.350000 ;
      RECT 66.500000 491.650000 108.500000 492.350000 ;
      RECT 29.500000 491.650000 58.500000 492.350000 ;
      RECT 0.000000 491.650000 16.500000 492.350000 ;
      RECT 1166.500000 490.350000 1186.000000 493.650000 ;
      RECT 1157.500000 490.350000 1158.500000 491.650000 ;
      RECT 716.500000 490.350000 723.500000 491.650000 ;
      RECT 707.500000 490.350000 708.500000 491.650000 ;
      RECT 666.500000 490.350000 699.500000 491.650000 ;
      RECT 657.500000 490.350000 658.500000 491.650000 ;
      RECT 616.500000 490.350000 649.500000 491.650000 ;
      RECT 607.500000 490.350000 608.500000 491.650000 ;
      RECT 566.500000 490.350000 599.500000 491.650000 ;
      RECT 557.500000 490.350000 558.500000 491.650000 ;
      RECT 516.500000 490.350000 549.500000 491.650000 ;
      RECT 507.500000 490.350000 508.500000 491.650000 ;
      RECT 466.500000 490.350000 499.500000 491.650000 ;
      RECT 457.500000 490.350000 458.500000 491.650000 ;
      RECT 416.500000 490.350000 449.500000 491.650000 ;
      RECT 407.500000 490.350000 408.500000 491.650000 ;
      RECT 372.500000 490.350000 399.500000 491.650000 ;
      RECT 357.500000 490.350000 358.500000 491.650000 ;
      RECT 316.500000 490.350000 349.500000 491.650000 ;
      RECT 307.500000 490.350000 308.500000 491.650000 ;
      RECT 266.500000 490.350000 299.500000 491.650000 ;
      RECT 257.500000 490.350000 258.500000 491.650000 ;
      RECT 216.500000 490.350000 249.500000 491.650000 ;
      RECT 207.500000 490.350000 208.500000 491.650000 ;
      RECT 166.500000 490.350000 199.500000 491.650000 ;
      RECT 157.500000 490.350000 158.500000 491.650000 ;
      RECT 116.500000 490.350000 149.500000 491.650000 ;
      RECT 107.500000 490.350000 108.500000 491.650000 ;
      RECT 66.500000 490.350000 99.500000 491.650000 ;
      RECT 57.500000 490.350000 58.500000 491.650000 ;
      RECT 29.500000 490.350000 49.500000 491.650000 ;
      RECT 15.500000 490.350000 16.500000 491.650000 ;
      RECT 1157.500000 489.650000 1186.000000 490.350000 ;
      RECT 707.500000 489.650000 723.500000 490.350000 ;
      RECT 657.500000 489.650000 699.500000 490.350000 ;
      RECT 607.500000 489.650000 649.500000 490.350000 ;
      RECT 557.500000 489.650000 599.500000 490.350000 ;
      RECT 507.500000 489.650000 549.500000 490.350000 ;
      RECT 457.500000 489.650000 499.500000 490.350000 ;
      RECT 407.500000 489.650000 449.500000 490.350000 ;
      RECT 357.500000 489.650000 399.500000 490.350000 ;
      RECT 307.500000 489.650000 349.500000 490.350000 ;
      RECT 257.500000 489.650000 299.500000 490.350000 ;
      RECT 207.500000 489.650000 249.500000 490.350000 ;
      RECT 157.500000 489.650000 199.500000 490.350000 ;
      RECT 107.500000 489.650000 149.500000 490.350000 ;
      RECT 57.500000 489.650000 99.500000 490.350000 ;
      RECT 15.500000 489.650000 49.500000 490.350000 ;
      RECT 1157.500000 488.350000 1158.500000 489.650000 ;
      RECT 1139.000000 488.350000 1149.500000 491.650000 ;
      RECT 736.500000 488.350000 739.000000 491.650000 ;
      RECT 722.500000 488.350000 723.500000 489.650000 ;
      RECT 707.500000 488.350000 708.500000 489.650000 ;
      RECT 666.500000 488.350000 699.500000 489.650000 ;
      RECT 657.500000 488.350000 658.500000 489.650000 ;
      RECT 616.500000 488.350000 649.500000 489.650000 ;
      RECT 607.500000 488.350000 608.500000 489.650000 ;
      RECT 566.500000 488.350000 599.500000 489.650000 ;
      RECT 557.500000 488.350000 558.500000 489.650000 ;
      RECT 516.500000 488.350000 549.500000 489.650000 ;
      RECT 507.500000 488.350000 508.500000 489.650000 ;
      RECT 466.500000 488.350000 499.500000 489.650000 ;
      RECT 457.500000 488.350000 458.500000 489.650000 ;
      RECT 416.500000 488.350000 449.500000 489.650000 ;
      RECT 407.500000 488.350000 408.500000 489.650000 ;
      RECT 372.500000 488.350000 399.500000 489.650000 ;
      RECT 357.500000 488.350000 359.500000 489.650000 ;
      RECT 316.500000 488.350000 349.500000 489.650000 ;
      RECT 307.500000 488.350000 308.500000 489.650000 ;
      RECT 266.500000 488.350000 299.500000 489.650000 ;
      RECT 257.500000 488.350000 258.500000 489.650000 ;
      RECT 216.500000 488.350000 249.500000 489.650000 ;
      RECT 207.500000 488.350000 208.500000 489.650000 ;
      RECT 166.500000 488.350000 199.500000 489.650000 ;
      RECT 157.500000 488.350000 158.500000 489.650000 ;
      RECT 116.500000 488.350000 149.500000 489.650000 ;
      RECT 107.500000 488.350000 108.500000 489.650000 ;
      RECT 66.500000 488.350000 99.500000 489.650000 ;
      RECT 57.500000 488.350000 58.500000 489.650000 ;
      RECT 29.500000 488.350000 49.500000 489.650000 ;
      RECT 15.500000 488.350000 16.500000 489.650000 ;
      RECT 0.000000 488.350000 2.500000 491.650000 ;
      RECT 1139.000000 487.650000 1158.500000 488.350000 ;
      RECT 722.500000 487.650000 739.000000 488.350000 ;
      RECT 666.500000 487.650000 708.500000 488.350000 ;
      RECT 616.500000 487.650000 658.500000 488.350000 ;
      RECT 566.500000 487.650000 608.500000 488.350000 ;
      RECT 516.500000 487.650000 558.500000 488.350000 ;
      RECT 466.500000 487.650000 508.500000 488.350000 ;
      RECT 416.500000 487.650000 458.500000 488.350000 ;
      RECT 372.500000 487.650000 408.500000 488.350000 ;
      RECT 316.500000 487.650000 359.500000 488.350000 ;
      RECT 266.500000 487.650000 308.500000 488.350000 ;
      RECT 216.500000 487.650000 258.500000 488.350000 ;
      RECT 166.500000 487.650000 208.500000 488.350000 ;
      RECT 116.500000 487.650000 158.500000 488.350000 ;
      RECT 66.500000 487.650000 108.500000 488.350000 ;
      RECT 29.500000 487.650000 58.500000 488.350000 ;
      RECT 0.000000 487.650000 16.500000 488.350000 ;
      RECT 0.000000 487.170000 2.500000 487.650000 ;
      RECT 1166.500000 487.165000 1186.000000 489.650000 ;
      RECT 1166.500000 486.350000 1183.980000 487.165000 ;
      RECT 1157.500000 486.350000 1158.500000 487.650000 ;
      RECT 722.500000 486.350000 723.500000 487.650000 ;
      RECT 707.500000 486.350000 708.500000 487.650000 ;
      RECT 666.500000 486.350000 699.500000 487.650000 ;
      RECT 657.500000 486.350000 658.500000 487.650000 ;
      RECT 616.500000 486.350000 649.500000 487.650000 ;
      RECT 607.500000 486.350000 608.500000 487.650000 ;
      RECT 566.500000 486.350000 599.500000 487.650000 ;
      RECT 557.500000 486.350000 558.500000 487.650000 ;
      RECT 516.500000 486.350000 549.500000 487.650000 ;
      RECT 507.500000 486.350000 508.500000 487.650000 ;
      RECT 466.500000 486.350000 499.500000 487.650000 ;
      RECT 457.500000 486.350000 458.500000 487.650000 ;
      RECT 416.500000 486.350000 449.500000 487.650000 ;
      RECT 407.500000 486.350000 408.500000 487.650000 ;
      RECT 372.500000 486.350000 399.500000 487.650000 ;
      RECT 357.500000 486.350000 359.500000 487.650000 ;
      RECT 316.500000 486.350000 349.500000 487.650000 ;
      RECT 307.500000 486.350000 308.500000 487.650000 ;
      RECT 266.500000 486.350000 299.500000 487.650000 ;
      RECT 257.500000 486.350000 258.500000 487.650000 ;
      RECT 216.500000 486.350000 249.500000 487.650000 ;
      RECT 207.500000 486.350000 208.500000 487.650000 ;
      RECT 166.500000 486.350000 199.500000 487.650000 ;
      RECT 157.500000 486.350000 158.500000 487.650000 ;
      RECT 116.500000 486.350000 149.500000 487.650000 ;
      RECT 107.500000 486.350000 108.500000 487.650000 ;
      RECT 66.500000 486.350000 99.500000 487.650000 ;
      RECT 57.500000 486.350000 58.500000 487.650000 ;
      RECT 29.500000 486.350000 49.500000 487.650000 ;
      RECT 15.500000 486.350000 16.500000 487.650000 ;
      RECT 1157.500000 485.650000 1183.980000 486.350000 ;
      RECT 707.500000 485.650000 723.500000 486.350000 ;
      RECT 657.500000 485.650000 699.500000 486.350000 ;
      RECT 607.500000 485.650000 649.500000 486.350000 ;
      RECT 557.500000 485.650000 599.500000 486.350000 ;
      RECT 507.500000 485.650000 549.500000 486.350000 ;
      RECT 457.500000 485.650000 499.500000 486.350000 ;
      RECT 407.500000 485.650000 449.500000 486.350000 ;
      RECT 357.500000 485.650000 399.500000 486.350000 ;
      RECT 307.500000 485.650000 349.500000 486.350000 ;
      RECT 257.500000 485.650000 299.500000 486.350000 ;
      RECT 207.500000 485.650000 249.500000 486.350000 ;
      RECT 157.500000 485.650000 199.500000 486.350000 ;
      RECT 107.500000 485.650000 149.500000 486.350000 ;
      RECT 57.500000 485.650000 99.500000 486.350000 ;
      RECT 15.500000 485.650000 49.500000 486.350000 ;
      RECT 1157.500000 484.350000 1158.500000 485.650000 ;
      RECT 1139.000000 484.350000 1149.500000 487.650000 ;
      RECT 736.500000 484.350000 739.000000 487.650000 ;
      RECT 722.500000 484.350000 723.500000 485.650000 ;
      RECT 707.500000 484.350000 708.500000 485.650000 ;
      RECT 666.500000 484.350000 699.500000 485.650000 ;
      RECT 657.500000 484.350000 658.500000 485.650000 ;
      RECT 616.500000 484.350000 649.500000 485.650000 ;
      RECT 607.500000 484.350000 608.500000 485.650000 ;
      RECT 566.500000 484.350000 599.500000 485.650000 ;
      RECT 557.500000 484.350000 558.500000 485.650000 ;
      RECT 516.500000 484.350000 549.500000 485.650000 ;
      RECT 507.500000 484.350000 508.500000 485.650000 ;
      RECT 466.500000 484.350000 499.500000 485.650000 ;
      RECT 457.500000 484.350000 458.500000 485.650000 ;
      RECT 416.500000 484.350000 449.500000 485.650000 ;
      RECT 407.500000 484.350000 408.500000 485.650000 ;
      RECT 372.500000 484.350000 399.500000 485.650000 ;
      RECT 357.500000 484.350000 359.500000 485.650000 ;
      RECT 316.500000 484.350000 349.500000 485.650000 ;
      RECT 307.500000 484.350000 308.500000 485.650000 ;
      RECT 266.500000 484.350000 299.500000 485.650000 ;
      RECT 257.500000 484.350000 258.500000 485.650000 ;
      RECT 216.500000 484.350000 249.500000 485.650000 ;
      RECT 207.500000 484.350000 208.500000 485.650000 ;
      RECT 166.500000 484.350000 199.500000 485.650000 ;
      RECT 157.500000 484.350000 158.500000 485.650000 ;
      RECT 116.500000 484.350000 149.500000 485.650000 ;
      RECT 107.500000 484.350000 108.500000 485.650000 ;
      RECT 66.500000 484.350000 99.500000 485.650000 ;
      RECT 57.500000 484.350000 58.500000 485.650000 ;
      RECT 29.500000 484.350000 49.500000 485.650000 ;
      RECT 15.500000 484.350000 16.500000 485.650000 ;
      RECT 2.020000 484.350000 2.500000 487.170000 ;
      RECT 2.020000 484.070000 16.500000 484.350000 ;
      RECT 1166.500000 484.065000 1183.980000 485.650000 ;
      RECT 1139.000000 483.650000 1158.500000 484.350000 ;
      RECT 722.500000 483.650000 739.000000 484.350000 ;
      RECT 666.500000 483.650000 708.500000 484.350000 ;
      RECT 616.500000 483.650000 658.500000 484.350000 ;
      RECT 566.500000 483.650000 608.500000 484.350000 ;
      RECT 516.500000 483.650000 558.500000 484.350000 ;
      RECT 466.500000 483.650000 508.500000 484.350000 ;
      RECT 416.500000 483.650000 458.500000 484.350000 ;
      RECT 372.500000 483.650000 408.500000 484.350000 ;
      RECT 316.500000 483.650000 359.500000 484.350000 ;
      RECT 266.500000 483.650000 308.500000 484.350000 ;
      RECT 216.500000 483.650000 258.500000 484.350000 ;
      RECT 166.500000 483.650000 208.500000 484.350000 ;
      RECT 116.500000 483.650000 158.500000 484.350000 ;
      RECT 66.500000 483.650000 108.500000 484.350000 ;
      RECT 29.500000 483.650000 58.500000 484.350000 ;
      RECT 0.000000 483.650000 16.500000 484.070000 ;
      RECT 1166.500000 482.350000 1186.000000 484.065000 ;
      RECT 1157.500000 482.350000 1158.500000 483.650000 ;
      RECT 722.500000 482.350000 723.500000 483.650000 ;
      RECT 707.500000 482.350000 708.500000 483.650000 ;
      RECT 666.500000 482.350000 699.500000 483.650000 ;
      RECT 657.500000 482.350000 658.500000 483.650000 ;
      RECT 616.500000 482.350000 649.500000 483.650000 ;
      RECT 607.500000 482.350000 608.500000 483.650000 ;
      RECT 566.500000 482.350000 599.500000 483.650000 ;
      RECT 557.500000 482.350000 558.500000 483.650000 ;
      RECT 516.500000 482.350000 549.500000 483.650000 ;
      RECT 507.500000 482.350000 508.500000 483.650000 ;
      RECT 466.500000 482.350000 499.500000 483.650000 ;
      RECT 457.500000 482.350000 458.500000 483.650000 ;
      RECT 416.500000 482.350000 449.500000 483.650000 ;
      RECT 407.500000 482.350000 408.500000 483.650000 ;
      RECT 372.500000 482.350000 399.500000 483.650000 ;
      RECT 357.500000 482.350000 359.500000 483.650000 ;
      RECT 316.500000 482.350000 349.500000 483.650000 ;
      RECT 307.500000 482.350000 308.500000 483.650000 ;
      RECT 266.500000 482.350000 299.500000 483.650000 ;
      RECT 257.500000 482.350000 258.500000 483.650000 ;
      RECT 216.500000 482.350000 249.500000 483.650000 ;
      RECT 207.500000 482.350000 208.500000 483.650000 ;
      RECT 166.500000 482.350000 199.500000 483.650000 ;
      RECT 157.500000 482.350000 158.500000 483.650000 ;
      RECT 116.500000 482.350000 149.500000 483.650000 ;
      RECT 107.500000 482.350000 108.500000 483.650000 ;
      RECT 66.500000 482.350000 99.500000 483.650000 ;
      RECT 57.500000 482.350000 58.500000 483.650000 ;
      RECT 29.500000 482.350000 49.500000 483.650000 ;
      RECT 15.500000 482.350000 16.500000 483.650000 ;
      RECT 1157.500000 481.650000 1186.000000 482.350000 ;
      RECT 707.500000 481.650000 723.500000 482.350000 ;
      RECT 657.500000 481.650000 699.500000 482.350000 ;
      RECT 607.500000 481.650000 649.500000 482.350000 ;
      RECT 557.500000 481.650000 599.500000 482.350000 ;
      RECT 507.500000 481.650000 549.500000 482.350000 ;
      RECT 457.500000 481.650000 499.500000 482.350000 ;
      RECT 407.500000 481.650000 449.500000 482.350000 ;
      RECT 357.500000 481.650000 399.500000 482.350000 ;
      RECT 307.500000 481.650000 349.500000 482.350000 ;
      RECT 257.500000 481.650000 299.500000 482.350000 ;
      RECT 207.500000 481.650000 249.500000 482.350000 ;
      RECT 157.500000 481.650000 199.500000 482.350000 ;
      RECT 107.500000 481.650000 149.500000 482.350000 ;
      RECT 57.500000 481.650000 99.500000 482.350000 ;
      RECT 15.500000 481.650000 49.500000 482.350000 ;
      RECT 1166.500000 481.485000 1186.000000 481.650000 ;
      RECT 1157.500000 480.350000 1158.500000 481.650000 ;
      RECT 1139.000000 480.350000 1149.500000 483.650000 ;
      RECT 736.500000 480.350000 739.000000 483.650000 ;
      RECT 722.500000 480.350000 723.500000 481.650000 ;
      RECT 707.500000 480.350000 708.500000 481.650000 ;
      RECT 666.500000 480.350000 699.500000 481.650000 ;
      RECT 657.500000 480.350000 658.500000 481.650000 ;
      RECT 616.500000 480.350000 649.500000 481.650000 ;
      RECT 607.500000 480.350000 608.500000 481.650000 ;
      RECT 566.500000 480.350000 599.500000 481.650000 ;
      RECT 557.500000 480.350000 558.500000 481.650000 ;
      RECT 516.500000 480.350000 549.500000 481.650000 ;
      RECT 507.500000 480.350000 508.500000 481.650000 ;
      RECT 466.500000 480.350000 499.500000 481.650000 ;
      RECT 457.500000 480.350000 458.500000 481.650000 ;
      RECT 416.500000 480.350000 449.500000 481.650000 ;
      RECT 407.500000 480.350000 408.500000 481.650000 ;
      RECT 372.500000 480.350000 399.500000 481.650000 ;
      RECT 357.500000 480.350000 359.500000 481.650000 ;
      RECT 316.500000 480.350000 349.500000 481.650000 ;
      RECT 307.500000 480.350000 308.500000 481.650000 ;
      RECT 266.500000 480.350000 299.500000 481.650000 ;
      RECT 257.500000 480.350000 258.500000 481.650000 ;
      RECT 216.500000 480.350000 249.500000 481.650000 ;
      RECT 207.500000 480.350000 208.500000 481.650000 ;
      RECT 166.500000 480.350000 199.500000 481.650000 ;
      RECT 157.500000 480.350000 158.500000 481.650000 ;
      RECT 116.500000 480.350000 149.500000 481.650000 ;
      RECT 107.500000 480.350000 108.500000 481.650000 ;
      RECT 66.500000 480.350000 99.500000 481.650000 ;
      RECT 57.500000 480.350000 58.500000 481.650000 ;
      RECT 29.500000 480.350000 49.500000 481.650000 ;
      RECT 15.500000 480.350000 16.500000 481.650000 ;
      RECT 0.000000 480.350000 2.500000 483.650000 ;
      RECT 1139.000000 479.650000 1158.500000 480.350000 ;
      RECT 722.500000 479.650000 739.000000 480.350000 ;
      RECT 666.500000 479.650000 708.500000 480.350000 ;
      RECT 616.500000 479.650000 658.500000 480.350000 ;
      RECT 566.500000 479.650000 608.500000 480.350000 ;
      RECT 516.500000 479.650000 558.500000 480.350000 ;
      RECT 466.500000 479.650000 508.500000 480.350000 ;
      RECT 416.500000 479.650000 458.500000 480.350000 ;
      RECT 372.500000 479.650000 408.500000 480.350000 ;
      RECT 316.500000 479.650000 359.500000 480.350000 ;
      RECT 266.500000 479.650000 308.500000 480.350000 ;
      RECT 216.500000 479.650000 258.500000 480.350000 ;
      RECT 166.500000 479.650000 208.500000 480.350000 ;
      RECT 116.500000 479.650000 158.500000 480.350000 ;
      RECT 66.500000 479.650000 108.500000 480.350000 ;
      RECT 29.500000 479.650000 58.500000 480.350000 ;
      RECT 0.000000 479.650000 16.500000 480.350000 ;
      RECT 1166.500000 478.385000 1183.980000 481.485000 ;
      RECT 1166.500000 478.350000 1186.000000 478.385000 ;
      RECT 1157.500000 478.350000 1158.500000 479.650000 ;
      RECT 722.500000 478.350000 723.500000 479.650000 ;
      RECT 707.500000 478.350000 708.500000 479.650000 ;
      RECT 666.500000 478.350000 699.500000 479.650000 ;
      RECT 657.500000 478.350000 658.500000 479.650000 ;
      RECT 616.500000 478.350000 649.500000 479.650000 ;
      RECT 607.500000 478.350000 608.500000 479.650000 ;
      RECT 566.500000 478.350000 599.500000 479.650000 ;
      RECT 557.500000 478.350000 558.500000 479.650000 ;
      RECT 516.500000 478.350000 549.500000 479.650000 ;
      RECT 507.500000 478.350000 508.500000 479.650000 ;
      RECT 466.500000 478.350000 499.500000 479.650000 ;
      RECT 457.500000 478.350000 458.500000 479.650000 ;
      RECT 416.500000 478.350000 449.500000 479.650000 ;
      RECT 407.500000 478.350000 408.500000 479.650000 ;
      RECT 372.500000 478.350000 399.500000 479.650000 ;
      RECT 357.500000 478.350000 359.500000 479.650000 ;
      RECT 316.500000 478.350000 349.500000 479.650000 ;
      RECT 307.500000 478.350000 308.500000 479.650000 ;
      RECT 266.500000 478.350000 299.500000 479.650000 ;
      RECT 257.500000 478.350000 258.500000 479.650000 ;
      RECT 216.500000 478.350000 249.500000 479.650000 ;
      RECT 207.500000 478.350000 208.500000 479.650000 ;
      RECT 166.500000 478.350000 199.500000 479.650000 ;
      RECT 157.500000 478.350000 158.500000 479.650000 ;
      RECT 116.500000 478.350000 149.500000 479.650000 ;
      RECT 107.500000 478.350000 108.500000 479.650000 ;
      RECT 66.500000 478.350000 99.500000 479.650000 ;
      RECT 57.500000 478.350000 58.500000 479.650000 ;
      RECT 29.500000 478.350000 49.500000 479.650000 ;
      RECT 15.500000 478.350000 16.500000 479.650000 ;
      RECT 1157.500000 477.650000 1186.000000 478.350000 ;
      RECT 707.500000 477.650000 723.500000 478.350000 ;
      RECT 657.500000 477.650000 699.500000 478.350000 ;
      RECT 607.500000 477.650000 649.500000 478.350000 ;
      RECT 557.500000 477.650000 599.500000 478.350000 ;
      RECT 507.500000 477.650000 549.500000 478.350000 ;
      RECT 457.500000 477.650000 499.500000 478.350000 ;
      RECT 407.500000 477.650000 449.500000 478.350000 ;
      RECT 357.500000 477.650000 399.500000 478.350000 ;
      RECT 307.500000 477.650000 349.500000 478.350000 ;
      RECT 257.500000 477.650000 299.500000 478.350000 ;
      RECT 207.500000 477.650000 249.500000 478.350000 ;
      RECT 157.500000 477.650000 199.500000 478.350000 ;
      RECT 107.500000 477.650000 149.500000 478.350000 ;
      RECT 57.500000 477.650000 99.500000 478.350000 ;
      RECT 15.500000 477.650000 49.500000 478.350000 ;
      RECT 1166.500000 477.525000 1186.000000 477.650000 ;
      RECT 0.000000 476.575000 2.500000 479.650000 ;
      RECT 1157.500000 476.350000 1158.500000 477.650000 ;
      RECT 1139.000000 476.350000 1149.500000 479.650000 ;
      RECT 736.500000 476.350000 739.000000 479.650000 ;
      RECT 722.500000 476.350000 723.500000 477.650000 ;
      RECT 707.500000 476.350000 708.500000 477.650000 ;
      RECT 666.500000 476.350000 699.500000 477.650000 ;
      RECT 657.500000 476.350000 658.500000 477.650000 ;
      RECT 616.500000 476.350000 649.500000 477.650000 ;
      RECT 607.500000 476.350000 608.500000 477.650000 ;
      RECT 566.500000 476.350000 599.500000 477.650000 ;
      RECT 557.500000 476.350000 558.500000 477.650000 ;
      RECT 516.500000 476.350000 549.500000 477.650000 ;
      RECT 507.500000 476.350000 508.500000 477.650000 ;
      RECT 466.500000 476.350000 499.500000 477.650000 ;
      RECT 457.500000 476.350000 458.500000 477.650000 ;
      RECT 416.500000 476.350000 449.500000 477.650000 ;
      RECT 407.500000 476.350000 408.500000 477.650000 ;
      RECT 370.000000 476.350000 399.500000 477.650000 ;
      RECT 357.500000 476.350000 362.000000 477.650000 ;
      RECT 316.500000 476.350000 349.500000 477.650000 ;
      RECT 307.500000 476.350000 308.500000 477.650000 ;
      RECT 266.500000 476.350000 299.500000 477.650000 ;
      RECT 257.500000 476.350000 258.500000 477.650000 ;
      RECT 216.500000 476.350000 249.500000 477.650000 ;
      RECT 207.500000 476.350000 208.500000 477.650000 ;
      RECT 166.500000 476.350000 199.500000 477.650000 ;
      RECT 157.500000 476.350000 158.500000 477.650000 ;
      RECT 116.500000 476.350000 149.500000 477.650000 ;
      RECT 107.500000 476.350000 108.500000 477.650000 ;
      RECT 66.500000 476.350000 99.500000 477.650000 ;
      RECT 57.500000 476.350000 58.500000 477.650000 ;
      RECT 29.500000 476.350000 49.500000 477.650000 ;
      RECT 15.500000 476.350000 16.500000 477.650000 ;
      RECT 2.020000 476.350000 2.500000 476.575000 ;
      RECT 1139.000000 475.650000 1158.500000 476.350000 ;
      RECT 722.500000 475.650000 739.000000 476.350000 ;
      RECT 666.500000 475.650000 708.500000 476.350000 ;
      RECT 616.500000 475.650000 658.500000 476.350000 ;
      RECT 566.500000 475.650000 608.500000 476.350000 ;
      RECT 516.500000 475.650000 558.500000 476.350000 ;
      RECT 466.500000 475.650000 508.500000 476.350000 ;
      RECT 416.500000 475.650000 458.500000 476.350000 ;
      RECT 370.000000 475.650000 408.500000 476.350000 ;
      RECT 316.500000 475.650000 362.000000 476.350000 ;
      RECT 266.500000 475.650000 308.500000 476.350000 ;
      RECT 216.500000 475.650000 258.500000 476.350000 ;
      RECT 166.500000 475.650000 208.500000 476.350000 ;
      RECT 116.500000 475.650000 158.500000 476.350000 ;
      RECT 66.500000 475.650000 108.500000 476.350000 ;
      RECT 29.500000 475.650000 58.500000 476.350000 ;
      RECT 2.020000 475.650000 16.500000 476.350000 ;
      RECT 1166.500000 474.425000 1183.980000 477.525000 ;
      RECT 1166.500000 474.350000 1186.000000 474.425000 ;
      RECT 1157.500000 474.350000 1158.500000 475.650000 ;
      RECT 722.500000 474.350000 723.500000 475.650000 ;
      RECT 707.500000 474.350000 708.500000 475.650000 ;
      RECT 666.500000 474.350000 699.500000 475.650000 ;
      RECT 657.500000 474.350000 658.500000 475.650000 ;
      RECT 616.500000 474.350000 649.500000 475.650000 ;
      RECT 607.500000 474.350000 608.500000 475.650000 ;
      RECT 566.500000 474.350000 599.500000 475.650000 ;
      RECT 557.500000 474.350000 558.500000 475.650000 ;
      RECT 516.500000 474.350000 549.500000 475.650000 ;
      RECT 507.500000 474.350000 508.500000 475.650000 ;
      RECT 466.500000 474.350000 499.500000 475.650000 ;
      RECT 457.500000 474.350000 458.500000 475.650000 ;
      RECT 416.500000 474.350000 449.500000 475.650000 ;
      RECT 407.500000 474.350000 408.500000 475.650000 ;
      RECT 370.000000 474.350000 399.500000 475.650000 ;
      RECT 357.500000 474.350000 362.000000 475.650000 ;
      RECT 316.500000 474.350000 349.500000 475.650000 ;
      RECT 307.500000 474.350000 308.500000 475.650000 ;
      RECT 266.500000 474.350000 299.500000 475.650000 ;
      RECT 257.500000 474.350000 258.500000 475.650000 ;
      RECT 216.500000 474.350000 249.500000 475.650000 ;
      RECT 207.500000 474.350000 208.500000 475.650000 ;
      RECT 166.500000 474.350000 199.500000 475.650000 ;
      RECT 157.500000 474.350000 158.500000 475.650000 ;
      RECT 116.500000 474.350000 149.500000 475.650000 ;
      RECT 107.500000 474.350000 108.500000 475.650000 ;
      RECT 66.500000 474.350000 99.500000 475.650000 ;
      RECT 57.500000 474.350000 58.500000 475.650000 ;
      RECT 29.500000 474.350000 49.500000 475.650000 ;
      RECT 15.500000 474.350000 16.500000 475.650000 ;
      RECT 1157.500000 473.650000 1186.000000 474.350000 ;
      RECT 707.500000 473.650000 723.500000 474.350000 ;
      RECT 657.500000 473.650000 699.500000 474.350000 ;
      RECT 607.500000 473.650000 649.500000 474.350000 ;
      RECT 557.500000 473.650000 599.500000 474.350000 ;
      RECT 507.500000 473.650000 549.500000 474.350000 ;
      RECT 457.500000 473.650000 499.500000 474.350000 ;
      RECT 407.500000 473.650000 449.500000 474.350000 ;
      RECT 357.500000 473.650000 399.500000 474.350000 ;
      RECT 307.500000 473.650000 349.500000 474.350000 ;
      RECT 257.500000 473.650000 299.500000 474.350000 ;
      RECT 207.500000 473.650000 249.500000 474.350000 ;
      RECT 157.500000 473.650000 199.500000 474.350000 ;
      RECT 107.500000 473.650000 149.500000 474.350000 ;
      RECT 57.500000 473.650000 99.500000 474.350000 ;
      RECT 15.500000 473.650000 49.500000 474.350000 ;
      RECT 2.020000 473.475000 2.500000 475.650000 ;
      RECT 0.000000 472.615000 2.500000 473.475000 ;
      RECT 1157.500000 472.350000 1158.500000 473.650000 ;
      RECT 1139.000000 472.350000 1149.500000 475.650000 ;
      RECT 736.500000 472.350000 739.000000 475.650000 ;
      RECT 722.500000 472.350000 723.500000 473.650000 ;
      RECT 707.500000 472.350000 708.500000 473.650000 ;
      RECT 666.500000 472.350000 699.500000 473.650000 ;
      RECT 657.500000 472.350000 658.500000 473.650000 ;
      RECT 616.500000 472.350000 649.500000 473.650000 ;
      RECT 607.500000 472.350000 608.500000 473.650000 ;
      RECT 566.500000 472.350000 599.500000 473.650000 ;
      RECT 557.500000 472.350000 558.500000 473.650000 ;
      RECT 516.500000 472.350000 549.500000 473.650000 ;
      RECT 507.500000 472.350000 508.500000 473.650000 ;
      RECT 466.500000 472.350000 499.500000 473.650000 ;
      RECT 457.500000 472.350000 458.500000 473.650000 ;
      RECT 416.500000 472.350000 449.500000 473.650000 ;
      RECT 407.500000 472.350000 408.500000 473.650000 ;
      RECT 370.000000 472.350000 399.500000 473.650000 ;
      RECT 357.500000 472.350000 358.500000 473.650000 ;
      RECT 316.500000 472.350000 349.500000 473.650000 ;
      RECT 307.500000 472.350000 308.500000 473.650000 ;
      RECT 266.500000 472.350000 299.500000 473.650000 ;
      RECT 257.500000 472.350000 258.500000 473.650000 ;
      RECT 216.500000 472.350000 249.500000 473.650000 ;
      RECT 207.500000 472.350000 208.500000 473.650000 ;
      RECT 166.500000 472.350000 199.500000 473.650000 ;
      RECT 157.500000 472.350000 158.500000 473.650000 ;
      RECT 116.500000 472.350000 149.500000 473.650000 ;
      RECT 107.500000 472.350000 108.500000 473.650000 ;
      RECT 66.500000 472.350000 99.500000 473.650000 ;
      RECT 57.500000 472.350000 58.500000 473.650000 ;
      RECT 29.500000 472.350000 49.500000 473.650000 ;
      RECT 15.500000 472.350000 16.500000 473.650000 ;
      RECT 2.020000 472.350000 2.500000 472.615000 ;
      RECT 1139.000000 471.650000 1158.500000 472.350000 ;
      RECT 722.500000 471.650000 739.000000 472.350000 ;
      RECT 666.500000 471.650000 708.500000 472.350000 ;
      RECT 616.500000 471.650000 658.500000 472.350000 ;
      RECT 566.500000 471.650000 608.500000 472.350000 ;
      RECT 516.500000 471.650000 558.500000 472.350000 ;
      RECT 466.500000 471.650000 508.500000 472.350000 ;
      RECT 416.500000 471.650000 458.500000 472.350000 ;
      RECT 370.000000 471.650000 408.500000 472.350000 ;
      RECT 316.500000 471.650000 358.500000 472.350000 ;
      RECT 266.500000 471.650000 308.500000 472.350000 ;
      RECT 216.500000 471.650000 258.500000 472.350000 ;
      RECT 166.500000 471.650000 208.500000 472.350000 ;
      RECT 116.500000 471.650000 158.500000 472.350000 ;
      RECT 66.500000 471.650000 108.500000 472.350000 ;
      RECT 29.500000 471.650000 58.500000 472.350000 ;
      RECT 2.020000 471.650000 16.500000 472.350000 ;
      RECT 1166.500000 470.350000 1186.000000 473.650000 ;
      RECT 1157.500000 470.350000 1158.500000 471.650000 ;
      RECT 722.500000 470.350000 723.500000 471.650000 ;
      RECT 707.500000 470.350000 708.500000 471.650000 ;
      RECT 666.500000 470.350000 699.500000 471.650000 ;
      RECT 657.500000 470.350000 658.500000 471.650000 ;
      RECT 616.500000 470.350000 649.500000 471.650000 ;
      RECT 607.500000 470.350000 608.500000 471.650000 ;
      RECT 566.500000 470.350000 599.500000 471.650000 ;
      RECT 557.500000 470.350000 558.500000 471.650000 ;
      RECT 516.500000 470.350000 549.500000 471.650000 ;
      RECT 507.500000 470.350000 508.500000 471.650000 ;
      RECT 466.500000 470.350000 499.500000 471.650000 ;
      RECT 457.500000 470.350000 458.500000 471.650000 ;
      RECT 416.500000 470.350000 449.500000 471.650000 ;
      RECT 407.500000 470.350000 408.500000 471.650000 ;
      RECT 370.000000 470.350000 399.500000 471.650000 ;
      RECT 357.500000 470.350000 358.500000 471.650000 ;
      RECT 316.500000 470.350000 349.500000 471.650000 ;
      RECT 307.500000 470.350000 308.500000 471.650000 ;
      RECT 266.500000 470.350000 299.500000 471.650000 ;
      RECT 257.500000 470.350000 258.500000 471.650000 ;
      RECT 216.500000 470.350000 249.500000 471.650000 ;
      RECT 207.500000 470.350000 208.500000 471.650000 ;
      RECT 166.500000 470.350000 199.500000 471.650000 ;
      RECT 157.500000 470.350000 158.500000 471.650000 ;
      RECT 116.500000 470.350000 149.500000 471.650000 ;
      RECT 107.500000 470.350000 108.500000 471.650000 ;
      RECT 66.500000 470.350000 99.500000 471.650000 ;
      RECT 57.500000 470.350000 58.500000 471.650000 ;
      RECT 29.500000 470.350000 49.500000 471.650000 ;
      RECT 15.500000 470.350000 16.500000 471.650000 ;
      RECT 1157.500000 469.650000 1186.000000 470.350000 ;
      RECT 707.500000 469.650000 723.500000 470.350000 ;
      RECT 657.500000 469.650000 699.500000 470.350000 ;
      RECT 607.500000 469.650000 649.500000 470.350000 ;
      RECT 557.500000 469.650000 599.500000 470.350000 ;
      RECT 507.500000 469.650000 549.500000 470.350000 ;
      RECT 457.500000 469.650000 499.500000 470.350000 ;
      RECT 407.500000 469.650000 449.500000 470.350000 ;
      RECT 357.500000 469.650000 399.500000 470.350000 ;
      RECT 307.500000 469.650000 349.500000 470.350000 ;
      RECT 257.500000 469.650000 299.500000 470.350000 ;
      RECT 207.500000 469.650000 249.500000 470.350000 ;
      RECT 157.500000 469.650000 199.500000 470.350000 ;
      RECT 107.500000 469.650000 149.500000 470.350000 ;
      RECT 57.500000 469.650000 99.500000 470.350000 ;
      RECT 15.500000 469.650000 49.500000 470.350000 ;
      RECT 2.020000 469.515000 2.500000 471.650000 ;
      RECT 1157.500000 468.350000 1158.500000 469.650000 ;
      RECT 1139.000000 468.350000 1149.500000 471.650000 ;
      RECT 736.500000 468.350000 739.000000 471.650000 ;
      RECT 722.500000 468.350000 723.500000 469.650000 ;
      RECT 707.500000 468.350000 708.500000 469.650000 ;
      RECT 666.500000 468.350000 699.500000 469.650000 ;
      RECT 657.500000 468.350000 658.500000 469.650000 ;
      RECT 616.500000 468.350000 649.500000 469.650000 ;
      RECT 607.500000 468.350000 608.500000 469.650000 ;
      RECT 566.500000 468.350000 599.500000 469.650000 ;
      RECT 557.500000 468.350000 558.500000 469.650000 ;
      RECT 516.500000 468.350000 549.500000 469.650000 ;
      RECT 507.500000 468.350000 508.500000 469.650000 ;
      RECT 466.500000 468.350000 499.500000 469.650000 ;
      RECT 457.500000 468.350000 458.500000 469.650000 ;
      RECT 416.500000 468.350000 449.500000 469.650000 ;
      RECT 407.500000 468.350000 408.500000 469.650000 ;
      RECT 366.500000 468.350000 399.500000 469.650000 ;
      RECT 357.500000 468.350000 358.500000 469.650000 ;
      RECT 316.500000 468.350000 349.500000 469.650000 ;
      RECT 307.500000 468.350000 308.500000 469.650000 ;
      RECT 266.500000 468.350000 299.500000 469.650000 ;
      RECT 257.500000 468.350000 258.500000 469.650000 ;
      RECT 216.500000 468.350000 249.500000 469.650000 ;
      RECT 207.500000 468.350000 208.500000 469.650000 ;
      RECT 166.500000 468.350000 199.500000 469.650000 ;
      RECT 157.500000 468.350000 158.500000 469.650000 ;
      RECT 116.500000 468.350000 149.500000 469.650000 ;
      RECT 107.500000 468.350000 108.500000 469.650000 ;
      RECT 66.500000 468.350000 99.500000 469.650000 ;
      RECT 57.500000 468.350000 58.500000 469.650000 ;
      RECT 29.500000 468.350000 49.500000 469.650000 ;
      RECT 15.500000 468.350000 16.500000 469.650000 ;
      RECT 0.000000 468.350000 2.500000 469.515000 ;
      RECT 1139.000000 467.650000 1158.500000 468.350000 ;
      RECT 722.500000 467.650000 739.000000 468.350000 ;
      RECT 666.500000 467.650000 708.500000 468.350000 ;
      RECT 616.500000 467.650000 658.500000 468.350000 ;
      RECT 566.500000 467.650000 608.500000 468.350000 ;
      RECT 516.500000 467.650000 558.500000 468.350000 ;
      RECT 466.500000 467.650000 508.500000 468.350000 ;
      RECT 416.500000 467.650000 458.500000 468.350000 ;
      RECT 366.500000 467.650000 408.500000 468.350000 ;
      RECT 316.500000 467.650000 358.500000 468.350000 ;
      RECT 266.500000 467.650000 308.500000 468.350000 ;
      RECT 216.500000 467.650000 258.500000 468.350000 ;
      RECT 166.500000 467.650000 208.500000 468.350000 ;
      RECT 116.500000 467.650000 158.500000 468.350000 ;
      RECT 66.500000 467.650000 108.500000 468.350000 ;
      RECT 29.500000 467.650000 58.500000 468.350000 ;
      RECT 0.000000 467.650000 16.500000 468.350000 ;
      RECT 0.000000 466.935000 2.500000 467.650000 ;
      RECT 1166.500000 466.930000 1186.000000 469.650000 ;
      RECT 1166.500000 466.350000 1183.980000 466.930000 ;
      RECT 1157.500000 466.350000 1158.500000 467.650000 ;
      RECT 722.500000 466.350000 723.500000 467.650000 ;
      RECT 707.500000 466.350000 708.500000 467.650000 ;
      RECT 666.500000 466.350000 699.500000 467.650000 ;
      RECT 657.500000 466.350000 658.500000 467.650000 ;
      RECT 616.500000 466.350000 649.500000 467.650000 ;
      RECT 607.500000 466.350000 608.500000 467.650000 ;
      RECT 566.500000 466.350000 599.500000 467.650000 ;
      RECT 557.500000 466.350000 558.500000 467.650000 ;
      RECT 516.500000 466.350000 549.500000 467.650000 ;
      RECT 507.500000 466.350000 508.500000 467.650000 ;
      RECT 466.500000 466.350000 499.500000 467.650000 ;
      RECT 457.500000 466.350000 458.500000 467.650000 ;
      RECT 416.500000 466.350000 449.500000 467.650000 ;
      RECT 407.500000 466.350000 408.500000 467.650000 ;
      RECT 366.500000 466.350000 399.500000 467.650000 ;
      RECT 357.500000 466.350000 358.500000 467.650000 ;
      RECT 316.500000 466.350000 349.500000 467.650000 ;
      RECT 307.500000 466.350000 308.500000 467.650000 ;
      RECT 266.500000 466.350000 299.500000 467.650000 ;
      RECT 257.500000 466.350000 258.500000 467.650000 ;
      RECT 216.500000 466.350000 249.500000 467.650000 ;
      RECT 207.500000 466.350000 208.500000 467.650000 ;
      RECT 166.500000 466.350000 199.500000 467.650000 ;
      RECT 157.500000 466.350000 158.500000 467.650000 ;
      RECT 116.500000 466.350000 149.500000 467.650000 ;
      RECT 107.500000 466.350000 108.500000 467.650000 ;
      RECT 66.500000 466.350000 99.500000 467.650000 ;
      RECT 57.500000 466.350000 58.500000 467.650000 ;
      RECT 29.500000 466.350000 49.500000 467.650000 ;
      RECT 15.500000 466.350000 16.500000 467.650000 ;
      RECT 1157.500000 465.650000 1183.980000 466.350000 ;
      RECT 707.500000 465.650000 723.500000 466.350000 ;
      RECT 657.500000 465.650000 699.500000 466.350000 ;
      RECT 607.500000 465.650000 649.500000 466.350000 ;
      RECT 557.500000 465.650000 599.500000 466.350000 ;
      RECT 507.500000 465.650000 549.500000 466.350000 ;
      RECT 457.500000 465.650000 499.500000 466.350000 ;
      RECT 407.500000 465.650000 449.500000 466.350000 ;
      RECT 357.500000 465.650000 399.500000 466.350000 ;
      RECT 307.500000 465.650000 349.500000 466.350000 ;
      RECT 257.500000 465.650000 299.500000 466.350000 ;
      RECT 207.500000 465.650000 249.500000 466.350000 ;
      RECT 157.500000 465.650000 199.500000 466.350000 ;
      RECT 107.500000 465.650000 149.500000 466.350000 ;
      RECT 57.500000 465.650000 99.500000 466.350000 ;
      RECT 15.500000 465.650000 49.500000 466.350000 ;
      RECT 1157.500000 464.350000 1158.500000 465.650000 ;
      RECT 1139.000000 464.350000 1149.500000 467.650000 ;
      RECT 736.500000 464.350000 739.000000 467.650000 ;
      RECT 722.500000 464.350000 723.500000 465.650000 ;
      RECT 707.500000 464.350000 708.500000 465.650000 ;
      RECT 666.500000 464.350000 699.500000 465.650000 ;
      RECT 657.500000 464.350000 658.500000 465.650000 ;
      RECT 616.500000 464.350000 649.500000 465.650000 ;
      RECT 607.500000 464.350000 608.500000 465.650000 ;
      RECT 566.500000 464.350000 599.500000 465.650000 ;
      RECT 557.500000 464.350000 558.500000 465.650000 ;
      RECT 516.500000 464.350000 549.500000 465.650000 ;
      RECT 507.500000 464.350000 508.500000 465.650000 ;
      RECT 466.500000 464.350000 499.500000 465.650000 ;
      RECT 457.500000 464.350000 458.500000 465.650000 ;
      RECT 416.500000 464.350000 449.500000 465.650000 ;
      RECT 407.500000 464.350000 408.500000 465.650000 ;
      RECT 366.500000 464.350000 399.500000 465.650000 ;
      RECT 357.500000 464.350000 358.500000 465.650000 ;
      RECT 316.500000 464.350000 349.500000 465.650000 ;
      RECT 307.500000 464.350000 308.500000 465.650000 ;
      RECT 266.500000 464.350000 299.500000 465.650000 ;
      RECT 257.500000 464.350000 258.500000 465.650000 ;
      RECT 216.500000 464.350000 249.500000 465.650000 ;
      RECT 207.500000 464.350000 208.500000 465.650000 ;
      RECT 166.500000 464.350000 199.500000 465.650000 ;
      RECT 157.500000 464.350000 158.500000 465.650000 ;
      RECT 116.500000 464.350000 149.500000 465.650000 ;
      RECT 107.500000 464.350000 108.500000 465.650000 ;
      RECT 66.500000 464.350000 99.500000 465.650000 ;
      RECT 57.500000 464.350000 58.500000 465.650000 ;
      RECT 29.500000 464.350000 49.500000 465.650000 ;
      RECT 15.500000 464.350000 16.500000 465.650000 ;
      RECT 2.020000 464.350000 2.500000 466.935000 ;
      RECT 2.020000 463.835000 16.500000 464.350000 ;
      RECT 1166.500000 463.830000 1183.980000 465.650000 ;
      RECT 1139.000000 463.650000 1158.500000 464.350000 ;
      RECT 722.500000 463.650000 739.000000 464.350000 ;
      RECT 666.500000 463.650000 708.500000 464.350000 ;
      RECT 616.500000 463.650000 658.500000 464.350000 ;
      RECT 566.500000 463.650000 608.500000 464.350000 ;
      RECT 516.500000 463.650000 558.500000 464.350000 ;
      RECT 466.500000 463.650000 508.500000 464.350000 ;
      RECT 416.500000 463.650000 458.500000 464.350000 ;
      RECT 366.500000 463.650000 408.500000 464.350000 ;
      RECT 316.500000 463.650000 358.500000 464.350000 ;
      RECT 266.500000 463.650000 308.500000 464.350000 ;
      RECT 216.500000 463.650000 258.500000 464.350000 ;
      RECT 166.500000 463.650000 208.500000 464.350000 ;
      RECT 116.500000 463.650000 158.500000 464.350000 ;
      RECT 66.500000 463.650000 108.500000 464.350000 ;
      RECT 29.500000 463.650000 58.500000 464.350000 ;
      RECT 0.000000 463.650000 16.500000 463.835000 ;
      RECT 1166.500000 462.350000 1186.000000 463.830000 ;
      RECT 1157.500000 462.350000 1158.500000 463.650000 ;
      RECT 722.500000 462.350000 723.500000 463.650000 ;
      RECT 707.500000 462.350000 708.500000 463.650000 ;
      RECT 666.500000 462.350000 699.500000 463.650000 ;
      RECT 657.500000 462.350000 658.500000 463.650000 ;
      RECT 616.500000 462.350000 649.500000 463.650000 ;
      RECT 607.500000 462.350000 608.500000 463.650000 ;
      RECT 566.500000 462.350000 599.500000 463.650000 ;
      RECT 557.500000 462.350000 558.500000 463.650000 ;
      RECT 516.500000 462.350000 549.500000 463.650000 ;
      RECT 507.500000 462.350000 508.500000 463.650000 ;
      RECT 466.500000 462.350000 499.500000 463.650000 ;
      RECT 457.500000 462.350000 458.500000 463.650000 ;
      RECT 416.500000 462.350000 449.500000 463.650000 ;
      RECT 407.500000 462.350000 408.500000 463.650000 ;
      RECT 366.500000 462.350000 399.500000 463.650000 ;
      RECT 357.500000 462.350000 358.500000 463.650000 ;
      RECT 316.500000 462.350000 349.500000 463.650000 ;
      RECT 307.500000 462.350000 308.500000 463.650000 ;
      RECT 266.500000 462.350000 299.500000 463.650000 ;
      RECT 257.500000 462.350000 258.500000 463.650000 ;
      RECT 216.500000 462.350000 249.500000 463.650000 ;
      RECT 207.500000 462.350000 208.500000 463.650000 ;
      RECT 166.500000 462.350000 199.500000 463.650000 ;
      RECT 157.500000 462.350000 158.500000 463.650000 ;
      RECT 116.500000 462.350000 149.500000 463.650000 ;
      RECT 107.500000 462.350000 108.500000 463.650000 ;
      RECT 66.500000 462.350000 99.500000 463.650000 ;
      RECT 57.500000 462.350000 58.500000 463.650000 ;
      RECT 29.500000 462.350000 49.500000 463.650000 ;
      RECT 15.500000 462.350000 16.500000 463.650000 ;
      RECT 1157.500000 461.650000 1186.000000 462.350000 ;
      RECT 707.500000 461.650000 723.500000 462.350000 ;
      RECT 657.500000 461.650000 699.500000 462.350000 ;
      RECT 607.500000 461.650000 649.500000 462.350000 ;
      RECT 557.500000 461.650000 599.500000 462.350000 ;
      RECT 507.500000 461.650000 549.500000 462.350000 ;
      RECT 457.500000 461.650000 499.500000 462.350000 ;
      RECT 407.500000 461.650000 449.500000 462.350000 ;
      RECT 357.500000 461.650000 399.500000 462.350000 ;
      RECT 307.500000 461.650000 349.500000 462.350000 ;
      RECT 207.500000 461.650000 249.500000 462.350000 ;
      RECT 107.500000 461.650000 149.500000 462.350000 ;
      RECT 57.500000 461.650000 99.500000 462.350000 ;
      RECT 15.500000 461.650000 49.500000 462.350000 ;
      RECT 1157.500000 460.350000 1158.500000 461.650000 ;
      RECT 1139.000000 460.350000 1149.500000 463.650000 ;
      RECT 736.500000 460.350000 739.000000 463.650000 ;
      RECT 722.500000 460.350000 723.500000 461.650000 ;
      RECT 707.500000 460.350000 708.500000 461.650000 ;
      RECT 666.500000 460.350000 699.500000 461.650000 ;
      RECT 657.500000 460.350000 658.500000 461.650000 ;
      RECT 616.500000 460.350000 649.500000 461.650000 ;
      RECT 607.500000 460.350000 608.500000 461.650000 ;
      RECT 566.500000 460.350000 599.500000 461.650000 ;
      RECT 557.500000 460.350000 558.500000 461.650000 ;
      RECT 516.500000 460.350000 549.500000 461.650000 ;
      RECT 507.500000 460.350000 508.500000 461.650000 ;
      RECT 466.500000 460.350000 499.500000 461.650000 ;
      RECT 457.500000 460.350000 458.500000 461.650000 ;
      RECT 416.500000 460.350000 449.500000 461.650000 ;
      RECT 407.500000 460.350000 408.500000 461.650000 ;
      RECT 366.500000 460.350000 399.500000 461.650000 ;
      RECT 357.500000 460.350000 358.500000 461.650000 ;
      RECT 316.500000 460.350000 349.500000 461.650000 ;
      RECT 307.500000 460.350000 308.500000 461.650000 ;
      RECT 257.500000 460.350000 299.500000 462.350000 ;
      RECT 216.500000 460.350000 249.500000 461.650000 ;
      RECT 207.500000 460.350000 208.500000 461.650000 ;
      RECT 157.500000 460.350000 199.500000 462.350000 ;
      RECT 116.500000 460.350000 149.500000 461.650000 ;
      RECT 107.500000 460.350000 108.500000 461.650000 ;
      RECT 66.500000 460.350000 99.500000 461.650000 ;
      RECT 57.500000 460.350000 58.500000 461.650000 ;
      RECT 29.500000 460.350000 49.500000 461.650000 ;
      RECT 15.500000 460.350000 16.500000 461.650000 ;
      RECT 0.000000 460.350000 2.500000 463.650000 ;
      RECT 1139.000000 459.650000 1158.500000 460.350000 ;
      RECT 722.500000 459.650000 739.000000 460.350000 ;
      RECT 666.500000 459.650000 708.500000 460.350000 ;
      RECT 616.500000 459.650000 658.500000 460.350000 ;
      RECT 566.500000 459.650000 608.500000 460.350000 ;
      RECT 516.500000 459.650000 558.500000 460.350000 ;
      RECT 466.500000 459.650000 508.500000 460.350000 ;
      RECT 416.500000 459.650000 458.500000 460.350000 ;
      RECT 366.500000 459.650000 408.500000 460.350000 ;
      RECT 316.500000 459.650000 358.500000 460.350000 ;
      RECT 216.500000 459.650000 308.500000 460.350000 ;
      RECT 116.500000 459.650000 208.500000 460.350000 ;
      RECT 66.500000 459.650000 108.500000 460.350000 ;
      RECT 29.500000 459.650000 58.500000 460.350000 ;
      RECT 0.000000 459.650000 16.500000 460.350000 ;
      RECT 1166.500000 458.350000 1186.000000 461.650000 ;
      RECT 1157.500000 458.350000 1158.500000 459.650000 ;
      RECT 722.500000 458.350000 723.500000 459.650000 ;
      RECT 707.500000 458.350000 708.500000 459.650000 ;
      RECT 666.500000 458.350000 699.500000 459.650000 ;
      RECT 657.500000 458.350000 658.500000 459.650000 ;
      RECT 616.500000 458.350000 649.500000 459.650000 ;
      RECT 607.500000 458.350000 608.500000 459.650000 ;
      RECT 566.500000 458.350000 599.500000 459.650000 ;
      RECT 557.500000 458.350000 558.500000 459.650000 ;
      RECT 516.500000 458.350000 549.500000 459.650000 ;
      RECT 507.500000 458.350000 508.500000 459.650000 ;
      RECT 466.500000 458.350000 499.500000 459.650000 ;
      RECT 457.500000 458.350000 458.500000 459.650000 ;
      RECT 416.500000 458.350000 449.500000 459.650000 ;
      RECT 407.500000 458.350000 408.500000 459.650000 ;
      RECT 366.500000 458.350000 399.500000 459.650000 ;
      RECT 357.500000 458.350000 358.500000 459.650000 ;
      RECT 316.500000 458.350000 349.500000 459.650000 ;
      RECT 307.500000 458.350000 308.500000 459.650000 ;
      RECT 216.500000 458.350000 249.500000 459.650000 ;
      RECT 207.500000 458.350000 208.500000 459.650000 ;
      RECT 116.500000 458.350000 149.500000 459.650000 ;
      RECT 107.500000 458.350000 108.500000 459.650000 ;
      RECT 66.500000 458.350000 99.500000 459.650000 ;
      RECT 57.500000 458.350000 58.500000 459.650000 ;
      RECT 29.500000 458.350000 49.500000 459.650000 ;
      RECT 15.500000 458.350000 16.500000 459.650000 ;
      RECT 1157.500000 457.650000 1186.000000 458.350000 ;
      RECT 707.500000 457.650000 723.500000 458.350000 ;
      RECT 657.500000 457.650000 699.500000 458.350000 ;
      RECT 607.500000 457.650000 649.500000 458.350000 ;
      RECT 557.500000 457.650000 599.500000 458.350000 ;
      RECT 507.500000 457.650000 549.500000 458.350000 ;
      RECT 457.500000 457.650000 499.500000 458.350000 ;
      RECT 407.500000 457.650000 449.500000 458.350000 ;
      RECT 357.500000 457.650000 399.500000 458.350000 ;
      RECT 307.500000 457.650000 349.500000 458.350000 ;
      RECT 207.500000 457.650000 249.500000 458.350000 ;
      RECT 107.500000 457.650000 149.500000 458.350000 ;
      RECT 57.500000 457.650000 99.500000 458.350000 ;
      RECT 15.500000 457.650000 49.500000 458.350000 ;
      RECT 1157.500000 456.350000 1158.500000 457.650000 ;
      RECT 1139.000000 456.350000 1149.500000 459.650000 ;
      RECT 736.500000 456.350000 739.000000 459.650000 ;
      RECT 722.500000 456.350000 723.500000 457.650000 ;
      RECT 707.500000 456.350000 708.500000 457.650000 ;
      RECT 666.500000 456.350000 699.500000 457.650000 ;
      RECT 657.500000 456.350000 658.500000 457.650000 ;
      RECT 616.500000 456.350000 649.500000 457.650000 ;
      RECT 607.500000 456.350000 608.500000 457.650000 ;
      RECT 566.500000 456.350000 599.500000 457.650000 ;
      RECT 557.500000 456.350000 558.500000 457.650000 ;
      RECT 516.500000 456.350000 549.500000 457.650000 ;
      RECT 507.500000 456.350000 508.500000 457.650000 ;
      RECT 466.500000 456.350000 499.500000 457.650000 ;
      RECT 457.500000 456.350000 458.500000 457.650000 ;
      RECT 416.500000 456.350000 449.500000 457.650000 ;
      RECT 407.500000 456.350000 408.500000 457.650000 ;
      RECT 366.500000 456.350000 399.500000 457.650000 ;
      RECT 357.500000 456.350000 358.500000 457.650000 ;
      RECT 316.500000 456.350000 349.500000 457.650000 ;
      RECT 307.500000 456.350000 308.500000 457.650000 ;
      RECT 257.500000 456.350000 299.500000 459.650000 ;
      RECT 216.500000 456.350000 249.500000 457.650000 ;
      RECT 207.500000 456.350000 208.500000 457.650000 ;
      RECT 157.500000 456.350000 199.500000 459.650000 ;
      RECT 116.500000 456.350000 149.500000 457.650000 ;
      RECT 107.500000 456.350000 108.500000 457.650000 ;
      RECT 66.500000 456.350000 99.500000 457.650000 ;
      RECT 57.500000 456.350000 58.500000 457.650000 ;
      RECT 29.500000 456.350000 49.500000 457.650000 ;
      RECT 15.500000 456.350000 16.500000 457.650000 ;
      RECT 0.000000 456.350000 2.500000 459.650000 ;
      RECT 1139.000000 455.650000 1158.500000 456.350000 ;
      RECT 722.500000 455.650000 739.000000 456.350000 ;
      RECT 666.500000 455.650000 708.500000 456.350000 ;
      RECT 616.500000 455.650000 658.500000 456.350000 ;
      RECT 566.500000 455.650000 608.500000 456.350000 ;
      RECT 516.500000 455.650000 558.500000 456.350000 ;
      RECT 466.500000 455.650000 508.500000 456.350000 ;
      RECT 416.500000 455.650000 458.500000 456.350000 ;
      RECT 366.500000 455.650000 408.500000 456.350000 ;
      RECT 316.500000 455.650000 358.500000 456.350000 ;
      RECT 216.500000 455.650000 308.500000 456.350000 ;
      RECT 116.500000 455.650000 208.500000 456.350000 ;
      RECT 66.500000 455.650000 108.500000 456.350000 ;
      RECT 29.500000 455.650000 58.500000 456.350000 ;
      RECT 0.000000 455.650000 16.500000 456.350000 ;
      RECT 1166.500000 454.350000 1186.000000 457.650000 ;
      RECT 1157.500000 454.350000 1158.500000 455.650000 ;
      RECT 722.500000 454.350000 723.500000 455.650000 ;
      RECT 707.500000 454.350000 708.500000 455.650000 ;
      RECT 666.500000 454.350000 699.500000 455.650000 ;
      RECT 657.500000 454.350000 658.500000 455.650000 ;
      RECT 616.500000 454.350000 649.500000 455.650000 ;
      RECT 607.500000 454.350000 608.500000 455.650000 ;
      RECT 566.500000 454.350000 599.500000 455.650000 ;
      RECT 557.500000 454.350000 558.500000 455.650000 ;
      RECT 516.500000 454.350000 549.500000 455.650000 ;
      RECT 507.500000 454.350000 508.500000 455.650000 ;
      RECT 466.500000 454.350000 499.500000 455.650000 ;
      RECT 457.500000 454.350000 458.500000 455.650000 ;
      RECT 416.500000 454.350000 449.500000 455.650000 ;
      RECT 407.500000 454.350000 408.500000 455.650000 ;
      RECT 366.500000 454.350000 399.500000 455.650000 ;
      RECT 357.500000 454.350000 358.500000 455.650000 ;
      RECT 316.500000 454.350000 349.500000 455.650000 ;
      RECT 307.500000 454.350000 308.500000 455.650000 ;
      RECT 216.500000 454.350000 249.500000 455.650000 ;
      RECT 207.500000 454.350000 208.500000 455.650000 ;
      RECT 116.500000 454.350000 149.500000 455.650000 ;
      RECT 107.500000 454.350000 108.500000 455.650000 ;
      RECT 66.500000 454.350000 99.500000 455.650000 ;
      RECT 57.500000 454.350000 58.500000 455.650000 ;
      RECT 29.500000 454.350000 49.500000 455.650000 ;
      RECT 15.500000 454.350000 16.500000 455.650000 ;
      RECT 1157.500000 453.650000 1186.000000 454.350000 ;
      RECT 707.500000 453.650000 723.500000 454.350000 ;
      RECT 657.500000 453.650000 699.500000 454.350000 ;
      RECT 607.500000 453.650000 649.500000 454.350000 ;
      RECT 557.500000 453.650000 599.500000 454.350000 ;
      RECT 507.500000 453.650000 549.500000 454.350000 ;
      RECT 457.500000 453.650000 499.500000 454.350000 ;
      RECT 407.500000 453.650000 449.500000 454.350000 ;
      RECT 357.500000 453.650000 399.500000 454.350000 ;
      RECT 307.500000 453.650000 349.500000 454.350000 ;
      RECT 207.500000 453.650000 249.500000 454.350000 ;
      RECT 107.500000 453.650000 149.500000 454.350000 ;
      RECT 57.500000 453.650000 99.500000 454.350000 ;
      RECT 15.500000 453.650000 49.500000 454.350000 ;
      RECT 1157.500000 452.350000 1158.500000 453.650000 ;
      RECT 1139.000000 452.350000 1149.500000 455.650000 ;
      RECT 736.500000 452.350000 739.000000 455.650000 ;
      RECT 722.500000 452.350000 723.500000 453.650000 ;
      RECT 707.500000 452.350000 708.500000 453.650000 ;
      RECT 666.500000 452.350000 699.500000 453.650000 ;
      RECT 657.500000 452.350000 658.500000 453.650000 ;
      RECT 616.500000 452.350000 649.500000 453.650000 ;
      RECT 607.500000 452.350000 608.500000 453.650000 ;
      RECT 566.500000 452.350000 599.500000 453.650000 ;
      RECT 557.500000 452.350000 558.500000 453.650000 ;
      RECT 516.500000 452.350000 549.500000 453.650000 ;
      RECT 507.500000 452.350000 508.500000 453.650000 ;
      RECT 466.500000 452.350000 499.500000 453.650000 ;
      RECT 457.500000 452.350000 458.500000 453.650000 ;
      RECT 416.500000 452.350000 449.500000 453.650000 ;
      RECT 407.500000 452.350000 408.500000 453.650000 ;
      RECT 366.500000 452.350000 399.500000 453.650000 ;
      RECT 357.500000 452.350000 358.500000 453.650000 ;
      RECT 316.500000 452.350000 349.500000 453.650000 ;
      RECT 307.500000 452.350000 308.500000 453.650000 ;
      RECT 257.500000 452.350000 299.500000 455.650000 ;
      RECT 216.500000 452.350000 249.500000 453.650000 ;
      RECT 207.500000 452.350000 208.500000 453.650000 ;
      RECT 157.500000 452.350000 199.500000 455.650000 ;
      RECT 116.500000 452.350000 149.500000 453.650000 ;
      RECT 107.500000 452.350000 108.500000 453.650000 ;
      RECT 66.500000 452.350000 99.500000 453.650000 ;
      RECT 57.500000 452.350000 58.500000 453.650000 ;
      RECT 29.500000 452.350000 49.500000 453.650000 ;
      RECT 15.500000 452.350000 16.500000 453.650000 ;
      RECT 0.000000 452.350000 2.500000 455.650000 ;
      RECT 1139.000000 451.650000 1158.500000 452.350000 ;
      RECT 722.500000 451.650000 739.000000 452.350000 ;
      RECT 666.500000 451.650000 708.500000 452.350000 ;
      RECT 616.500000 451.650000 658.500000 452.350000 ;
      RECT 566.500000 451.650000 608.500000 452.350000 ;
      RECT 516.500000 451.650000 558.500000 452.350000 ;
      RECT 466.500000 451.650000 508.500000 452.350000 ;
      RECT 416.500000 451.650000 458.500000 452.350000 ;
      RECT 366.500000 451.650000 408.500000 452.350000 ;
      RECT 316.500000 451.650000 358.500000 452.350000 ;
      RECT 216.500000 451.650000 308.500000 452.350000 ;
      RECT 116.500000 451.650000 208.500000 452.350000 ;
      RECT 66.500000 451.650000 108.500000 452.350000 ;
      RECT 29.500000 451.650000 58.500000 452.350000 ;
      RECT 0.000000 451.650000 16.500000 452.350000 ;
      RECT 1166.500000 450.350000 1186.000000 453.650000 ;
      RECT 1157.500000 450.350000 1158.500000 451.650000 ;
      RECT 722.500000 450.350000 723.500000 451.650000 ;
      RECT 707.500000 450.350000 708.500000 451.650000 ;
      RECT 666.500000 450.350000 699.500000 451.650000 ;
      RECT 657.500000 450.350000 658.500000 451.650000 ;
      RECT 616.500000 450.350000 649.500000 451.650000 ;
      RECT 607.500000 450.350000 608.500000 451.650000 ;
      RECT 566.500000 450.350000 599.500000 451.650000 ;
      RECT 557.500000 450.350000 558.500000 451.650000 ;
      RECT 516.500000 450.350000 549.500000 451.650000 ;
      RECT 507.500000 450.350000 508.500000 451.650000 ;
      RECT 466.500000 450.350000 499.500000 451.650000 ;
      RECT 457.500000 450.350000 458.500000 451.650000 ;
      RECT 416.500000 450.350000 449.500000 451.650000 ;
      RECT 407.500000 450.350000 408.500000 451.650000 ;
      RECT 366.500000 450.350000 399.500000 451.650000 ;
      RECT 357.500000 450.350000 358.500000 451.650000 ;
      RECT 316.500000 450.350000 349.500000 451.650000 ;
      RECT 307.500000 450.350000 308.500000 451.650000 ;
      RECT 216.500000 450.350000 299.500000 451.650000 ;
      RECT 207.500000 450.350000 208.500000 451.650000 ;
      RECT 116.500000 450.350000 199.500000 451.650000 ;
      RECT 107.500000 450.350000 108.500000 451.650000 ;
      RECT 66.500000 450.350000 99.500000 451.650000 ;
      RECT 57.500000 450.350000 58.500000 451.650000 ;
      RECT 29.500000 450.350000 49.500000 451.650000 ;
      RECT 15.500000 450.350000 16.500000 451.650000 ;
      RECT 1157.500000 449.650000 1186.000000 450.350000 ;
      RECT 707.500000 449.650000 723.500000 450.350000 ;
      RECT 657.500000 449.650000 699.500000 450.350000 ;
      RECT 607.500000 449.650000 649.500000 450.350000 ;
      RECT 557.500000 449.650000 599.500000 450.350000 ;
      RECT 507.500000 449.650000 549.500000 450.350000 ;
      RECT 457.500000 449.650000 499.500000 450.350000 ;
      RECT 407.500000 449.650000 449.500000 450.350000 ;
      RECT 357.500000 449.650000 399.500000 450.350000 ;
      RECT 307.500000 449.650000 349.500000 450.350000 ;
      RECT 207.500000 449.650000 299.500000 450.350000 ;
      RECT 107.500000 449.650000 199.500000 450.350000 ;
      RECT 57.500000 449.650000 99.500000 450.350000 ;
      RECT 15.500000 449.650000 49.500000 450.350000 ;
      RECT 1157.500000 448.350000 1158.500000 449.650000 ;
      RECT 1139.000000 448.350000 1149.500000 451.650000 ;
      RECT 736.500000 448.350000 739.000000 451.650000 ;
      RECT 722.500000 448.350000 723.500000 449.650000 ;
      RECT 707.500000 448.350000 708.500000 449.650000 ;
      RECT 666.500000 448.350000 699.500000 449.650000 ;
      RECT 657.500000 448.350000 658.500000 449.650000 ;
      RECT 616.500000 448.350000 649.500000 449.650000 ;
      RECT 607.500000 448.350000 608.500000 449.650000 ;
      RECT 566.500000 448.350000 599.500000 449.650000 ;
      RECT 557.500000 448.350000 558.500000 449.650000 ;
      RECT 516.500000 448.350000 549.500000 449.650000 ;
      RECT 507.500000 448.350000 508.500000 449.650000 ;
      RECT 466.500000 448.350000 499.500000 449.650000 ;
      RECT 457.500000 448.350000 458.500000 449.650000 ;
      RECT 416.500000 448.350000 449.500000 449.650000 ;
      RECT 407.500000 448.350000 408.500000 449.650000 ;
      RECT 366.500000 448.350000 399.500000 449.650000 ;
      RECT 357.500000 448.350000 358.500000 449.650000 ;
      RECT 316.500000 448.350000 349.500000 449.650000 ;
      RECT 307.500000 448.350000 308.500000 449.650000 ;
      RECT 216.500000 448.350000 299.500000 449.650000 ;
      RECT 207.500000 448.350000 208.500000 449.650000 ;
      RECT 116.500000 448.350000 199.500000 449.650000 ;
      RECT 107.500000 448.350000 108.500000 449.650000 ;
      RECT 66.500000 448.350000 99.500000 449.650000 ;
      RECT 57.500000 448.350000 58.500000 449.650000 ;
      RECT 29.500000 448.350000 49.500000 449.650000 ;
      RECT 15.500000 448.350000 16.500000 449.650000 ;
      RECT 0.000000 448.350000 2.500000 451.650000 ;
      RECT 1139.000000 447.650000 1158.500000 448.350000 ;
      RECT 722.500000 447.650000 739.000000 448.350000 ;
      RECT 666.500000 447.650000 708.500000 448.350000 ;
      RECT 616.500000 447.650000 658.500000 448.350000 ;
      RECT 566.500000 447.650000 608.500000 448.350000 ;
      RECT 516.500000 447.650000 558.500000 448.350000 ;
      RECT 466.500000 447.650000 508.500000 448.350000 ;
      RECT 416.500000 447.650000 458.500000 448.350000 ;
      RECT 366.500000 447.650000 408.500000 448.350000 ;
      RECT 316.500000 447.650000 358.500000 448.350000 ;
      RECT 216.500000 447.650000 308.500000 448.350000 ;
      RECT 116.500000 447.650000 208.500000 448.350000 ;
      RECT 66.500000 447.650000 108.500000 448.350000 ;
      RECT 29.500000 447.650000 58.500000 448.350000 ;
      RECT 0.000000 447.650000 16.500000 448.350000 ;
      RECT 1166.500000 446.350000 1186.000000 449.650000 ;
      RECT 1157.500000 446.350000 1158.500000 447.650000 ;
      RECT 722.500000 446.350000 723.500000 447.650000 ;
      RECT 707.500000 446.350000 708.500000 447.650000 ;
      RECT 666.500000 446.350000 699.500000 447.650000 ;
      RECT 657.500000 446.350000 658.500000 447.650000 ;
      RECT 616.500000 446.350000 649.500000 447.650000 ;
      RECT 607.500000 446.350000 608.500000 447.650000 ;
      RECT 566.500000 446.350000 599.500000 447.650000 ;
      RECT 557.500000 446.350000 558.500000 447.650000 ;
      RECT 516.500000 446.350000 549.500000 447.650000 ;
      RECT 507.500000 446.350000 508.500000 447.650000 ;
      RECT 466.500000 446.350000 499.500000 447.650000 ;
      RECT 457.500000 446.350000 458.500000 447.650000 ;
      RECT 416.500000 446.350000 449.500000 447.650000 ;
      RECT 407.500000 446.350000 408.500000 447.650000 ;
      RECT 366.500000 446.350000 399.500000 447.650000 ;
      RECT 357.500000 446.350000 358.500000 447.650000 ;
      RECT 316.500000 446.350000 349.500000 447.650000 ;
      RECT 307.500000 446.350000 308.500000 447.650000 ;
      RECT 216.500000 446.350000 299.500000 447.650000 ;
      RECT 207.500000 446.350000 208.500000 447.650000 ;
      RECT 116.500000 446.350000 199.500000 447.650000 ;
      RECT 107.500000 446.350000 108.500000 447.650000 ;
      RECT 66.500000 446.350000 99.500000 447.650000 ;
      RECT 57.500000 446.350000 58.500000 447.650000 ;
      RECT 29.500000 446.350000 49.500000 447.650000 ;
      RECT 15.500000 446.350000 16.500000 447.650000 ;
      RECT 1139.000000 446.000000 1149.500000 447.650000 ;
      RECT 736.500000 446.000000 739.000000 447.650000 ;
      RECT 1157.500000 445.650000 1186.000000 446.350000 ;
      RECT 1060.750000 445.650000 1149.500000 446.000000 ;
      RECT 999.630000 445.650000 1009.115000 446.000000 ;
      RECT 876.205000 445.650000 996.530000 446.000000 ;
      RECT 736.500000 445.650000 868.305000 446.000000 ;
      RECT 707.500000 445.650000 723.500000 446.350000 ;
      RECT 657.500000 445.650000 699.500000 446.350000 ;
      RECT 607.500000 445.650000 649.500000 446.350000 ;
      RECT 557.500000 445.650000 599.500000 446.350000 ;
      RECT 507.500000 445.650000 549.500000 446.350000 ;
      RECT 457.500000 445.650000 499.500000 446.350000 ;
      RECT 407.500000 445.650000 449.500000 446.350000 ;
      RECT 357.500000 445.650000 399.500000 446.350000 ;
      RECT 307.500000 445.650000 349.500000 446.350000 ;
      RECT 207.500000 445.650000 299.500000 446.350000 ;
      RECT 107.500000 445.650000 199.500000 446.350000 ;
      RECT 57.500000 445.650000 99.500000 446.350000 ;
      RECT 15.500000 445.650000 49.500000 446.350000 ;
      RECT 1157.500000 444.350000 1158.500000 445.650000 ;
      RECT 1116.500000 444.350000 1149.500000 445.650000 ;
      RECT 736.500000 444.350000 758.500000 445.650000 ;
      RECT 722.500000 444.350000 723.500000 445.650000 ;
      RECT 707.500000 444.350000 708.500000 445.650000 ;
      RECT 666.500000 444.350000 699.500000 445.650000 ;
      RECT 657.500000 444.350000 658.500000 445.650000 ;
      RECT 616.500000 444.350000 649.500000 445.650000 ;
      RECT 607.500000 444.350000 608.500000 445.650000 ;
      RECT 566.500000 444.350000 599.500000 445.650000 ;
      RECT 557.500000 444.350000 558.500000 445.650000 ;
      RECT 516.500000 444.350000 549.500000 445.650000 ;
      RECT 507.500000 444.350000 508.500000 445.650000 ;
      RECT 466.500000 444.350000 499.500000 445.650000 ;
      RECT 457.500000 444.350000 458.500000 445.650000 ;
      RECT 416.500000 444.350000 449.500000 445.650000 ;
      RECT 407.500000 444.350000 408.500000 445.650000 ;
      RECT 366.500000 444.350000 399.500000 445.650000 ;
      RECT 357.500000 444.350000 358.500000 445.650000 ;
      RECT 316.500000 444.350000 349.500000 445.650000 ;
      RECT 307.500000 444.350000 308.500000 445.650000 ;
      RECT 216.500000 444.350000 299.500000 445.650000 ;
      RECT 207.500000 444.350000 208.500000 445.650000 ;
      RECT 116.500000 444.350000 199.500000 445.650000 ;
      RECT 107.500000 444.350000 108.500000 445.650000 ;
      RECT 66.500000 444.350000 99.500000 445.650000 ;
      RECT 57.500000 444.350000 58.500000 445.650000 ;
      RECT 29.500000 444.350000 49.500000 445.650000 ;
      RECT 15.500000 444.350000 16.500000 445.650000 ;
      RECT 0.000000 444.350000 2.500000 447.650000 ;
      RECT 1029.110000 443.980000 1040.755000 446.000000 ;
      RECT 999.630000 443.980000 1008.500000 445.650000 ;
      RECT 966.500000 443.980000 996.530000 445.650000 ;
      RECT 876.205000 443.980000 908.500000 445.650000 ;
      RECT 866.500000 443.980000 868.305000 445.650000 ;
      RECT 1166.500000 443.650000 1186.000000 445.650000 ;
      RECT 1116.500000 443.650000 1158.500000 444.350000 ;
      RECT 1066.500000 443.650000 1108.500000 445.650000 ;
      RECT 1016.500000 443.650000 1058.500000 443.980000 ;
      RECT 966.500000 443.650000 1008.500000 443.980000 ;
      RECT 916.500000 443.650000 958.500000 445.650000 ;
      RECT 866.500000 443.650000 908.500000 443.980000 ;
      RECT 816.500000 443.650000 858.500000 445.650000 ;
      RECT 766.500000 443.650000 808.500000 445.650000 ;
      RECT 722.500000 443.650000 758.500000 444.350000 ;
      RECT 666.500000 443.650000 708.500000 444.350000 ;
      RECT 616.500000 443.650000 658.500000 444.350000 ;
      RECT 566.500000 443.650000 608.500000 444.350000 ;
      RECT 516.500000 443.650000 558.500000 444.350000 ;
      RECT 466.500000 443.650000 508.500000 444.350000 ;
      RECT 416.500000 443.650000 458.500000 444.350000 ;
      RECT 366.500000 443.650000 408.500000 444.350000 ;
      RECT 316.500000 443.650000 358.500000 444.350000 ;
      RECT 216.500000 443.650000 308.500000 444.350000 ;
      RECT 116.500000 443.650000 208.500000 444.350000 ;
      RECT 66.500000 443.650000 108.500000 444.350000 ;
      RECT 29.500000 443.650000 58.500000 444.350000 ;
      RECT 0.000000 443.650000 16.500000 444.350000 ;
      RECT 1166.500000 442.350000 1170.500000 443.650000 ;
      RECT 1157.500000 442.350000 1158.500000 443.650000 ;
      RECT 1116.500000 442.350000 1149.500000 443.650000 ;
      RECT 1107.500000 442.350000 1108.500000 443.650000 ;
      RECT 1066.500000 442.350000 1099.500000 443.650000 ;
      RECT 1057.500000 442.350000 1058.500000 443.650000 ;
      RECT 1016.500000 442.350000 1049.500000 443.650000 ;
      RECT 1007.500000 442.350000 1008.500000 443.650000 ;
      RECT 966.500000 442.350000 999.500000 443.650000 ;
      RECT 957.500000 442.350000 958.500000 443.650000 ;
      RECT 916.500000 442.350000 949.500000 443.650000 ;
      RECT 907.500000 442.350000 908.500000 443.650000 ;
      RECT 866.500000 442.350000 899.500000 443.650000 ;
      RECT 857.500000 442.350000 858.500000 443.650000 ;
      RECT 816.500000 442.350000 849.500000 443.650000 ;
      RECT 807.500000 442.350000 808.500000 443.650000 ;
      RECT 766.500000 442.350000 799.500000 443.650000 ;
      RECT 757.500000 442.350000 758.500000 443.650000 ;
      RECT 722.500000 442.350000 723.500000 443.650000 ;
      RECT 707.500000 442.350000 708.500000 443.650000 ;
      RECT 666.500000 442.350000 699.500000 443.650000 ;
      RECT 657.500000 442.350000 658.500000 443.650000 ;
      RECT 616.500000 442.350000 649.500000 443.650000 ;
      RECT 607.500000 442.350000 608.500000 443.650000 ;
      RECT 566.500000 442.350000 599.500000 443.650000 ;
      RECT 557.500000 442.350000 558.500000 443.650000 ;
      RECT 516.500000 442.350000 549.500000 443.650000 ;
      RECT 507.500000 442.350000 508.500000 443.650000 ;
      RECT 466.500000 442.350000 499.500000 443.650000 ;
      RECT 457.500000 442.350000 458.500000 443.650000 ;
      RECT 416.500000 442.350000 449.500000 443.650000 ;
      RECT 407.500000 442.350000 408.500000 443.650000 ;
      RECT 366.500000 442.350000 399.500000 443.650000 ;
      RECT 357.500000 442.350000 358.500000 443.650000 ;
      RECT 316.500000 442.350000 349.500000 443.650000 ;
      RECT 307.500000 442.350000 308.500000 443.650000 ;
      RECT 216.500000 442.350000 299.500000 443.650000 ;
      RECT 207.500000 442.350000 208.500000 443.650000 ;
      RECT 116.500000 442.350000 199.500000 443.650000 ;
      RECT 107.500000 442.350000 108.500000 443.650000 ;
      RECT 66.500000 442.350000 99.500000 443.650000 ;
      RECT 57.500000 442.350000 58.500000 443.650000 ;
      RECT 29.500000 442.350000 49.500000 443.650000 ;
      RECT 15.500000 442.350000 16.500000 443.650000 ;
      RECT 1157.500000 441.650000 1170.500000 442.350000 ;
      RECT 1107.500000 441.650000 1149.500000 442.350000 ;
      RECT 1057.500000 441.650000 1099.500000 442.350000 ;
      RECT 1007.500000 441.650000 1049.500000 442.350000 ;
      RECT 957.500000 441.650000 999.500000 442.350000 ;
      RECT 907.500000 441.650000 949.500000 442.350000 ;
      RECT 857.500000 441.650000 899.500000 442.350000 ;
      RECT 807.500000 441.650000 849.500000 442.350000 ;
      RECT 757.500000 441.650000 799.500000 442.350000 ;
      RECT 707.500000 441.650000 723.500000 442.350000 ;
      RECT 657.500000 441.650000 699.500000 442.350000 ;
      RECT 607.500000 441.650000 649.500000 442.350000 ;
      RECT 557.500000 441.650000 599.500000 442.350000 ;
      RECT 507.500000 441.650000 549.500000 442.350000 ;
      RECT 457.500000 441.650000 499.500000 442.350000 ;
      RECT 407.500000 441.650000 449.500000 442.350000 ;
      RECT 357.500000 441.650000 399.500000 442.350000 ;
      RECT 307.500000 441.650000 349.500000 442.350000 ;
      RECT 207.500000 441.650000 299.500000 442.350000 ;
      RECT 107.500000 441.650000 199.500000 442.350000 ;
      RECT 57.500000 441.650000 99.500000 442.350000 ;
      RECT 15.500000 441.650000 49.500000 442.350000 ;
      RECT 1183.500000 440.350000 1186.000000 443.650000 ;
      RECT 1166.500000 440.350000 1170.500000 441.650000 ;
      RECT 1157.500000 440.350000 1158.500000 441.650000 ;
      RECT 1116.500000 440.350000 1149.500000 441.650000 ;
      RECT 1107.500000 440.350000 1108.500000 441.650000 ;
      RECT 1066.500000 440.350000 1099.500000 441.650000 ;
      RECT 1057.500000 440.350000 1058.500000 441.650000 ;
      RECT 1016.500000 440.350000 1049.500000 441.650000 ;
      RECT 1007.500000 440.350000 1008.500000 441.650000 ;
      RECT 966.500000 440.350000 999.500000 441.650000 ;
      RECT 957.500000 440.350000 958.500000 441.650000 ;
      RECT 916.500000 440.350000 949.500000 441.650000 ;
      RECT 907.500000 440.350000 908.500000 441.650000 ;
      RECT 866.500000 440.350000 899.500000 441.650000 ;
      RECT 857.500000 440.350000 858.500000 441.650000 ;
      RECT 816.500000 440.350000 849.500000 441.650000 ;
      RECT 807.500000 440.350000 808.500000 441.650000 ;
      RECT 766.500000 440.350000 799.500000 441.650000 ;
      RECT 757.500000 440.350000 758.500000 441.650000 ;
      RECT 736.500000 440.350000 749.500000 443.650000 ;
      RECT 722.500000 440.350000 723.500000 441.650000 ;
      RECT 707.500000 440.350000 708.500000 441.650000 ;
      RECT 666.500000 440.350000 699.500000 441.650000 ;
      RECT 657.500000 440.350000 658.500000 441.650000 ;
      RECT 616.500000 440.350000 649.500000 441.650000 ;
      RECT 607.500000 440.350000 608.500000 441.650000 ;
      RECT 566.500000 440.350000 599.500000 441.650000 ;
      RECT 557.500000 440.350000 558.500000 441.650000 ;
      RECT 516.500000 440.350000 549.500000 441.650000 ;
      RECT 507.500000 440.350000 508.500000 441.650000 ;
      RECT 466.500000 440.350000 499.500000 441.650000 ;
      RECT 457.500000 440.350000 458.500000 441.650000 ;
      RECT 416.500000 440.350000 449.500000 441.650000 ;
      RECT 407.500000 440.350000 408.500000 441.650000 ;
      RECT 366.500000 440.350000 399.500000 441.650000 ;
      RECT 357.500000 440.350000 358.500000 441.650000 ;
      RECT 316.500000 440.350000 349.500000 441.650000 ;
      RECT 307.500000 440.350000 308.500000 441.650000 ;
      RECT 216.500000 440.350000 299.500000 441.650000 ;
      RECT 207.500000 440.350000 208.500000 441.650000 ;
      RECT 116.500000 440.350000 199.500000 441.650000 ;
      RECT 107.500000 440.350000 108.500000 441.650000 ;
      RECT 66.500000 440.350000 99.500000 441.650000 ;
      RECT 57.500000 440.350000 58.500000 441.650000 ;
      RECT 29.500000 440.350000 49.500000 441.650000 ;
      RECT 15.500000 440.350000 16.500000 441.650000 ;
      RECT 0.000000 440.350000 2.500000 443.650000 ;
      RECT 1166.500000 439.650000 1186.000000 440.350000 ;
      RECT 1116.500000 439.650000 1158.500000 440.350000 ;
      RECT 1066.500000 439.650000 1108.500000 440.350000 ;
      RECT 1016.500000 439.650000 1058.500000 440.350000 ;
      RECT 966.500000 439.650000 1008.500000 440.350000 ;
      RECT 916.500000 439.650000 958.500000 440.350000 ;
      RECT 866.500000 439.650000 908.500000 440.350000 ;
      RECT 816.500000 439.650000 858.500000 440.350000 ;
      RECT 766.500000 439.650000 808.500000 440.350000 ;
      RECT 722.500000 439.650000 758.500000 440.350000 ;
      RECT 666.500000 439.650000 708.500000 440.350000 ;
      RECT 616.500000 439.650000 658.500000 440.350000 ;
      RECT 566.500000 439.650000 608.500000 440.350000 ;
      RECT 516.500000 439.650000 558.500000 440.350000 ;
      RECT 466.500000 439.650000 508.500000 440.350000 ;
      RECT 416.500000 439.650000 458.500000 440.350000 ;
      RECT 366.500000 439.650000 408.500000 440.350000 ;
      RECT 316.500000 439.650000 358.500000 440.350000 ;
      RECT 216.500000 439.650000 308.500000 440.350000 ;
      RECT 116.500000 439.650000 208.500000 440.350000 ;
      RECT 66.500000 439.650000 108.500000 440.350000 ;
      RECT 29.500000 439.650000 58.500000 440.350000 ;
      RECT 0.000000 439.650000 16.500000 440.350000 ;
      RECT 1166.500000 438.350000 1170.500000 439.650000 ;
      RECT 1157.500000 438.350000 1158.500000 439.650000 ;
      RECT 1116.500000 438.350000 1149.500000 439.650000 ;
      RECT 1107.500000 438.350000 1108.500000 439.650000 ;
      RECT 1066.500000 438.350000 1099.500000 439.650000 ;
      RECT 1057.500000 438.350000 1058.500000 439.650000 ;
      RECT 1016.500000 438.350000 1049.500000 439.650000 ;
      RECT 1007.500000 438.350000 1008.500000 439.650000 ;
      RECT 966.500000 438.350000 999.500000 439.650000 ;
      RECT 957.500000 438.350000 958.500000 439.650000 ;
      RECT 916.500000 438.350000 949.500000 439.650000 ;
      RECT 907.500000 438.350000 908.500000 439.650000 ;
      RECT 866.500000 438.350000 899.500000 439.650000 ;
      RECT 857.500000 438.350000 858.500000 439.650000 ;
      RECT 816.500000 438.350000 849.500000 439.650000 ;
      RECT 807.500000 438.350000 808.500000 439.650000 ;
      RECT 766.500000 438.350000 799.500000 439.650000 ;
      RECT 757.500000 438.350000 758.500000 439.650000 ;
      RECT 722.500000 438.350000 723.500000 439.650000 ;
      RECT 707.500000 438.350000 708.500000 439.650000 ;
      RECT 666.500000 438.350000 699.500000 439.650000 ;
      RECT 657.500000 438.350000 658.500000 439.650000 ;
      RECT 616.500000 438.350000 649.500000 439.650000 ;
      RECT 607.500000 438.350000 608.500000 439.650000 ;
      RECT 566.500000 438.350000 599.500000 439.650000 ;
      RECT 557.500000 438.350000 558.500000 439.650000 ;
      RECT 516.500000 438.350000 549.500000 439.650000 ;
      RECT 507.500000 438.350000 508.500000 439.650000 ;
      RECT 466.500000 438.350000 499.500000 439.650000 ;
      RECT 457.500000 438.350000 458.500000 439.650000 ;
      RECT 416.500000 438.350000 449.500000 439.650000 ;
      RECT 407.500000 438.350000 408.500000 439.650000 ;
      RECT 366.500000 438.350000 399.500000 439.650000 ;
      RECT 357.500000 438.350000 358.500000 439.650000 ;
      RECT 316.500000 438.350000 349.500000 439.650000 ;
      RECT 307.500000 438.350000 308.500000 439.650000 ;
      RECT 216.500000 438.350000 299.500000 439.650000 ;
      RECT 207.500000 438.350000 208.500000 439.650000 ;
      RECT 116.500000 438.350000 199.500000 439.650000 ;
      RECT 107.500000 438.350000 108.500000 439.650000 ;
      RECT 66.500000 438.350000 99.500000 439.650000 ;
      RECT 57.500000 438.350000 58.500000 439.650000 ;
      RECT 29.500000 438.350000 49.500000 439.650000 ;
      RECT 15.500000 438.350000 16.500000 439.650000 ;
      RECT 1157.500000 437.650000 1170.500000 438.350000 ;
      RECT 1107.500000 437.650000 1149.500000 438.350000 ;
      RECT 1057.500000 437.650000 1099.500000 438.350000 ;
      RECT 1007.500000 437.650000 1049.500000 438.350000 ;
      RECT 957.500000 437.650000 999.500000 438.350000 ;
      RECT 907.500000 437.650000 949.500000 438.350000 ;
      RECT 857.500000 437.650000 899.500000 438.350000 ;
      RECT 807.500000 437.650000 849.500000 438.350000 ;
      RECT 757.500000 437.650000 799.500000 438.350000 ;
      RECT 707.500000 437.650000 723.500000 438.350000 ;
      RECT 657.500000 437.650000 699.500000 438.350000 ;
      RECT 607.500000 437.650000 649.500000 438.350000 ;
      RECT 557.500000 437.650000 599.500000 438.350000 ;
      RECT 507.500000 437.650000 549.500000 438.350000 ;
      RECT 457.500000 437.650000 499.500000 438.350000 ;
      RECT 407.500000 437.650000 449.500000 438.350000 ;
      RECT 357.500000 437.650000 399.500000 438.350000 ;
      RECT 307.500000 437.650000 349.500000 438.350000 ;
      RECT 207.500000 437.650000 299.500000 438.350000 ;
      RECT 107.500000 437.650000 199.500000 438.350000 ;
      RECT 57.500000 437.650000 99.500000 438.350000 ;
      RECT 15.500000 437.650000 49.500000 438.350000 ;
      RECT 1183.500000 436.350000 1186.000000 439.650000 ;
      RECT 1166.500000 436.350000 1170.500000 437.650000 ;
      RECT 1157.500000 436.350000 1158.500000 437.650000 ;
      RECT 1116.500000 436.350000 1149.500000 437.650000 ;
      RECT 1107.500000 436.350000 1108.500000 437.650000 ;
      RECT 1066.500000 436.350000 1099.500000 437.650000 ;
      RECT 1057.500000 436.350000 1058.500000 437.650000 ;
      RECT 1016.500000 436.350000 1049.500000 437.650000 ;
      RECT 1007.500000 436.350000 1008.500000 437.650000 ;
      RECT 966.500000 436.350000 999.500000 437.650000 ;
      RECT 957.500000 436.350000 958.500000 437.650000 ;
      RECT 916.500000 436.350000 949.500000 437.650000 ;
      RECT 907.500000 436.350000 908.500000 437.650000 ;
      RECT 866.500000 436.350000 899.500000 437.650000 ;
      RECT 857.500000 436.350000 858.500000 437.650000 ;
      RECT 816.500000 436.350000 849.500000 437.650000 ;
      RECT 807.500000 436.350000 808.500000 437.650000 ;
      RECT 766.500000 436.350000 799.500000 437.650000 ;
      RECT 757.500000 436.350000 758.500000 437.650000 ;
      RECT 736.500000 436.350000 749.500000 439.650000 ;
      RECT 722.500000 436.350000 723.500000 437.650000 ;
      RECT 707.500000 436.350000 708.500000 437.650000 ;
      RECT 666.500000 436.350000 699.500000 437.650000 ;
      RECT 657.500000 436.350000 658.500000 437.650000 ;
      RECT 616.500000 436.350000 649.500000 437.650000 ;
      RECT 607.500000 436.350000 608.500000 437.650000 ;
      RECT 566.500000 436.350000 599.500000 437.650000 ;
      RECT 557.500000 436.350000 558.500000 437.650000 ;
      RECT 516.500000 436.350000 549.500000 437.650000 ;
      RECT 507.500000 436.350000 508.500000 437.650000 ;
      RECT 466.500000 436.350000 499.500000 437.650000 ;
      RECT 457.500000 436.350000 458.500000 437.650000 ;
      RECT 416.500000 436.350000 449.500000 437.650000 ;
      RECT 407.500000 436.350000 408.500000 437.650000 ;
      RECT 366.500000 436.350000 399.500000 437.650000 ;
      RECT 357.500000 436.350000 358.500000 437.650000 ;
      RECT 316.500000 436.350000 349.500000 437.650000 ;
      RECT 307.500000 436.350000 308.500000 437.650000 ;
      RECT 216.500000 436.350000 299.500000 437.650000 ;
      RECT 207.500000 436.350000 208.500000 437.650000 ;
      RECT 116.500000 436.350000 199.500000 437.650000 ;
      RECT 107.500000 436.350000 108.500000 437.650000 ;
      RECT 66.500000 436.350000 99.500000 437.650000 ;
      RECT 57.500000 436.350000 58.500000 437.650000 ;
      RECT 29.500000 436.350000 49.500000 437.650000 ;
      RECT 15.500000 436.350000 16.500000 437.650000 ;
      RECT 0.000000 436.350000 2.500000 439.650000 ;
      RECT 1166.500000 435.650000 1186.000000 436.350000 ;
      RECT 1116.500000 435.650000 1158.500000 436.350000 ;
      RECT 1066.500000 435.650000 1108.500000 436.350000 ;
      RECT 1016.500000 435.650000 1058.500000 436.350000 ;
      RECT 966.500000 435.650000 1008.500000 436.350000 ;
      RECT 916.500000 435.650000 958.500000 436.350000 ;
      RECT 866.500000 435.650000 908.500000 436.350000 ;
      RECT 816.500000 435.650000 858.500000 436.350000 ;
      RECT 766.500000 435.650000 808.500000 436.350000 ;
      RECT 722.500000 435.650000 758.500000 436.350000 ;
      RECT 666.500000 435.650000 708.500000 436.350000 ;
      RECT 616.500000 435.650000 658.500000 436.350000 ;
      RECT 566.500000 435.650000 608.500000 436.350000 ;
      RECT 516.500000 435.650000 558.500000 436.350000 ;
      RECT 466.500000 435.650000 508.500000 436.350000 ;
      RECT 416.500000 435.650000 458.500000 436.350000 ;
      RECT 366.500000 435.650000 408.500000 436.350000 ;
      RECT 316.500000 435.650000 358.500000 436.350000 ;
      RECT 216.500000 435.650000 308.500000 436.350000 ;
      RECT 116.500000 435.650000 208.500000 436.350000 ;
      RECT 66.500000 435.650000 108.500000 436.350000 ;
      RECT 29.500000 435.650000 58.500000 436.350000 ;
      RECT 0.000000 435.650000 16.500000 436.350000 ;
      RECT 1166.500000 434.350000 1170.500000 435.650000 ;
      RECT 1157.500000 434.350000 1158.500000 435.650000 ;
      RECT 1116.500000 434.350000 1149.500000 435.650000 ;
      RECT 1107.500000 434.350000 1108.500000 435.650000 ;
      RECT 1066.500000 434.350000 1099.500000 435.650000 ;
      RECT 1057.500000 434.350000 1058.500000 435.650000 ;
      RECT 1016.500000 434.350000 1049.500000 435.650000 ;
      RECT 1007.500000 434.350000 1008.500000 435.650000 ;
      RECT 966.500000 434.350000 999.500000 435.650000 ;
      RECT 957.500000 434.350000 958.500000 435.650000 ;
      RECT 916.500000 434.350000 949.500000 435.650000 ;
      RECT 907.500000 434.350000 908.500000 435.650000 ;
      RECT 866.500000 434.350000 899.500000 435.650000 ;
      RECT 857.500000 434.350000 858.500000 435.650000 ;
      RECT 816.500000 434.350000 849.500000 435.650000 ;
      RECT 807.500000 434.350000 808.500000 435.650000 ;
      RECT 766.500000 434.350000 799.500000 435.650000 ;
      RECT 757.500000 434.350000 758.500000 435.650000 ;
      RECT 722.500000 434.350000 723.500000 435.650000 ;
      RECT 707.500000 434.350000 708.500000 435.650000 ;
      RECT 666.500000 434.350000 699.500000 435.650000 ;
      RECT 657.500000 434.350000 658.500000 435.650000 ;
      RECT 616.500000 434.350000 649.500000 435.650000 ;
      RECT 607.500000 434.350000 608.500000 435.650000 ;
      RECT 566.500000 434.350000 599.500000 435.650000 ;
      RECT 557.500000 434.350000 558.500000 435.650000 ;
      RECT 516.500000 434.350000 549.500000 435.650000 ;
      RECT 507.500000 434.350000 508.500000 435.650000 ;
      RECT 466.500000 434.350000 499.500000 435.650000 ;
      RECT 457.500000 434.350000 458.500000 435.650000 ;
      RECT 416.500000 434.350000 449.500000 435.650000 ;
      RECT 407.500000 434.350000 408.500000 435.650000 ;
      RECT 366.500000 434.350000 399.500000 435.650000 ;
      RECT 357.500000 434.350000 358.500000 435.650000 ;
      RECT 316.500000 434.350000 349.500000 435.650000 ;
      RECT 307.500000 434.350000 308.500000 435.650000 ;
      RECT 216.500000 434.350000 299.500000 435.650000 ;
      RECT 207.500000 434.350000 208.500000 435.650000 ;
      RECT 116.500000 434.350000 199.500000 435.650000 ;
      RECT 107.500000 434.350000 108.500000 435.650000 ;
      RECT 66.500000 434.350000 99.500000 435.650000 ;
      RECT 57.500000 434.350000 58.500000 435.650000 ;
      RECT 29.500000 434.350000 49.500000 435.650000 ;
      RECT 15.500000 434.350000 16.500000 435.650000 ;
      RECT 1157.500000 433.650000 1170.500000 434.350000 ;
      RECT 1107.500000 433.650000 1149.500000 434.350000 ;
      RECT 1057.500000 433.650000 1099.500000 434.350000 ;
      RECT 1007.500000 433.650000 1049.500000 434.350000 ;
      RECT 957.500000 433.650000 999.500000 434.350000 ;
      RECT 907.500000 433.650000 949.500000 434.350000 ;
      RECT 857.500000 433.650000 899.500000 434.350000 ;
      RECT 807.500000 433.650000 849.500000 434.350000 ;
      RECT 757.500000 433.650000 799.500000 434.350000 ;
      RECT 707.500000 433.650000 723.500000 434.350000 ;
      RECT 657.500000 433.650000 699.500000 434.350000 ;
      RECT 607.500000 433.650000 649.500000 434.350000 ;
      RECT 557.500000 433.650000 599.500000 434.350000 ;
      RECT 507.500000 433.650000 549.500000 434.350000 ;
      RECT 457.500000 433.650000 499.500000 434.350000 ;
      RECT 407.500000 433.650000 449.500000 434.350000 ;
      RECT 357.500000 433.650000 399.500000 434.350000 ;
      RECT 307.500000 433.650000 349.500000 434.350000 ;
      RECT 207.500000 433.650000 299.500000 434.350000 ;
      RECT 107.500000 433.650000 199.500000 434.350000 ;
      RECT 57.500000 433.650000 99.500000 434.350000 ;
      RECT 15.500000 433.650000 49.500000 434.350000 ;
      RECT 1183.500000 432.350000 1186.000000 435.650000 ;
      RECT 1166.500000 432.350000 1170.500000 433.650000 ;
      RECT 1157.500000 432.350000 1158.500000 433.650000 ;
      RECT 1116.500000 432.350000 1149.500000 433.650000 ;
      RECT 1107.500000 432.350000 1108.500000 433.650000 ;
      RECT 1066.500000 432.350000 1099.500000 433.650000 ;
      RECT 1057.500000 432.350000 1058.500000 433.650000 ;
      RECT 1016.500000 432.350000 1049.500000 433.650000 ;
      RECT 1007.500000 432.350000 1008.500000 433.650000 ;
      RECT 966.500000 432.350000 999.500000 433.650000 ;
      RECT 957.500000 432.350000 958.500000 433.650000 ;
      RECT 916.500000 432.350000 949.500000 433.650000 ;
      RECT 907.500000 432.350000 908.500000 433.650000 ;
      RECT 866.500000 432.350000 899.500000 433.650000 ;
      RECT 857.500000 432.350000 858.500000 433.650000 ;
      RECT 816.500000 432.350000 849.500000 433.650000 ;
      RECT 807.500000 432.350000 808.500000 433.650000 ;
      RECT 766.500000 432.350000 799.500000 433.650000 ;
      RECT 757.500000 432.350000 758.500000 433.650000 ;
      RECT 736.500000 432.350000 749.500000 435.650000 ;
      RECT 722.500000 432.350000 723.500000 433.650000 ;
      RECT 707.500000 432.350000 708.500000 433.650000 ;
      RECT 666.500000 432.350000 699.500000 433.650000 ;
      RECT 657.500000 432.350000 658.500000 433.650000 ;
      RECT 616.500000 432.350000 649.500000 433.650000 ;
      RECT 607.500000 432.350000 608.500000 433.650000 ;
      RECT 566.500000 432.350000 599.500000 433.650000 ;
      RECT 557.500000 432.350000 558.500000 433.650000 ;
      RECT 516.500000 432.350000 549.500000 433.650000 ;
      RECT 507.500000 432.350000 508.500000 433.650000 ;
      RECT 466.500000 432.350000 499.500000 433.650000 ;
      RECT 457.500000 432.350000 458.500000 433.650000 ;
      RECT 416.500000 432.350000 449.500000 433.650000 ;
      RECT 407.500000 432.350000 408.500000 433.650000 ;
      RECT 366.500000 432.350000 399.500000 433.650000 ;
      RECT 357.500000 432.350000 358.500000 433.650000 ;
      RECT 316.500000 432.350000 349.500000 433.650000 ;
      RECT 307.500000 432.350000 308.500000 433.650000 ;
      RECT 216.500000 432.350000 299.500000 433.650000 ;
      RECT 207.500000 432.350000 208.500000 433.650000 ;
      RECT 116.500000 432.350000 199.500000 433.650000 ;
      RECT 107.500000 432.350000 108.500000 433.650000 ;
      RECT 66.500000 432.350000 99.500000 433.650000 ;
      RECT 57.500000 432.350000 58.500000 433.650000 ;
      RECT 29.500000 432.350000 49.500000 433.650000 ;
      RECT 15.500000 432.350000 16.500000 433.650000 ;
      RECT 0.000000 432.350000 2.500000 435.650000 ;
      RECT 1166.500000 431.650000 1186.000000 432.350000 ;
      RECT 1116.500000 431.650000 1158.500000 432.350000 ;
      RECT 1066.500000 431.650000 1108.500000 432.350000 ;
      RECT 1016.500000 431.650000 1058.500000 432.350000 ;
      RECT 966.500000 431.650000 1008.500000 432.350000 ;
      RECT 916.500000 431.650000 958.500000 432.350000 ;
      RECT 866.500000 431.650000 908.500000 432.350000 ;
      RECT 816.500000 431.650000 858.500000 432.350000 ;
      RECT 766.500000 431.650000 808.500000 432.350000 ;
      RECT 722.500000 431.650000 758.500000 432.350000 ;
      RECT 666.500000 431.650000 708.500000 432.350000 ;
      RECT 616.500000 431.650000 658.500000 432.350000 ;
      RECT 566.500000 431.650000 608.500000 432.350000 ;
      RECT 516.500000 431.650000 558.500000 432.350000 ;
      RECT 466.500000 431.650000 508.500000 432.350000 ;
      RECT 416.500000 431.650000 458.500000 432.350000 ;
      RECT 366.500000 431.650000 408.500000 432.350000 ;
      RECT 316.500000 431.650000 358.500000 432.350000 ;
      RECT 216.500000 431.650000 308.500000 432.350000 ;
      RECT 116.500000 431.650000 208.500000 432.350000 ;
      RECT 66.500000 431.650000 108.500000 432.350000 ;
      RECT 29.500000 431.650000 58.500000 432.350000 ;
      RECT 0.000000 431.650000 16.500000 432.350000 ;
      RECT 1166.500000 430.350000 1170.500000 431.650000 ;
      RECT 1157.500000 430.350000 1158.500000 431.650000 ;
      RECT 1116.500000 430.350000 1149.500000 431.650000 ;
      RECT 1107.500000 430.350000 1108.500000 431.650000 ;
      RECT 1066.500000 430.350000 1099.500000 431.650000 ;
      RECT 1057.500000 430.350000 1058.500000 431.650000 ;
      RECT 1016.500000 430.350000 1049.500000 431.650000 ;
      RECT 1007.500000 430.350000 1008.500000 431.650000 ;
      RECT 966.500000 430.350000 999.500000 431.650000 ;
      RECT 957.500000 430.350000 958.500000 431.650000 ;
      RECT 916.500000 430.350000 949.500000 431.650000 ;
      RECT 907.500000 430.350000 908.500000 431.650000 ;
      RECT 866.500000 430.350000 899.500000 431.650000 ;
      RECT 857.500000 430.350000 858.500000 431.650000 ;
      RECT 816.500000 430.350000 849.500000 431.650000 ;
      RECT 807.500000 430.350000 808.500000 431.650000 ;
      RECT 766.500000 430.350000 799.500000 431.650000 ;
      RECT 757.500000 430.350000 758.500000 431.650000 ;
      RECT 722.500000 430.350000 749.500000 431.650000 ;
      RECT 707.500000 430.350000 708.500000 431.650000 ;
      RECT 666.500000 430.350000 699.500000 431.650000 ;
      RECT 657.500000 430.350000 658.500000 431.650000 ;
      RECT 616.500000 430.350000 649.500000 431.650000 ;
      RECT 607.500000 430.350000 608.500000 431.650000 ;
      RECT 566.500000 430.350000 599.500000 431.650000 ;
      RECT 557.500000 430.350000 558.500000 431.650000 ;
      RECT 516.500000 430.350000 549.500000 431.650000 ;
      RECT 507.500000 430.350000 508.500000 431.650000 ;
      RECT 466.500000 430.350000 499.500000 431.650000 ;
      RECT 457.500000 430.350000 458.500000 431.650000 ;
      RECT 416.500000 430.350000 449.500000 431.650000 ;
      RECT 407.500000 430.350000 408.500000 431.650000 ;
      RECT 366.500000 430.350000 399.500000 431.650000 ;
      RECT 357.500000 430.350000 358.500000 431.650000 ;
      RECT 316.500000 430.350000 349.500000 431.650000 ;
      RECT 307.500000 430.350000 308.500000 431.650000 ;
      RECT 216.500000 430.350000 299.500000 431.650000 ;
      RECT 207.500000 430.350000 208.500000 431.650000 ;
      RECT 116.500000 430.350000 199.500000 431.650000 ;
      RECT 107.500000 430.350000 108.500000 431.650000 ;
      RECT 66.500000 430.350000 99.500000 431.650000 ;
      RECT 57.500000 430.350000 58.500000 431.650000 ;
      RECT 29.500000 430.350000 49.500000 431.650000 ;
      RECT 15.500000 430.350000 16.500000 431.650000 ;
      RECT 1157.500000 429.650000 1170.500000 430.350000 ;
      RECT 1107.500000 429.650000 1149.500000 430.350000 ;
      RECT 1057.500000 429.650000 1099.500000 430.350000 ;
      RECT 1007.500000 429.650000 1049.500000 430.350000 ;
      RECT 957.500000 429.650000 999.500000 430.350000 ;
      RECT 907.500000 429.650000 949.500000 430.350000 ;
      RECT 857.500000 429.650000 899.500000 430.350000 ;
      RECT 807.500000 429.650000 849.500000 430.350000 ;
      RECT 757.500000 429.650000 799.500000 430.350000 ;
      RECT 707.500000 429.650000 749.500000 430.350000 ;
      RECT 657.500000 429.650000 699.500000 430.350000 ;
      RECT 607.500000 429.650000 649.500000 430.350000 ;
      RECT 557.500000 429.650000 599.500000 430.350000 ;
      RECT 507.500000 429.650000 549.500000 430.350000 ;
      RECT 457.500000 429.650000 499.500000 430.350000 ;
      RECT 407.500000 429.650000 449.500000 430.350000 ;
      RECT 357.500000 429.650000 399.500000 430.350000 ;
      RECT 307.500000 429.650000 349.500000 430.350000 ;
      RECT 207.500000 429.650000 299.500000 430.350000 ;
      RECT 107.500000 429.650000 199.500000 430.350000 ;
      RECT 57.500000 429.650000 99.500000 430.350000 ;
      RECT 15.500000 429.650000 49.500000 430.350000 ;
      RECT 1183.500000 428.350000 1186.000000 431.650000 ;
      RECT 1169.500000 428.350000 1170.500000 429.650000 ;
      RECT 1116.500000 428.350000 1149.500000 429.650000 ;
      RECT 1107.500000 428.350000 1108.500000 429.650000 ;
      RECT 1066.500000 428.350000 1099.500000 429.650000 ;
      RECT 1057.500000 428.350000 1058.500000 429.650000 ;
      RECT 1016.500000 428.350000 1049.500000 429.650000 ;
      RECT 1007.500000 428.350000 1008.500000 429.650000 ;
      RECT 966.500000 428.350000 999.500000 429.650000 ;
      RECT 957.500000 428.350000 958.500000 429.650000 ;
      RECT 916.500000 428.350000 949.500000 429.650000 ;
      RECT 907.500000 428.350000 908.500000 429.650000 ;
      RECT 866.500000 428.350000 899.500000 429.650000 ;
      RECT 857.500000 428.350000 858.500000 429.650000 ;
      RECT 816.500000 428.350000 849.500000 429.650000 ;
      RECT 807.500000 428.350000 808.500000 429.650000 ;
      RECT 766.500000 428.350000 799.500000 429.650000 ;
      RECT 757.500000 428.350000 758.500000 429.650000 ;
      RECT 722.500000 428.350000 749.500000 429.650000 ;
      RECT 707.500000 428.350000 709.500000 429.650000 ;
      RECT 666.500000 428.350000 699.500000 429.650000 ;
      RECT 657.500000 428.350000 658.500000 429.650000 ;
      RECT 616.500000 428.350000 649.500000 429.650000 ;
      RECT 607.500000 428.350000 608.500000 429.650000 ;
      RECT 566.500000 428.350000 599.500000 429.650000 ;
      RECT 557.500000 428.350000 558.500000 429.650000 ;
      RECT 516.500000 428.350000 549.500000 429.650000 ;
      RECT 507.500000 428.350000 508.500000 429.650000 ;
      RECT 466.500000 428.350000 499.500000 429.650000 ;
      RECT 457.500000 428.350000 458.500000 429.650000 ;
      RECT 416.500000 428.350000 449.500000 429.650000 ;
      RECT 407.500000 428.350000 408.500000 429.650000 ;
      RECT 366.500000 428.350000 399.500000 429.650000 ;
      RECT 357.500000 428.350000 358.500000 429.650000 ;
      RECT 316.500000 428.350000 349.500000 429.650000 ;
      RECT 307.500000 428.350000 308.500000 429.650000 ;
      RECT 216.500000 428.350000 299.500000 429.650000 ;
      RECT 207.500000 428.350000 208.500000 429.650000 ;
      RECT 116.500000 428.350000 199.500000 429.650000 ;
      RECT 107.500000 428.350000 108.500000 429.650000 ;
      RECT 66.500000 428.350000 99.500000 429.650000 ;
      RECT 57.500000 428.350000 58.500000 429.650000 ;
      RECT 29.500000 428.350000 49.500000 429.650000 ;
      RECT 15.500000 428.350000 16.500000 429.650000 ;
      RECT 0.000000 428.350000 2.500000 431.650000 ;
      RECT 1169.500000 427.650000 1186.000000 428.350000 ;
      RECT 1116.500000 427.650000 1156.500000 428.350000 ;
      RECT 1066.500000 427.650000 1108.500000 428.350000 ;
      RECT 1016.500000 427.650000 1058.500000 428.350000 ;
      RECT 966.500000 427.650000 1008.500000 428.350000 ;
      RECT 916.500000 427.650000 958.500000 428.350000 ;
      RECT 866.500000 427.650000 908.500000 428.350000 ;
      RECT 816.500000 427.650000 858.500000 428.350000 ;
      RECT 766.500000 427.650000 808.500000 428.350000 ;
      RECT 722.500000 427.650000 758.500000 428.350000 ;
      RECT 666.500000 427.650000 709.500000 428.350000 ;
      RECT 616.500000 427.650000 658.500000 428.350000 ;
      RECT 566.500000 427.650000 608.500000 428.350000 ;
      RECT 516.500000 427.650000 558.500000 428.350000 ;
      RECT 466.500000 427.650000 508.500000 428.350000 ;
      RECT 416.500000 427.650000 458.500000 428.350000 ;
      RECT 366.500000 427.650000 408.500000 428.350000 ;
      RECT 316.500000 427.650000 358.500000 428.350000 ;
      RECT 216.500000 427.650000 308.500000 428.350000 ;
      RECT 116.500000 427.650000 208.500000 428.350000 ;
      RECT 66.500000 427.650000 108.500000 428.350000 ;
      RECT 29.500000 427.650000 58.500000 428.350000 ;
      RECT 0.000000 427.650000 16.500000 428.350000 ;
      RECT 1169.500000 426.350000 1170.500000 427.650000 ;
      RECT 1116.500000 426.350000 1149.500000 427.650000 ;
      RECT 1107.500000 426.350000 1108.500000 427.650000 ;
      RECT 1066.500000 426.350000 1099.500000 427.650000 ;
      RECT 1057.500000 426.350000 1058.500000 427.650000 ;
      RECT 1016.500000 426.350000 1049.500000 427.650000 ;
      RECT 1007.500000 426.350000 1008.500000 427.650000 ;
      RECT 966.500000 426.350000 999.500000 427.650000 ;
      RECT 957.500000 426.350000 958.500000 427.650000 ;
      RECT 916.500000 426.350000 949.500000 427.650000 ;
      RECT 907.500000 426.350000 908.500000 427.650000 ;
      RECT 866.500000 426.350000 899.500000 427.650000 ;
      RECT 857.500000 426.350000 858.500000 427.650000 ;
      RECT 816.500000 426.350000 849.500000 427.650000 ;
      RECT 807.500000 426.350000 808.500000 427.650000 ;
      RECT 766.500000 426.350000 799.500000 427.650000 ;
      RECT 757.500000 426.350000 758.500000 427.650000 ;
      RECT 722.500000 426.350000 749.500000 427.650000 ;
      RECT 707.500000 426.350000 709.500000 427.650000 ;
      RECT 666.500000 426.350000 699.500000 427.650000 ;
      RECT 657.500000 426.350000 658.500000 427.650000 ;
      RECT 616.500000 426.350000 649.500000 427.650000 ;
      RECT 607.500000 426.350000 608.500000 427.650000 ;
      RECT 566.500000 426.350000 599.500000 427.650000 ;
      RECT 557.500000 426.350000 558.500000 427.650000 ;
      RECT 516.500000 426.350000 549.500000 427.650000 ;
      RECT 507.500000 426.350000 508.500000 427.650000 ;
      RECT 466.500000 426.350000 499.500000 427.650000 ;
      RECT 457.500000 426.350000 458.500000 427.650000 ;
      RECT 416.500000 426.350000 449.500000 427.650000 ;
      RECT 407.500000 426.350000 408.500000 427.650000 ;
      RECT 366.500000 426.350000 399.500000 427.650000 ;
      RECT 357.500000 426.350000 358.500000 427.650000 ;
      RECT 316.500000 426.350000 349.500000 427.650000 ;
      RECT 307.500000 426.350000 308.500000 427.650000 ;
      RECT 216.500000 426.350000 299.500000 427.650000 ;
      RECT 207.500000 426.350000 208.500000 427.650000 ;
      RECT 116.500000 426.350000 199.500000 427.650000 ;
      RECT 107.500000 426.350000 108.500000 427.650000 ;
      RECT 66.500000 426.350000 99.500000 427.650000 ;
      RECT 57.500000 426.350000 58.500000 427.650000 ;
      RECT 29.500000 426.350000 49.500000 427.650000 ;
      RECT 15.500000 426.350000 16.500000 427.650000 ;
      RECT 1157.500000 425.650000 1170.500000 426.350000 ;
      RECT 1107.500000 425.650000 1149.500000 426.350000 ;
      RECT 1057.500000 425.650000 1099.500000 426.350000 ;
      RECT 1007.500000 425.650000 1049.500000 426.350000 ;
      RECT 957.500000 425.650000 999.500000 426.350000 ;
      RECT 907.500000 425.650000 949.500000 426.350000 ;
      RECT 857.500000 425.650000 899.500000 426.350000 ;
      RECT 807.500000 425.650000 849.500000 426.350000 ;
      RECT 757.500000 425.650000 799.500000 426.350000 ;
      RECT 707.500000 425.650000 749.500000 426.350000 ;
      RECT 657.500000 425.650000 699.500000 426.350000 ;
      RECT 607.500000 425.650000 649.500000 426.350000 ;
      RECT 557.500000 425.650000 599.500000 426.350000 ;
      RECT 507.500000 425.650000 549.500000 426.350000 ;
      RECT 457.500000 425.650000 499.500000 426.350000 ;
      RECT 407.500000 425.650000 449.500000 426.350000 ;
      RECT 357.500000 425.650000 399.500000 426.350000 ;
      RECT 307.500000 425.650000 349.500000 426.350000 ;
      RECT 207.500000 425.650000 299.500000 426.350000 ;
      RECT 107.500000 425.650000 199.500000 426.350000 ;
      RECT 57.500000 425.650000 99.500000 426.350000 ;
      RECT 15.500000 425.650000 49.500000 426.350000 ;
      RECT 1183.500000 424.350000 1186.000000 427.650000 ;
      RECT 1169.500000 424.350000 1170.500000 425.650000 ;
      RECT 1116.500000 424.350000 1149.500000 425.650000 ;
      RECT 1107.500000 424.350000 1108.500000 425.650000 ;
      RECT 1066.500000 424.350000 1099.500000 425.650000 ;
      RECT 1057.500000 424.350000 1058.500000 425.650000 ;
      RECT 1016.500000 424.350000 1049.500000 425.650000 ;
      RECT 1007.500000 424.350000 1008.500000 425.650000 ;
      RECT 966.500000 424.350000 999.500000 425.650000 ;
      RECT 957.500000 424.350000 958.500000 425.650000 ;
      RECT 916.500000 424.350000 949.500000 425.650000 ;
      RECT 907.500000 424.350000 908.500000 425.650000 ;
      RECT 866.500000 424.350000 899.500000 425.650000 ;
      RECT 857.500000 424.350000 858.500000 425.650000 ;
      RECT 816.500000 424.350000 849.500000 425.650000 ;
      RECT 807.500000 424.350000 808.500000 425.650000 ;
      RECT 766.500000 424.350000 799.500000 425.650000 ;
      RECT 757.500000 424.350000 758.500000 425.650000 ;
      RECT 722.500000 424.350000 749.500000 425.650000 ;
      RECT 707.500000 424.350000 709.500000 425.650000 ;
      RECT 666.500000 424.350000 699.500000 425.650000 ;
      RECT 657.500000 424.350000 658.500000 425.650000 ;
      RECT 616.500000 424.350000 649.500000 425.650000 ;
      RECT 607.500000 424.350000 608.500000 425.650000 ;
      RECT 566.500000 424.350000 599.500000 425.650000 ;
      RECT 557.500000 424.350000 558.500000 425.650000 ;
      RECT 516.500000 424.350000 549.500000 425.650000 ;
      RECT 507.500000 424.350000 508.500000 425.650000 ;
      RECT 466.500000 424.350000 499.500000 425.650000 ;
      RECT 457.500000 424.350000 458.500000 425.650000 ;
      RECT 416.500000 424.350000 449.500000 425.650000 ;
      RECT 407.500000 424.350000 408.500000 425.650000 ;
      RECT 366.500000 424.350000 399.500000 425.650000 ;
      RECT 357.500000 424.350000 358.500000 425.650000 ;
      RECT 316.500000 424.350000 349.500000 425.650000 ;
      RECT 307.500000 424.350000 308.500000 425.650000 ;
      RECT 216.500000 424.350000 299.500000 425.650000 ;
      RECT 207.500000 424.350000 208.500000 425.650000 ;
      RECT 116.500000 424.350000 199.500000 425.650000 ;
      RECT 107.500000 424.350000 108.500000 425.650000 ;
      RECT 66.500000 424.350000 99.500000 425.650000 ;
      RECT 57.500000 424.350000 58.500000 425.650000 ;
      RECT 29.500000 424.350000 49.500000 425.650000 ;
      RECT 15.500000 424.350000 16.500000 425.650000 ;
      RECT 0.000000 424.350000 2.500000 427.650000 ;
      RECT 1169.500000 423.650000 1186.000000 424.350000 ;
      RECT 1116.500000 423.650000 1156.500000 424.350000 ;
      RECT 1066.500000 423.650000 1108.500000 424.350000 ;
      RECT 1016.500000 423.650000 1058.500000 424.350000 ;
      RECT 966.500000 423.650000 1008.500000 424.350000 ;
      RECT 916.500000 423.650000 958.500000 424.350000 ;
      RECT 866.500000 423.650000 908.500000 424.350000 ;
      RECT 816.500000 423.650000 858.500000 424.350000 ;
      RECT 766.500000 423.650000 808.500000 424.350000 ;
      RECT 722.500000 423.650000 758.500000 424.350000 ;
      RECT 666.500000 423.650000 709.500000 424.350000 ;
      RECT 616.500000 423.650000 658.500000 424.350000 ;
      RECT 566.500000 423.650000 608.500000 424.350000 ;
      RECT 516.500000 423.650000 558.500000 424.350000 ;
      RECT 466.500000 423.650000 508.500000 424.350000 ;
      RECT 416.500000 423.650000 458.500000 424.350000 ;
      RECT 366.500000 423.650000 408.500000 424.350000 ;
      RECT 316.500000 423.650000 358.500000 424.350000 ;
      RECT 216.500000 423.650000 308.500000 424.350000 ;
      RECT 116.500000 423.650000 208.500000 424.350000 ;
      RECT 66.500000 423.650000 108.500000 424.350000 ;
      RECT 29.500000 423.650000 58.500000 424.350000 ;
      RECT 0.000000 423.650000 16.500000 424.350000 ;
      RECT 1169.500000 422.350000 1170.500000 423.650000 ;
      RECT 1116.500000 422.350000 1149.500000 423.650000 ;
      RECT 1107.500000 422.350000 1108.500000 423.650000 ;
      RECT 1066.500000 422.350000 1099.500000 423.650000 ;
      RECT 1057.500000 422.350000 1058.500000 423.650000 ;
      RECT 1016.500000 422.350000 1049.500000 423.650000 ;
      RECT 1007.500000 422.350000 1008.500000 423.650000 ;
      RECT 966.500000 422.350000 999.500000 423.650000 ;
      RECT 957.500000 422.350000 958.500000 423.650000 ;
      RECT 916.500000 422.350000 949.500000 423.650000 ;
      RECT 907.500000 422.350000 908.500000 423.650000 ;
      RECT 866.500000 422.350000 899.500000 423.650000 ;
      RECT 857.500000 422.350000 858.500000 423.650000 ;
      RECT 816.500000 422.350000 849.500000 423.650000 ;
      RECT 807.500000 422.350000 808.500000 423.650000 ;
      RECT 766.500000 422.350000 799.500000 423.650000 ;
      RECT 757.500000 422.350000 758.500000 423.650000 ;
      RECT 722.500000 422.350000 749.500000 423.650000 ;
      RECT 707.500000 422.350000 709.500000 423.650000 ;
      RECT 666.500000 422.350000 699.500000 423.650000 ;
      RECT 657.500000 422.350000 658.500000 423.650000 ;
      RECT 616.500000 422.350000 649.500000 423.650000 ;
      RECT 607.500000 422.350000 608.500000 423.650000 ;
      RECT 566.500000 422.350000 599.500000 423.650000 ;
      RECT 557.500000 422.350000 558.500000 423.650000 ;
      RECT 516.500000 422.350000 549.500000 423.650000 ;
      RECT 507.500000 422.350000 508.500000 423.650000 ;
      RECT 466.500000 422.350000 499.500000 423.650000 ;
      RECT 457.500000 422.350000 458.500000 423.650000 ;
      RECT 416.500000 422.350000 449.500000 423.650000 ;
      RECT 407.500000 422.350000 408.500000 423.650000 ;
      RECT 366.500000 422.350000 399.500000 423.650000 ;
      RECT 357.500000 422.350000 358.500000 423.650000 ;
      RECT 316.500000 422.350000 349.500000 423.650000 ;
      RECT 307.500000 422.350000 308.500000 423.650000 ;
      RECT 216.500000 422.350000 299.500000 423.650000 ;
      RECT 207.500000 422.350000 208.500000 423.650000 ;
      RECT 116.500000 422.350000 199.500000 423.650000 ;
      RECT 107.500000 422.350000 108.500000 423.650000 ;
      RECT 66.500000 422.350000 99.500000 423.650000 ;
      RECT 57.500000 422.350000 58.500000 423.650000 ;
      RECT 29.500000 422.350000 49.500000 423.650000 ;
      RECT 15.500000 422.350000 16.500000 423.650000 ;
      RECT 1157.500000 421.650000 1170.500000 422.350000 ;
      RECT 1107.500000 421.650000 1149.500000 422.350000 ;
      RECT 1057.500000 421.650000 1099.500000 422.350000 ;
      RECT 1007.500000 421.650000 1049.500000 422.350000 ;
      RECT 957.500000 421.650000 999.500000 422.350000 ;
      RECT 907.500000 421.650000 949.500000 422.350000 ;
      RECT 857.500000 421.650000 899.500000 422.350000 ;
      RECT 807.500000 421.650000 849.500000 422.350000 ;
      RECT 757.500000 421.650000 799.500000 422.350000 ;
      RECT 707.500000 421.650000 749.500000 422.350000 ;
      RECT 657.500000 421.650000 699.500000 422.350000 ;
      RECT 607.500000 421.650000 649.500000 422.350000 ;
      RECT 557.500000 421.650000 599.500000 422.350000 ;
      RECT 507.500000 421.650000 549.500000 422.350000 ;
      RECT 457.500000 421.650000 499.500000 422.350000 ;
      RECT 407.500000 421.650000 449.500000 422.350000 ;
      RECT 357.500000 421.650000 399.500000 422.350000 ;
      RECT 307.500000 421.650000 349.500000 422.350000 ;
      RECT 207.500000 421.650000 299.500000 422.350000 ;
      RECT 107.500000 421.650000 199.500000 422.350000 ;
      RECT 57.500000 421.650000 99.500000 422.350000 ;
      RECT 15.500000 421.650000 49.500000 422.350000 ;
      RECT 1183.500000 420.350000 1186.000000 423.650000 ;
      RECT 1169.500000 420.350000 1170.500000 421.650000 ;
      RECT 1116.500000 420.350000 1149.500000 421.650000 ;
      RECT 1107.500000 420.350000 1108.500000 421.650000 ;
      RECT 1066.500000 420.350000 1099.500000 421.650000 ;
      RECT 1057.500000 420.350000 1058.500000 421.650000 ;
      RECT 1016.500000 420.350000 1049.500000 421.650000 ;
      RECT 1007.500000 420.350000 1008.500000 421.650000 ;
      RECT 966.500000 420.350000 999.500000 421.650000 ;
      RECT 957.500000 420.350000 958.500000 421.650000 ;
      RECT 916.500000 420.350000 949.500000 421.650000 ;
      RECT 907.500000 420.350000 908.500000 421.650000 ;
      RECT 866.500000 420.350000 899.500000 421.650000 ;
      RECT 857.500000 420.350000 858.500000 421.650000 ;
      RECT 816.500000 420.350000 849.500000 421.650000 ;
      RECT 807.500000 420.350000 808.500000 421.650000 ;
      RECT 766.500000 420.350000 799.500000 421.650000 ;
      RECT 757.500000 420.350000 758.500000 421.650000 ;
      RECT 722.500000 420.350000 749.500000 421.650000 ;
      RECT 707.500000 420.350000 709.500000 421.650000 ;
      RECT 666.500000 420.350000 699.500000 421.650000 ;
      RECT 657.500000 420.350000 658.500000 421.650000 ;
      RECT 616.500000 420.350000 649.500000 421.650000 ;
      RECT 607.500000 420.350000 608.500000 421.650000 ;
      RECT 566.500000 420.350000 599.500000 421.650000 ;
      RECT 557.500000 420.350000 558.500000 421.650000 ;
      RECT 516.500000 420.350000 549.500000 421.650000 ;
      RECT 507.500000 420.350000 508.500000 421.650000 ;
      RECT 466.500000 420.350000 499.500000 421.650000 ;
      RECT 457.500000 420.350000 458.500000 421.650000 ;
      RECT 416.500000 420.350000 449.500000 421.650000 ;
      RECT 407.500000 420.350000 408.500000 421.650000 ;
      RECT 366.500000 420.350000 399.500000 421.650000 ;
      RECT 357.500000 420.350000 358.500000 421.650000 ;
      RECT 316.500000 420.350000 349.500000 421.650000 ;
      RECT 307.500000 420.350000 308.500000 421.650000 ;
      RECT 216.500000 420.350000 299.500000 421.650000 ;
      RECT 207.500000 420.350000 208.500000 421.650000 ;
      RECT 116.500000 420.350000 199.500000 421.650000 ;
      RECT 107.500000 420.350000 108.500000 421.650000 ;
      RECT 66.500000 420.350000 99.500000 421.650000 ;
      RECT 57.500000 420.350000 58.500000 421.650000 ;
      RECT 29.500000 420.350000 49.500000 421.650000 ;
      RECT 15.500000 420.350000 16.500000 421.650000 ;
      RECT 0.000000 420.350000 2.500000 423.650000 ;
      RECT 1169.500000 419.650000 1186.000000 420.350000 ;
      RECT 1116.500000 419.650000 1156.500000 420.350000 ;
      RECT 1066.500000 419.650000 1108.500000 420.350000 ;
      RECT 1016.500000 419.650000 1058.500000 420.350000 ;
      RECT 966.500000 419.650000 1008.500000 420.350000 ;
      RECT 916.500000 419.650000 958.500000 420.350000 ;
      RECT 866.500000 419.650000 908.500000 420.350000 ;
      RECT 816.500000 419.650000 858.500000 420.350000 ;
      RECT 766.500000 419.650000 808.500000 420.350000 ;
      RECT 722.500000 419.650000 758.500000 420.350000 ;
      RECT 666.500000 419.650000 709.500000 420.350000 ;
      RECT 616.500000 419.650000 658.500000 420.350000 ;
      RECT 566.500000 419.650000 608.500000 420.350000 ;
      RECT 516.500000 419.650000 558.500000 420.350000 ;
      RECT 466.500000 419.650000 508.500000 420.350000 ;
      RECT 366.500000 419.650000 408.500000 420.350000 ;
      RECT 316.500000 419.650000 358.500000 420.350000 ;
      RECT 216.500000 419.650000 308.500000 420.350000 ;
      RECT 116.500000 419.650000 208.500000 420.350000 ;
      RECT 66.500000 419.650000 108.500000 420.350000 ;
      RECT 29.500000 419.650000 58.500000 420.350000 ;
      RECT 0.000000 419.650000 16.500000 420.350000 ;
      RECT 1169.500000 418.350000 1170.500000 419.650000 ;
      RECT 1116.500000 418.350000 1149.500000 419.650000 ;
      RECT 1107.500000 418.350000 1108.500000 419.650000 ;
      RECT 1066.500000 418.350000 1099.500000 419.650000 ;
      RECT 1057.500000 418.350000 1058.500000 419.650000 ;
      RECT 1016.500000 418.350000 1049.500000 419.650000 ;
      RECT 1007.500000 418.350000 1008.500000 419.650000 ;
      RECT 966.500000 418.350000 999.500000 419.650000 ;
      RECT 957.500000 418.350000 958.500000 419.650000 ;
      RECT 916.500000 418.350000 949.500000 419.650000 ;
      RECT 907.500000 418.350000 908.500000 419.650000 ;
      RECT 866.500000 418.350000 899.500000 419.650000 ;
      RECT 857.500000 418.350000 858.500000 419.650000 ;
      RECT 816.500000 418.350000 849.500000 419.650000 ;
      RECT 807.500000 418.350000 808.500000 419.650000 ;
      RECT 766.500000 418.350000 799.500000 419.650000 ;
      RECT 757.500000 418.350000 758.500000 419.650000 ;
      RECT 722.500000 418.350000 749.500000 419.650000 ;
      RECT 707.500000 418.350000 709.500000 419.650000 ;
      RECT 666.500000 418.350000 699.500000 419.650000 ;
      RECT 657.500000 418.350000 658.500000 419.650000 ;
      RECT 616.500000 418.350000 649.500000 419.650000 ;
      RECT 607.500000 418.350000 608.500000 419.650000 ;
      RECT 566.500000 418.350000 599.500000 419.650000 ;
      RECT 557.500000 418.350000 558.500000 419.650000 ;
      RECT 516.500000 418.350000 549.500000 419.650000 ;
      RECT 507.500000 418.350000 508.500000 419.650000 ;
      RECT 466.500000 418.350000 499.500000 419.650000 ;
      RECT 416.500000 418.350000 458.500000 420.350000 ;
      RECT 407.500000 418.350000 408.500000 419.650000 ;
      RECT 366.500000 418.350000 399.500000 419.650000 ;
      RECT 357.500000 418.350000 358.500000 419.650000 ;
      RECT 316.500000 418.350000 349.500000 419.650000 ;
      RECT 307.500000 418.350000 308.500000 419.650000 ;
      RECT 216.500000 418.350000 299.500000 419.650000 ;
      RECT 207.500000 418.350000 208.500000 419.650000 ;
      RECT 116.500000 418.350000 199.500000 419.650000 ;
      RECT 107.500000 418.350000 108.500000 419.650000 ;
      RECT 66.500000 418.350000 99.500000 419.650000 ;
      RECT 57.500000 418.350000 58.500000 419.650000 ;
      RECT 29.500000 418.350000 49.500000 419.650000 ;
      RECT 15.500000 418.350000 16.500000 419.650000 ;
      RECT 1157.500000 417.650000 1170.500000 418.350000 ;
      RECT 1107.500000 417.650000 1149.500000 418.350000 ;
      RECT 1057.500000 417.650000 1099.500000 418.350000 ;
      RECT 1007.500000 417.650000 1049.500000 418.350000 ;
      RECT 957.500000 417.650000 999.500000 418.350000 ;
      RECT 907.500000 417.650000 949.500000 418.350000 ;
      RECT 857.500000 417.650000 899.500000 418.350000 ;
      RECT 807.500000 417.650000 849.500000 418.350000 ;
      RECT 757.500000 417.650000 799.500000 418.350000 ;
      RECT 707.500000 417.650000 749.500000 418.350000 ;
      RECT 657.500000 417.650000 699.500000 418.350000 ;
      RECT 607.500000 417.650000 649.500000 418.350000 ;
      RECT 557.500000 417.650000 599.500000 418.350000 ;
      RECT 507.500000 417.650000 549.500000 418.350000 ;
      RECT 407.500000 417.650000 499.500000 418.350000 ;
      RECT 357.500000 417.650000 399.500000 418.350000 ;
      RECT 307.500000 417.650000 349.500000 418.350000 ;
      RECT 207.500000 417.650000 299.500000 418.350000 ;
      RECT 107.500000 417.650000 199.500000 418.350000 ;
      RECT 57.500000 417.650000 99.500000 418.350000 ;
      RECT 15.500000 417.650000 49.500000 418.350000 ;
      RECT 1183.500000 416.350000 1186.000000 419.650000 ;
      RECT 1169.500000 416.350000 1170.500000 417.650000 ;
      RECT 1116.500000 416.350000 1149.500000 417.650000 ;
      RECT 1107.500000 416.350000 1108.500000 417.650000 ;
      RECT 1066.500000 416.350000 1099.500000 417.650000 ;
      RECT 1057.500000 416.350000 1058.500000 417.650000 ;
      RECT 1016.500000 416.350000 1049.500000 417.650000 ;
      RECT 1007.500000 416.350000 1008.500000 417.650000 ;
      RECT 966.500000 416.350000 999.500000 417.650000 ;
      RECT 957.500000 416.350000 958.500000 417.650000 ;
      RECT 916.500000 416.350000 949.500000 417.650000 ;
      RECT 907.500000 416.350000 908.500000 417.650000 ;
      RECT 866.500000 416.350000 899.500000 417.650000 ;
      RECT 857.500000 416.350000 858.500000 417.650000 ;
      RECT 816.500000 416.350000 849.500000 417.650000 ;
      RECT 807.500000 416.350000 808.500000 417.650000 ;
      RECT 766.500000 416.350000 799.500000 417.650000 ;
      RECT 757.500000 416.350000 758.500000 417.650000 ;
      RECT 720.000000 416.350000 749.500000 417.650000 ;
      RECT 707.500000 416.350000 712.000000 417.650000 ;
      RECT 666.500000 416.350000 699.500000 417.650000 ;
      RECT 657.500000 416.350000 658.500000 417.650000 ;
      RECT 616.500000 416.350000 649.500000 417.650000 ;
      RECT 607.500000 416.350000 608.500000 417.650000 ;
      RECT 566.500000 416.350000 599.500000 417.650000 ;
      RECT 557.500000 416.350000 558.500000 417.650000 ;
      RECT 516.500000 416.350000 549.500000 417.650000 ;
      RECT 507.500000 416.350000 508.500000 417.650000 ;
      RECT 416.500000 416.350000 499.500000 417.650000 ;
      RECT 407.500000 416.350000 408.500000 417.650000 ;
      RECT 366.500000 416.350000 399.500000 417.650000 ;
      RECT 357.500000 416.350000 358.500000 417.650000 ;
      RECT 316.500000 416.350000 349.500000 417.650000 ;
      RECT 307.500000 416.350000 308.500000 417.650000 ;
      RECT 216.500000 416.350000 299.500000 417.650000 ;
      RECT 207.500000 416.350000 208.500000 417.650000 ;
      RECT 116.500000 416.350000 199.500000 417.650000 ;
      RECT 107.500000 416.350000 108.500000 417.650000 ;
      RECT 66.500000 416.350000 99.500000 417.650000 ;
      RECT 57.500000 416.350000 58.500000 417.650000 ;
      RECT 29.500000 416.350000 49.500000 417.650000 ;
      RECT 15.500000 416.350000 16.500000 417.650000 ;
      RECT 0.000000 416.350000 2.500000 419.650000 ;
      RECT 1169.500000 415.650000 1186.000000 416.350000 ;
      RECT 1116.500000 415.650000 1156.500000 416.350000 ;
      RECT 1066.500000 415.650000 1108.500000 416.350000 ;
      RECT 1016.500000 415.650000 1058.500000 416.350000 ;
      RECT 966.500000 415.650000 1008.500000 416.350000 ;
      RECT 916.500000 415.650000 958.500000 416.350000 ;
      RECT 866.500000 415.650000 908.500000 416.350000 ;
      RECT 816.500000 415.650000 858.500000 416.350000 ;
      RECT 766.500000 415.650000 808.500000 416.350000 ;
      RECT 720.000000 415.650000 758.500000 416.350000 ;
      RECT 666.500000 415.650000 712.000000 416.350000 ;
      RECT 616.500000 415.650000 658.500000 416.350000 ;
      RECT 566.500000 415.650000 608.500000 416.350000 ;
      RECT 516.500000 415.650000 558.500000 416.350000 ;
      RECT 416.500000 415.650000 508.500000 416.350000 ;
      RECT 366.500000 415.650000 408.500000 416.350000 ;
      RECT 316.500000 415.650000 358.500000 416.350000 ;
      RECT 216.500000 415.650000 308.500000 416.350000 ;
      RECT 116.500000 415.650000 208.500000 416.350000 ;
      RECT 66.500000 415.650000 108.500000 416.350000 ;
      RECT 29.500000 415.650000 58.500000 416.350000 ;
      RECT 0.000000 415.650000 16.500000 416.350000 ;
      RECT 1169.500000 414.350000 1170.500000 415.650000 ;
      RECT 1116.500000 414.350000 1149.500000 415.650000 ;
      RECT 1107.500000 414.350000 1108.500000 415.650000 ;
      RECT 1066.500000 414.350000 1099.500000 415.650000 ;
      RECT 1057.500000 414.350000 1058.500000 415.650000 ;
      RECT 1016.500000 414.350000 1049.500000 415.650000 ;
      RECT 1007.500000 414.350000 1008.500000 415.650000 ;
      RECT 966.500000 414.350000 999.500000 415.650000 ;
      RECT 957.500000 414.350000 958.500000 415.650000 ;
      RECT 916.500000 414.350000 949.500000 415.650000 ;
      RECT 907.500000 414.350000 908.500000 415.650000 ;
      RECT 866.500000 414.350000 899.500000 415.650000 ;
      RECT 857.500000 414.350000 858.500000 415.650000 ;
      RECT 816.500000 414.350000 849.500000 415.650000 ;
      RECT 807.500000 414.350000 808.500000 415.650000 ;
      RECT 766.500000 414.350000 799.500000 415.650000 ;
      RECT 757.500000 414.350000 758.500000 415.650000 ;
      RECT 720.000000 414.350000 749.500000 415.650000 ;
      RECT 707.500000 414.350000 712.000000 415.650000 ;
      RECT 666.500000 414.350000 699.500000 415.650000 ;
      RECT 657.500000 414.350000 658.500000 415.650000 ;
      RECT 616.500000 414.350000 649.500000 415.650000 ;
      RECT 607.500000 414.350000 608.500000 415.650000 ;
      RECT 566.500000 414.350000 599.500000 415.650000 ;
      RECT 557.500000 414.350000 558.500000 415.650000 ;
      RECT 516.500000 414.350000 549.500000 415.650000 ;
      RECT 507.500000 414.350000 508.500000 415.650000 ;
      RECT 416.500000 414.350000 499.500000 415.650000 ;
      RECT 407.500000 414.350000 408.500000 415.650000 ;
      RECT 366.500000 414.350000 399.500000 415.650000 ;
      RECT 357.500000 414.350000 358.500000 415.650000 ;
      RECT 316.500000 414.350000 349.500000 415.650000 ;
      RECT 307.500000 414.350000 308.500000 415.650000 ;
      RECT 216.500000 414.350000 299.500000 415.650000 ;
      RECT 207.500000 414.350000 208.500000 415.650000 ;
      RECT 116.500000 414.350000 199.500000 415.650000 ;
      RECT 107.500000 414.350000 108.500000 415.650000 ;
      RECT 66.500000 414.350000 99.500000 415.650000 ;
      RECT 57.500000 414.350000 58.500000 415.650000 ;
      RECT 29.500000 414.350000 49.500000 415.650000 ;
      RECT 15.500000 414.350000 16.500000 415.650000 ;
      RECT 1157.500000 413.650000 1170.500000 414.350000 ;
      RECT 1107.500000 413.650000 1149.500000 414.350000 ;
      RECT 1057.500000 413.650000 1099.500000 414.350000 ;
      RECT 1007.500000 413.650000 1049.500000 414.350000 ;
      RECT 957.500000 413.650000 999.500000 414.350000 ;
      RECT 907.500000 413.650000 949.500000 414.350000 ;
      RECT 857.500000 413.650000 899.500000 414.350000 ;
      RECT 807.500000 413.650000 849.500000 414.350000 ;
      RECT 757.500000 413.650000 799.500000 414.350000 ;
      RECT 707.500000 413.650000 749.500000 414.350000 ;
      RECT 657.500000 413.650000 699.500000 414.350000 ;
      RECT 607.500000 413.650000 649.500000 414.350000 ;
      RECT 557.500000 413.650000 599.500000 414.350000 ;
      RECT 507.500000 413.650000 549.500000 414.350000 ;
      RECT 407.500000 413.650000 499.500000 414.350000 ;
      RECT 357.500000 413.650000 399.500000 414.350000 ;
      RECT 307.500000 413.650000 349.500000 414.350000 ;
      RECT 207.500000 413.650000 299.500000 414.350000 ;
      RECT 107.500000 413.650000 199.500000 414.350000 ;
      RECT 57.500000 413.650000 99.500000 414.350000 ;
      RECT 15.500000 413.650000 49.500000 414.350000 ;
      RECT 1183.500000 412.350000 1186.000000 415.650000 ;
      RECT 1169.500000 412.350000 1170.500000 413.650000 ;
      RECT 1116.500000 412.350000 1149.500000 413.650000 ;
      RECT 1107.500000 412.350000 1108.500000 413.650000 ;
      RECT 1066.500000 412.350000 1099.500000 413.650000 ;
      RECT 1057.500000 412.350000 1058.500000 413.650000 ;
      RECT 1016.500000 412.350000 1049.500000 413.650000 ;
      RECT 1007.500000 412.350000 1008.500000 413.650000 ;
      RECT 966.500000 412.350000 999.500000 413.650000 ;
      RECT 957.500000 412.350000 958.500000 413.650000 ;
      RECT 916.500000 412.350000 949.500000 413.650000 ;
      RECT 907.500000 412.350000 908.500000 413.650000 ;
      RECT 866.500000 412.350000 899.500000 413.650000 ;
      RECT 857.500000 412.350000 858.500000 413.650000 ;
      RECT 816.500000 412.350000 849.500000 413.650000 ;
      RECT 807.500000 412.350000 808.500000 413.650000 ;
      RECT 766.500000 412.350000 799.500000 413.650000 ;
      RECT 757.500000 412.350000 758.500000 413.650000 ;
      RECT 720.000000 412.350000 749.500000 413.650000 ;
      RECT 707.500000 412.350000 708.500000 413.650000 ;
      RECT 666.500000 412.350000 699.500000 413.650000 ;
      RECT 657.500000 412.350000 658.500000 413.650000 ;
      RECT 616.500000 412.350000 649.500000 413.650000 ;
      RECT 607.500000 412.350000 608.500000 413.650000 ;
      RECT 566.500000 412.350000 599.500000 413.650000 ;
      RECT 557.500000 412.350000 558.500000 413.650000 ;
      RECT 516.500000 412.350000 549.500000 413.650000 ;
      RECT 507.500000 412.350000 508.500000 413.650000 ;
      RECT 416.500000 412.350000 499.500000 413.650000 ;
      RECT 407.500000 412.350000 408.500000 413.650000 ;
      RECT 366.500000 412.350000 399.500000 413.650000 ;
      RECT 357.500000 412.350000 358.500000 413.650000 ;
      RECT 316.500000 412.350000 349.500000 413.650000 ;
      RECT 307.500000 412.350000 308.500000 413.650000 ;
      RECT 216.500000 412.350000 299.500000 413.650000 ;
      RECT 207.500000 412.350000 208.500000 413.650000 ;
      RECT 116.500000 412.350000 199.500000 413.650000 ;
      RECT 107.500000 412.350000 108.500000 413.650000 ;
      RECT 66.500000 412.350000 99.500000 413.650000 ;
      RECT 57.500000 412.350000 58.500000 413.650000 ;
      RECT 29.500000 412.350000 49.500000 413.650000 ;
      RECT 15.500000 412.350000 16.500000 413.650000 ;
      RECT 0.000000 412.350000 2.500000 415.650000 ;
      RECT 1169.500000 411.650000 1186.000000 412.350000 ;
      RECT 1116.500000 411.650000 1156.500000 412.350000 ;
      RECT 1066.500000 411.650000 1108.500000 412.350000 ;
      RECT 1016.500000 411.650000 1058.500000 412.350000 ;
      RECT 966.500000 411.650000 1008.500000 412.350000 ;
      RECT 916.500000 411.650000 958.500000 412.350000 ;
      RECT 866.500000 411.650000 908.500000 412.350000 ;
      RECT 816.500000 411.650000 858.500000 412.350000 ;
      RECT 766.500000 411.650000 808.500000 412.350000 ;
      RECT 720.000000 411.650000 758.500000 412.350000 ;
      RECT 666.500000 411.650000 708.500000 412.350000 ;
      RECT 616.500000 411.650000 658.500000 412.350000 ;
      RECT 566.500000 411.650000 608.500000 412.350000 ;
      RECT 516.500000 411.650000 558.500000 412.350000 ;
      RECT 416.500000 411.650000 508.500000 412.350000 ;
      RECT 366.500000 411.650000 408.500000 412.350000 ;
      RECT 316.500000 411.650000 358.500000 412.350000 ;
      RECT 216.500000 411.650000 308.500000 412.350000 ;
      RECT 116.500000 411.650000 208.500000 412.350000 ;
      RECT 66.500000 411.650000 108.500000 412.350000 ;
      RECT 29.500000 411.650000 58.500000 412.350000 ;
      RECT 0.000000 411.650000 16.500000 412.350000 ;
      RECT 1169.500000 410.350000 1170.500000 411.650000 ;
      RECT 1116.500000 410.350000 1149.500000 411.650000 ;
      RECT 1107.500000 410.350000 1108.500000 411.650000 ;
      RECT 1066.500000 410.350000 1099.500000 411.650000 ;
      RECT 1057.500000 410.350000 1058.500000 411.650000 ;
      RECT 1016.500000 410.350000 1049.500000 411.650000 ;
      RECT 1007.500000 410.350000 1008.500000 411.650000 ;
      RECT 966.500000 410.350000 999.500000 411.650000 ;
      RECT 957.500000 410.350000 958.500000 411.650000 ;
      RECT 916.500000 410.350000 949.500000 411.650000 ;
      RECT 907.500000 410.350000 908.500000 411.650000 ;
      RECT 866.500000 410.350000 899.500000 411.650000 ;
      RECT 857.500000 410.350000 858.500000 411.650000 ;
      RECT 816.500000 410.350000 849.500000 411.650000 ;
      RECT 807.500000 410.350000 808.500000 411.650000 ;
      RECT 766.500000 410.350000 799.500000 411.650000 ;
      RECT 757.500000 410.350000 758.500000 411.650000 ;
      RECT 720.000000 410.350000 749.500000 411.650000 ;
      RECT 707.500000 410.350000 708.500000 411.650000 ;
      RECT 666.500000 410.350000 699.500000 411.650000 ;
      RECT 657.500000 410.350000 658.500000 411.650000 ;
      RECT 616.500000 410.350000 649.500000 411.650000 ;
      RECT 607.500000 410.350000 608.500000 411.650000 ;
      RECT 566.500000 410.350000 599.500000 411.650000 ;
      RECT 557.500000 410.350000 558.500000 411.650000 ;
      RECT 516.500000 410.350000 549.500000 411.650000 ;
      RECT 507.500000 410.350000 508.500000 411.650000 ;
      RECT 416.500000 410.350000 499.500000 411.650000 ;
      RECT 407.500000 410.350000 408.500000 411.650000 ;
      RECT 366.500000 410.350000 399.500000 411.650000 ;
      RECT 357.500000 410.350000 358.500000 411.650000 ;
      RECT 316.500000 410.350000 349.500000 411.650000 ;
      RECT 307.500000 410.350000 308.500000 411.650000 ;
      RECT 216.500000 410.350000 299.500000 411.650000 ;
      RECT 207.500000 410.350000 208.500000 411.650000 ;
      RECT 116.500000 410.350000 199.500000 411.650000 ;
      RECT 107.500000 410.350000 108.500000 411.650000 ;
      RECT 66.500000 410.350000 99.500000 411.650000 ;
      RECT 57.500000 410.350000 58.500000 411.650000 ;
      RECT 29.500000 410.350000 49.500000 411.650000 ;
      RECT 15.500000 410.350000 16.500000 411.650000 ;
      RECT 1157.500000 409.650000 1170.500000 410.350000 ;
      RECT 1107.500000 409.650000 1149.500000 410.350000 ;
      RECT 1057.500000 409.650000 1099.500000 410.350000 ;
      RECT 1007.500000 409.650000 1049.500000 410.350000 ;
      RECT 957.500000 409.650000 999.500000 410.350000 ;
      RECT 907.500000 409.650000 949.500000 410.350000 ;
      RECT 857.500000 409.650000 899.500000 410.350000 ;
      RECT 807.500000 409.650000 849.500000 410.350000 ;
      RECT 757.500000 409.650000 799.500000 410.350000 ;
      RECT 707.500000 409.650000 749.500000 410.350000 ;
      RECT 657.500000 409.650000 699.500000 410.350000 ;
      RECT 607.500000 409.650000 649.500000 410.350000 ;
      RECT 557.500000 409.650000 599.500000 410.350000 ;
      RECT 507.500000 409.650000 549.500000 410.350000 ;
      RECT 407.500000 409.650000 499.500000 410.350000 ;
      RECT 357.500000 409.650000 399.500000 410.350000 ;
      RECT 307.500000 409.650000 349.500000 410.350000 ;
      RECT 207.500000 409.650000 299.500000 410.350000 ;
      RECT 107.500000 409.650000 199.500000 410.350000 ;
      RECT 57.500000 409.650000 99.500000 410.350000 ;
      RECT 15.500000 409.650000 49.500000 410.350000 ;
      RECT 1183.500000 408.350000 1186.000000 411.650000 ;
      RECT 1169.500000 408.350000 1170.500000 409.650000 ;
      RECT 1116.500000 408.350000 1149.500000 409.650000 ;
      RECT 1107.500000 408.350000 1108.500000 409.650000 ;
      RECT 1066.500000 408.350000 1099.500000 409.650000 ;
      RECT 1057.500000 408.350000 1058.500000 409.650000 ;
      RECT 1016.500000 408.350000 1049.500000 409.650000 ;
      RECT 1007.500000 408.350000 1008.500000 409.650000 ;
      RECT 966.500000 408.350000 999.500000 409.650000 ;
      RECT 957.500000 408.350000 958.500000 409.650000 ;
      RECT 916.500000 408.350000 949.500000 409.650000 ;
      RECT 907.500000 408.350000 908.500000 409.650000 ;
      RECT 866.500000 408.350000 899.500000 409.650000 ;
      RECT 857.500000 408.350000 858.500000 409.650000 ;
      RECT 816.500000 408.350000 849.500000 409.650000 ;
      RECT 807.500000 408.350000 808.500000 409.650000 ;
      RECT 766.500000 408.350000 799.500000 409.650000 ;
      RECT 757.500000 408.350000 758.500000 409.650000 ;
      RECT 716.500000 408.350000 749.500000 409.650000 ;
      RECT 707.500000 408.350000 708.500000 409.650000 ;
      RECT 666.500000 408.350000 699.500000 409.650000 ;
      RECT 657.500000 408.350000 658.500000 409.650000 ;
      RECT 616.500000 408.350000 649.500000 409.650000 ;
      RECT 607.500000 408.350000 608.500000 409.650000 ;
      RECT 566.500000 408.350000 599.500000 409.650000 ;
      RECT 557.500000 408.350000 558.500000 409.650000 ;
      RECT 516.500000 408.350000 549.500000 409.650000 ;
      RECT 507.500000 408.350000 508.500000 409.650000 ;
      RECT 416.500000 408.350000 499.500000 409.650000 ;
      RECT 407.500000 408.350000 408.500000 409.650000 ;
      RECT 366.500000 408.350000 399.500000 409.650000 ;
      RECT 357.500000 408.350000 358.500000 409.650000 ;
      RECT 316.500000 408.350000 349.500000 409.650000 ;
      RECT 307.500000 408.350000 308.500000 409.650000 ;
      RECT 216.500000 408.350000 299.500000 409.650000 ;
      RECT 207.500000 408.350000 208.500000 409.650000 ;
      RECT 116.500000 408.350000 199.500000 409.650000 ;
      RECT 107.500000 408.350000 108.500000 409.650000 ;
      RECT 66.500000 408.350000 99.500000 409.650000 ;
      RECT 57.500000 408.350000 58.500000 409.650000 ;
      RECT 29.500000 408.350000 49.500000 409.650000 ;
      RECT 15.500000 408.350000 16.500000 409.650000 ;
      RECT 0.000000 408.350000 2.500000 411.650000 ;
      RECT 1169.500000 407.650000 1186.000000 408.350000 ;
      RECT 1116.500000 407.650000 1156.500000 408.350000 ;
      RECT 1066.500000 407.650000 1108.500000 408.350000 ;
      RECT 1016.500000 407.650000 1058.500000 408.350000 ;
      RECT 966.500000 407.650000 1008.500000 408.350000 ;
      RECT 916.500000 407.650000 958.500000 408.350000 ;
      RECT 866.500000 407.650000 908.500000 408.350000 ;
      RECT 816.500000 407.650000 858.500000 408.350000 ;
      RECT 766.500000 407.650000 808.500000 408.350000 ;
      RECT 716.500000 407.650000 758.500000 408.350000 ;
      RECT 666.500000 407.650000 708.500000 408.350000 ;
      RECT 616.500000 407.650000 658.500000 408.350000 ;
      RECT 566.500000 407.650000 608.500000 408.350000 ;
      RECT 516.500000 407.650000 558.500000 408.350000 ;
      RECT 416.500000 407.650000 508.500000 408.350000 ;
      RECT 366.500000 407.650000 408.500000 408.350000 ;
      RECT 316.500000 407.650000 358.500000 408.350000 ;
      RECT 216.500000 407.650000 308.500000 408.350000 ;
      RECT 116.500000 407.650000 208.500000 408.350000 ;
      RECT 66.500000 407.650000 108.500000 408.350000 ;
      RECT 29.500000 407.650000 58.500000 408.350000 ;
      RECT 0.000000 407.650000 16.500000 408.350000 ;
      RECT 1169.500000 406.350000 1170.500000 407.650000 ;
      RECT 1116.500000 406.350000 1149.500000 407.650000 ;
      RECT 1107.500000 406.350000 1108.500000 407.650000 ;
      RECT 1066.500000 406.350000 1099.500000 407.650000 ;
      RECT 1057.500000 406.350000 1058.500000 407.650000 ;
      RECT 1016.500000 406.350000 1049.500000 407.650000 ;
      RECT 1007.500000 406.350000 1008.500000 407.650000 ;
      RECT 966.500000 406.350000 999.500000 407.650000 ;
      RECT 957.500000 406.350000 958.500000 407.650000 ;
      RECT 916.500000 406.350000 949.500000 407.650000 ;
      RECT 907.500000 406.350000 908.500000 407.650000 ;
      RECT 866.500000 406.350000 899.500000 407.650000 ;
      RECT 857.500000 406.350000 858.500000 407.650000 ;
      RECT 816.500000 406.350000 849.500000 407.650000 ;
      RECT 807.500000 406.350000 808.500000 407.650000 ;
      RECT 766.500000 406.350000 799.500000 407.650000 ;
      RECT 757.500000 406.350000 758.500000 407.650000 ;
      RECT 716.500000 406.350000 749.500000 407.650000 ;
      RECT 707.500000 406.350000 708.500000 407.650000 ;
      RECT 666.500000 406.350000 699.500000 407.650000 ;
      RECT 657.500000 406.350000 658.500000 407.650000 ;
      RECT 616.500000 406.350000 649.500000 407.650000 ;
      RECT 607.500000 406.350000 608.500000 407.650000 ;
      RECT 566.500000 406.350000 599.500000 407.650000 ;
      RECT 557.500000 406.350000 558.500000 407.650000 ;
      RECT 516.500000 406.350000 549.500000 407.650000 ;
      RECT 507.500000 406.350000 508.500000 407.650000 ;
      RECT 416.500000 406.350000 499.500000 407.650000 ;
      RECT 407.500000 406.350000 408.500000 407.650000 ;
      RECT 366.500000 406.350000 399.500000 407.650000 ;
      RECT 357.500000 406.350000 358.500000 407.650000 ;
      RECT 316.500000 406.350000 349.500000 407.650000 ;
      RECT 307.500000 406.350000 308.500000 407.650000 ;
      RECT 216.500000 406.350000 299.500000 407.650000 ;
      RECT 207.500000 406.350000 208.500000 407.650000 ;
      RECT 116.500000 406.350000 199.500000 407.650000 ;
      RECT 107.500000 406.350000 108.500000 407.650000 ;
      RECT 66.500000 406.350000 99.500000 407.650000 ;
      RECT 57.500000 406.350000 58.500000 407.650000 ;
      RECT 29.500000 406.350000 49.500000 407.650000 ;
      RECT 15.500000 406.350000 16.500000 407.650000 ;
      RECT 1157.500000 405.650000 1170.500000 406.350000 ;
      RECT 1107.500000 405.650000 1149.500000 406.350000 ;
      RECT 1057.500000 405.650000 1099.500000 406.350000 ;
      RECT 1007.500000 405.650000 1049.500000 406.350000 ;
      RECT 957.500000 405.650000 999.500000 406.350000 ;
      RECT 907.500000 405.650000 949.500000 406.350000 ;
      RECT 857.500000 405.650000 899.500000 406.350000 ;
      RECT 807.500000 405.650000 849.500000 406.350000 ;
      RECT 757.500000 405.650000 799.500000 406.350000 ;
      RECT 707.500000 405.650000 749.500000 406.350000 ;
      RECT 657.500000 405.650000 699.500000 406.350000 ;
      RECT 607.500000 405.650000 649.500000 406.350000 ;
      RECT 557.500000 405.650000 599.500000 406.350000 ;
      RECT 507.500000 405.650000 549.500000 406.350000 ;
      RECT 407.500000 405.650000 499.500000 406.350000 ;
      RECT 357.500000 405.650000 399.500000 406.350000 ;
      RECT 307.500000 405.650000 349.500000 406.350000 ;
      RECT 207.500000 405.650000 299.500000 406.350000 ;
      RECT 107.500000 405.650000 199.500000 406.350000 ;
      RECT 57.500000 405.650000 99.500000 406.350000 ;
      RECT 15.500000 405.650000 49.500000 406.350000 ;
      RECT 1183.500000 404.350000 1186.000000 407.650000 ;
      RECT 1169.500000 404.350000 1170.500000 405.650000 ;
      RECT 1116.500000 404.350000 1149.500000 405.650000 ;
      RECT 1107.500000 404.350000 1108.500000 405.650000 ;
      RECT 1066.500000 404.350000 1099.500000 405.650000 ;
      RECT 1057.500000 404.350000 1058.500000 405.650000 ;
      RECT 1016.500000 404.350000 1049.500000 405.650000 ;
      RECT 1007.500000 404.350000 1008.500000 405.650000 ;
      RECT 966.500000 404.350000 999.500000 405.650000 ;
      RECT 957.500000 404.350000 958.500000 405.650000 ;
      RECT 916.500000 404.350000 949.500000 405.650000 ;
      RECT 907.500000 404.350000 908.500000 405.650000 ;
      RECT 866.500000 404.350000 899.500000 405.650000 ;
      RECT 857.500000 404.350000 858.500000 405.650000 ;
      RECT 816.500000 404.350000 849.500000 405.650000 ;
      RECT 807.500000 404.350000 808.500000 405.650000 ;
      RECT 766.500000 404.350000 799.500000 405.650000 ;
      RECT 757.500000 404.350000 758.500000 405.650000 ;
      RECT 716.500000 404.350000 749.500000 405.650000 ;
      RECT 707.500000 404.350000 708.500000 405.650000 ;
      RECT 666.500000 404.350000 699.500000 405.650000 ;
      RECT 657.500000 404.350000 658.500000 405.650000 ;
      RECT 616.500000 404.350000 649.500000 405.650000 ;
      RECT 607.500000 404.350000 608.500000 405.650000 ;
      RECT 566.500000 404.350000 599.500000 405.650000 ;
      RECT 557.500000 404.350000 558.500000 405.650000 ;
      RECT 516.500000 404.350000 549.500000 405.650000 ;
      RECT 507.500000 404.350000 508.500000 405.650000 ;
      RECT 416.500000 404.350000 499.500000 405.650000 ;
      RECT 407.500000 404.350000 408.500000 405.650000 ;
      RECT 366.500000 404.350000 399.500000 405.650000 ;
      RECT 357.500000 404.350000 358.500000 405.650000 ;
      RECT 316.500000 404.350000 349.500000 405.650000 ;
      RECT 307.500000 404.350000 308.500000 405.650000 ;
      RECT 216.500000 404.350000 299.500000 405.650000 ;
      RECT 207.500000 404.350000 208.500000 405.650000 ;
      RECT 116.500000 404.350000 199.500000 405.650000 ;
      RECT 107.500000 404.350000 108.500000 405.650000 ;
      RECT 66.500000 404.350000 99.500000 405.650000 ;
      RECT 57.500000 404.350000 58.500000 405.650000 ;
      RECT 29.500000 404.350000 49.500000 405.650000 ;
      RECT 15.500000 404.350000 16.500000 405.650000 ;
      RECT 0.000000 404.350000 2.500000 407.650000 ;
      RECT 1169.500000 403.650000 1186.000000 404.350000 ;
      RECT 1116.500000 403.650000 1156.500000 404.350000 ;
      RECT 1066.500000 403.650000 1108.500000 404.350000 ;
      RECT 1016.500000 403.650000 1058.500000 404.350000 ;
      RECT 966.500000 403.650000 1008.500000 404.350000 ;
      RECT 916.500000 403.650000 958.500000 404.350000 ;
      RECT 866.500000 403.650000 908.500000 404.350000 ;
      RECT 816.500000 403.650000 858.500000 404.350000 ;
      RECT 766.500000 403.650000 808.500000 404.350000 ;
      RECT 716.500000 403.650000 758.500000 404.350000 ;
      RECT 666.500000 403.650000 708.500000 404.350000 ;
      RECT 616.500000 403.650000 658.500000 404.350000 ;
      RECT 566.500000 403.650000 608.500000 404.350000 ;
      RECT 516.500000 403.650000 558.500000 404.350000 ;
      RECT 416.500000 403.650000 508.500000 404.350000 ;
      RECT 366.500000 403.650000 408.500000 404.350000 ;
      RECT 316.500000 403.650000 358.500000 404.350000 ;
      RECT 216.500000 403.650000 308.500000 404.350000 ;
      RECT 116.500000 403.650000 208.500000 404.350000 ;
      RECT 66.500000 403.650000 108.500000 404.350000 ;
      RECT 29.500000 403.650000 58.500000 404.350000 ;
      RECT 0.000000 403.650000 16.500000 404.350000 ;
      RECT 1169.500000 402.350000 1170.500000 403.650000 ;
      RECT 1116.500000 402.350000 1149.500000 403.650000 ;
      RECT 1107.500000 402.350000 1108.500000 403.650000 ;
      RECT 1066.500000 402.350000 1099.500000 403.650000 ;
      RECT 1057.500000 402.350000 1058.500000 403.650000 ;
      RECT 1016.500000 402.350000 1049.500000 403.650000 ;
      RECT 1007.500000 402.350000 1008.500000 403.650000 ;
      RECT 966.500000 402.350000 999.500000 403.650000 ;
      RECT 957.500000 402.350000 958.500000 403.650000 ;
      RECT 916.500000 402.350000 949.500000 403.650000 ;
      RECT 907.500000 402.350000 908.500000 403.650000 ;
      RECT 866.500000 402.350000 899.500000 403.650000 ;
      RECT 857.500000 402.350000 858.500000 403.650000 ;
      RECT 816.500000 402.350000 849.500000 403.650000 ;
      RECT 807.500000 402.350000 808.500000 403.650000 ;
      RECT 766.500000 402.350000 799.500000 403.650000 ;
      RECT 757.500000 402.350000 758.500000 403.650000 ;
      RECT 716.500000 402.350000 749.500000 403.650000 ;
      RECT 707.500000 402.350000 708.500000 403.650000 ;
      RECT 666.500000 402.350000 699.500000 403.650000 ;
      RECT 657.500000 402.350000 658.500000 403.650000 ;
      RECT 616.500000 402.350000 649.500000 403.650000 ;
      RECT 607.500000 402.350000 608.500000 403.650000 ;
      RECT 566.500000 402.350000 599.500000 403.650000 ;
      RECT 557.500000 402.350000 558.500000 403.650000 ;
      RECT 516.500000 402.350000 549.500000 403.650000 ;
      RECT 507.500000 402.350000 508.500000 403.650000 ;
      RECT 416.500000 402.350000 499.500000 403.650000 ;
      RECT 407.500000 402.350000 408.500000 403.650000 ;
      RECT 366.500000 402.350000 399.500000 403.650000 ;
      RECT 357.500000 402.350000 358.500000 403.650000 ;
      RECT 316.500000 402.350000 349.500000 403.650000 ;
      RECT 307.500000 402.350000 308.500000 403.650000 ;
      RECT 216.500000 402.350000 249.500000 403.650000 ;
      RECT 207.500000 402.350000 208.500000 403.650000 ;
      RECT 116.500000 402.350000 149.500000 403.650000 ;
      RECT 107.500000 402.350000 108.500000 403.650000 ;
      RECT 66.500000 402.350000 99.500000 403.650000 ;
      RECT 57.500000 402.350000 58.500000 403.650000 ;
      RECT 29.500000 402.350000 49.500000 403.650000 ;
      RECT 15.500000 402.350000 16.500000 403.650000 ;
      RECT 1157.500000 401.650000 1170.500000 402.350000 ;
      RECT 1107.500000 401.650000 1149.500000 402.350000 ;
      RECT 1057.500000 401.650000 1099.500000 402.350000 ;
      RECT 1007.500000 401.650000 1049.500000 402.350000 ;
      RECT 957.500000 401.650000 999.500000 402.350000 ;
      RECT 907.500000 401.650000 949.500000 402.350000 ;
      RECT 857.500000 401.650000 899.500000 402.350000 ;
      RECT 807.500000 401.650000 849.500000 402.350000 ;
      RECT 757.500000 401.650000 799.500000 402.350000 ;
      RECT 707.500000 401.650000 749.500000 402.350000 ;
      RECT 657.500000 401.650000 699.500000 402.350000 ;
      RECT 607.500000 401.650000 649.500000 402.350000 ;
      RECT 557.500000 401.650000 599.500000 402.350000 ;
      RECT 507.500000 401.650000 549.500000 402.350000 ;
      RECT 407.500000 401.650000 499.500000 402.350000 ;
      RECT 357.500000 401.650000 399.500000 402.350000 ;
      RECT 307.500000 401.650000 349.500000 402.350000 ;
      RECT 257.500000 401.650000 299.500000 403.650000 ;
      RECT 207.500000 401.650000 249.500000 402.350000 ;
      RECT 157.500000 401.650000 199.500000 403.650000 ;
      RECT 107.500000 401.650000 149.500000 402.350000 ;
      RECT 57.500000 401.650000 99.500000 402.350000 ;
      RECT 15.500000 401.650000 49.500000 402.350000 ;
      RECT 1183.500000 400.350000 1186.000000 403.650000 ;
      RECT 1169.500000 400.350000 1170.500000 401.650000 ;
      RECT 1116.500000 400.350000 1149.500000 401.650000 ;
      RECT 1107.500000 400.350000 1108.500000 401.650000 ;
      RECT 1066.500000 400.350000 1099.500000 401.650000 ;
      RECT 1057.500000 400.350000 1058.500000 401.650000 ;
      RECT 1016.500000 400.350000 1049.500000 401.650000 ;
      RECT 1007.500000 400.350000 1008.500000 401.650000 ;
      RECT 966.500000 400.350000 999.500000 401.650000 ;
      RECT 957.500000 400.350000 958.500000 401.650000 ;
      RECT 916.500000 400.350000 949.500000 401.650000 ;
      RECT 907.500000 400.350000 908.500000 401.650000 ;
      RECT 866.500000 400.350000 899.500000 401.650000 ;
      RECT 857.500000 400.350000 858.500000 401.650000 ;
      RECT 816.500000 400.350000 849.500000 401.650000 ;
      RECT 807.500000 400.350000 808.500000 401.650000 ;
      RECT 766.500000 400.350000 799.500000 401.650000 ;
      RECT 757.500000 400.350000 758.500000 401.650000 ;
      RECT 716.500000 400.350000 749.500000 401.650000 ;
      RECT 707.500000 400.350000 708.500000 401.650000 ;
      RECT 666.500000 400.350000 699.500000 401.650000 ;
      RECT 657.500000 400.350000 658.500000 401.650000 ;
      RECT 616.500000 400.350000 649.500000 401.650000 ;
      RECT 607.500000 400.350000 608.500000 401.650000 ;
      RECT 566.500000 400.350000 599.500000 401.650000 ;
      RECT 557.500000 400.350000 558.500000 401.650000 ;
      RECT 516.500000 400.350000 549.500000 401.650000 ;
      RECT 507.500000 400.350000 508.500000 401.650000 ;
      RECT 416.500000 400.350000 499.500000 401.650000 ;
      RECT 407.500000 400.350000 408.500000 401.650000 ;
      RECT 366.500000 400.350000 399.500000 401.650000 ;
      RECT 357.500000 400.350000 358.500000 401.650000 ;
      RECT 316.500000 400.350000 349.500000 401.650000 ;
      RECT 307.500000 400.350000 308.500000 401.650000 ;
      RECT 266.500000 400.350000 299.500000 401.650000 ;
      RECT 257.500000 400.350000 258.500000 401.650000 ;
      RECT 216.500000 400.350000 249.500000 401.650000 ;
      RECT 207.500000 400.350000 208.500000 401.650000 ;
      RECT 166.500000 400.350000 199.500000 401.650000 ;
      RECT 157.500000 400.350000 158.500000 401.650000 ;
      RECT 116.500000 400.350000 149.500000 401.650000 ;
      RECT 107.500000 400.350000 108.500000 401.650000 ;
      RECT 66.500000 400.350000 99.500000 401.650000 ;
      RECT 57.500000 400.350000 58.500000 401.650000 ;
      RECT 29.500000 400.350000 49.500000 401.650000 ;
      RECT 15.500000 400.350000 16.500000 401.650000 ;
      RECT 0.000000 400.350000 2.500000 403.650000 ;
      RECT 1169.500000 399.650000 1186.000000 400.350000 ;
      RECT 1116.500000 399.650000 1156.500000 400.350000 ;
      RECT 1066.500000 399.650000 1108.500000 400.350000 ;
      RECT 1016.500000 399.650000 1058.500000 400.350000 ;
      RECT 966.500000 399.650000 1008.500000 400.350000 ;
      RECT 916.500000 399.650000 958.500000 400.350000 ;
      RECT 866.500000 399.650000 908.500000 400.350000 ;
      RECT 816.500000 399.650000 858.500000 400.350000 ;
      RECT 766.500000 399.650000 808.500000 400.350000 ;
      RECT 716.500000 399.650000 758.500000 400.350000 ;
      RECT 666.500000 399.650000 708.500000 400.350000 ;
      RECT 616.500000 399.650000 658.500000 400.350000 ;
      RECT 566.500000 399.650000 608.500000 400.350000 ;
      RECT 516.500000 399.650000 558.500000 400.350000 ;
      RECT 416.500000 399.650000 508.500000 400.350000 ;
      RECT 366.500000 399.650000 408.500000 400.350000 ;
      RECT 316.500000 399.650000 358.500000 400.350000 ;
      RECT 266.500000 399.650000 308.500000 400.350000 ;
      RECT 216.500000 399.650000 258.500000 400.350000 ;
      RECT 166.500000 399.650000 208.500000 400.350000 ;
      RECT 116.500000 399.650000 158.500000 400.350000 ;
      RECT 66.500000 399.650000 108.500000 400.350000 ;
      RECT 29.500000 399.650000 58.500000 400.350000 ;
      RECT 0.000000 399.650000 16.500000 400.350000 ;
      RECT 0.000000 399.170000 2.500000 399.650000 ;
      RECT 1183.500000 399.165000 1186.000000 399.650000 ;
      RECT 1169.500000 398.350000 1170.500000 399.650000 ;
      RECT 1116.500000 398.350000 1149.500000 399.650000 ;
      RECT 1107.500000 398.350000 1108.500000 399.650000 ;
      RECT 1066.500000 398.350000 1099.500000 399.650000 ;
      RECT 1057.500000 398.350000 1058.500000 399.650000 ;
      RECT 1016.500000 398.350000 1049.500000 399.650000 ;
      RECT 1007.500000 398.350000 1008.500000 399.650000 ;
      RECT 966.500000 398.350000 999.500000 399.650000 ;
      RECT 957.500000 398.350000 958.500000 399.650000 ;
      RECT 916.500000 398.350000 949.500000 399.650000 ;
      RECT 907.500000 398.350000 908.500000 399.650000 ;
      RECT 866.500000 398.350000 899.500000 399.650000 ;
      RECT 857.500000 398.350000 858.500000 399.650000 ;
      RECT 816.500000 398.350000 849.500000 399.650000 ;
      RECT 807.500000 398.350000 808.500000 399.650000 ;
      RECT 766.500000 398.350000 799.500000 399.650000 ;
      RECT 757.500000 398.350000 758.500000 399.650000 ;
      RECT 716.500000 398.350000 749.500000 399.650000 ;
      RECT 707.500000 398.350000 708.500000 399.650000 ;
      RECT 666.500000 398.350000 699.500000 399.650000 ;
      RECT 657.500000 398.350000 658.500000 399.650000 ;
      RECT 616.500000 398.350000 649.500000 399.650000 ;
      RECT 607.500000 398.350000 608.500000 399.650000 ;
      RECT 566.500000 398.350000 599.500000 399.650000 ;
      RECT 557.500000 398.350000 558.500000 399.650000 ;
      RECT 516.500000 398.350000 549.500000 399.650000 ;
      RECT 507.500000 398.350000 508.500000 399.650000 ;
      RECT 416.500000 398.350000 449.500000 399.650000 ;
      RECT 407.500000 398.350000 408.500000 399.650000 ;
      RECT 366.500000 398.350000 399.500000 399.650000 ;
      RECT 357.500000 398.350000 358.500000 399.650000 ;
      RECT 316.500000 398.350000 349.500000 399.650000 ;
      RECT 307.500000 398.350000 308.500000 399.650000 ;
      RECT 266.500000 398.350000 299.500000 399.650000 ;
      RECT 257.500000 398.350000 258.500000 399.650000 ;
      RECT 216.500000 398.350000 249.500000 399.650000 ;
      RECT 207.500000 398.350000 208.500000 399.650000 ;
      RECT 166.500000 398.350000 199.500000 399.650000 ;
      RECT 157.500000 398.350000 158.500000 399.650000 ;
      RECT 116.500000 398.350000 149.500000 399.650000 ;
      RECT 107.500000 398.350000 108.500000 399.650000 ;
      RECT 66.500000 398.350000 99.500000 399.650000 ;
      RECT 57.500000 398.350000 58.500000 399.650000 ;
      RECT 29.500000 398.350000 49.500000 399.650000 ;
      RECT 15.500000 398.350000 16.500000 399.650000 ;
      RECT 1157.500000 397.650000 1170.500000 398.350000 ;
      RECT 1107.500000 397.650000 1149.500000 398.350000 ;
      RECT 1057.500000 397.650000 1099.500000 398.350000 ;
      RECT 1007.500000 397.650000 1049.500000 398.350000 ;
      RECT 957.500000 397.650000 999.500000 398.350000 ;
      RECT 907.500000 397.650000 949.500000 398.350000 ;
      RECT 857.500000 397.650000 899.500000 398.350000 ;
      RECT 807.500000 397.650000 849.500000 398.350000 ;
      RECT 757.500000 397.650000 799.500000 398.350000 ;
      RECT 707.500000 397.650000 749.500000 398.350000 ;
      RECT 657.500000 397.650000 699.500000 398.350000 ;
      RECT 607.500000 397.650000 649.500000 398.350000 ;
      RECT 557.500000 397.650000 599.500000 398.350000 ;
      RECT 507.500000 397.650000 549.500000 398.350000 ;
      RECT 457.500000 397.650000 499.500000 399.650000 ;
      RECT 407.500000 397.650000 449.500000 398.350000 ;
      RECT 357.500000 397.650000 399.500000 398.350000 ;
      RECT 307.500000 397.650000 349.500000 398.350000 ;
      RECT 257.500000 397.650000 299.500000 398.350000 ;
      RECT 207.500000 397.650000 249.500000 398.350000 ;
      RECT 157.500000 397.650000 199.500000 398.350000 ;
      RECT 107.500000 397.650000 149.500000 398.350000 ;
      RECT 57.500000 397.650000 99.500000 398.350000 ;
      RECT 15.500000 397.650000 49.500000 398.350000 ;
      RECT 1183.500000 396.350000 1183.980000 399.165000 ;
      RECT 1169.500000 396.350000 1170.500000 397.650000 ;
      RECT 1116.500000 396.350000 1149.500000 397.650000 ;
      RECT 1107.500000 396.350000 1108.500000 397.650000 ;
      RECT 1066.500000 396.350000 1099.500000 397.650000 ;
      RECT 1057.500000 396.350000 1058.500000 397.650000 ;
      RECT 1016.500000 396.350000 1049.500000 397.650000 ;
      RECT 1007.500000 396.350000 1008.500000 397.650000 ;
      RECT 966.500000 396.350000 999.500000 397.650000 ;
      RECT 957.500000 396.350000 958.500000 397.650000 ;
      RECT 916.500000 396.350000 949.500000 397.650000 ;
      RECT 907.500000 396.350000 908.500000 397.650000 ;
      RECT 866.500000 396.350000 899.500000 397.650000 ;
      RECT 857.500000 396.350000 858.500000 397.650000 ;
      RECT 816.500000 396.350000 849.500000 397.650000 ;
      RECT 807.500000 396.350000 808.500000 397.650000 ;
      RECT 766.500000 396.350000 799.500000 397.650000 ;
      RECT 757.500000 396.350000 758.500000 397.650000 ;
      RECT 716.500000 396.350000 749.500000 397.650000 ;
      RECT 707.500000 396.350000 708.500000 397.650000 ;
      RECT 666.500000 396.350000 699.500000 397.650000 ;
      RECT 657.500000 396.350000 658.500000 397.650000 ;
      RECT 616.500000 396.350000 649.500000 397.650000 ;
      RECT 607.500000 396.350000 608.500000 397.650000 ;
      RECT 566.500000 396.350000 599.500000 397.650000 ;
      RECT 557.500000 396.350000 558.500000 397.650000 ;
      RECT 516.500000 396.350000 549.500000 397.650000 ;
      RECT 507.500000 396.350000 508.500000 397.650000 ;
      RECT 466.500000 396.350000 499.500000 397.650000 ;
      RECT 457.500000 396.350000 458.500000 397.650000 ;
      RECT 416.500000 396.350000 449.500000 397.650000 ;
      RECT 407.500000 396.350000 408.500000 397.650000 ;
      RECT 366.500000 396.350000 399.500000 397.650000 ;
      RECT 357.500000 396.350000 358.500000 397.650000 ;
      RECT 316.500000 396.350000 349.500000 397.650000 ;
      RECT 307.500000 396.350000 308.500000 397.650000 ;
      RECT 266.500000 396.350000 299.500000 397.650000 ;
      RECT 257.500000 396.350000 258.500000 397.650000 ;
      RECT 216.500000 396.350000 249.500000 397.650000 ;
      RECT 207.500000 396.350000 208.500000 397.650000 ;
      RECT 166.500000 396.350000 199.500000 397.650000 ;
      RECT 157.500000 396.350000 158.500000 397.650000 ;
      RECT 116.500000 396.350000 149.500000 397.650000 ;
      RECT 107.500000 396.350000 108.500000 397.650000 ;
      RECT 66.500000 396.350000 99.500000 397.650000 ;
      RECT 57.500000 396.350000 58.500000 397.650000 ;
      RECT 29.500000 396.350000 49.500000 397.650000 ;
      RECT 15.500000 396.350000 16.500000 397.650000 ;
      RECT 2.020000 396.350000 2.500000 399.170000 ;
      RECT 2.020000 396.070000 16.500000 396.350000 ;
      RECT 1169.500000 396.065000 1183.980000 396.350000 ;
      RECT 1169.500000 395.650000 1186.000000 396.065000 ;
      RECT 1116.500000 395.650000 1156.500000 396.350000 ;
      RECT 1066.500000 395.650000 1108.500000 396.350000 ;
      RECT 1016.500000 395.650000 1058.500000 396.350000 ;
      RECT 966.500000 395.650000 1008.500000 396.350000 ;
      RECT 916.500000 395.650000 958.500000 396.350000 ;
      RECT 866.500000 395.650000 908.500000 396.350000 ;
      RECT 816.500000 395.650000 858.500000 396.350000 ;
      RECT 766.500000 395.650000 808.500000 396.350000 ;
      RECT 716.500000 395.650000 758.500000 396.350000 ;
      RECT 666.500000 395.650000 708.500000 396.350000 ;
      RECT 616.500000 395.650000 658.500000 396.350000 ;
      RECT 566.500000 395.650000 608.500000 396.350000 ;
      RECT 516.500000 395.650000 558.500000 396.350000 ;
      RECT 466.500000 395.650000 508.500000 396.350000 ;
      RECT 416.500000 395.650000 458.500000 396.350000 ;
      RECT 366.500000 395.650000 408.500000 396.350000 ;
      RECT 316.500000 395.650000 358.500000 396.350000 ;
      RECT 266.500000 395.650000 308.500000 396.350000 ;
      RECT 216.500000 395.650000 258.500000 396.350000 ;
      RECT 166.500000 395.650000 208.500000 396.350000 ;
      RECT 116.500000 395.650000 158.500000 396.350000 ;
      RECT 66.500000 395.650000 108.500000 396.350000 ;
      RECT 29.500000 395.650000 58.500000 396.350000 ;
      RECT 0.000000 395.650000 16.500000 396.070000 ;
      RECT 1169.500000 394.350000 1170.500000 395.650000 ;
      RECT 1116.500000 394.350000 1149.500000 395.650000 ;
      RECT 1107.500000 394.350000 1108.500000 395.650000 ;
      RECT 1066.500000 394.350000 1099.500000 395.650000 ;
      RECT 1057.500000 394.350000 1058.500000 395.650000 ;
      RECT 1016.500000 394.350000 1049.500000 395.650000 ;
      RECT 1007.500000 394.350000 1008.500000 395.650000 ;
      RECT 966.500000 394.350000 999.500000 395.650000 ;
      RECT 957.500000 394.350000 958.500000 395.650000 ;
      RECT 916.500000 394.350000 949.500000 395.650000 ;
      RECT 907.500000 394.350000 908.500000 395.650000 ;
      RECT 866.500000 394.350000 899.500000 395.650000 ;
      RECT 857.500000 394.350000 858.500000 395.650000 ;
      RECT 816.500000 394.350000 849.500000 395.650000 ;
      RECT 807.500000 394.350000 808.500000 395.650000 ;
      RECT 766.500000 394.350000 799.500000 395.650000 ;
      RECT 757.500000 394.350000 758.500000 395.650000 ;
      RECT 716.500000 394.350000 749.500000 395.650000 ;
      RECT 707.500000 394.350000 708.500000 395.650000 ;
      RECT 666.500000 394.350000 699.500000 395.650000 ;
      RECT 657.500000 394.350000 658.500000 395.650000 ;
      RECT 616.500000 394.350000 649.500000 395.650000 ;
      RECT 607.500000 394.350000 608.500000 395.650000 ;
      RECT 566.500000 394.350000 599.500000 395.650000 ;
      RECT 557.500000 394.350000 558.500000 395.650000 ;
      RECT 516.500000 394.350000 549.500000 395.650000 ;
      RECT 507.500000 394.350000 508.500000 395.650000 ;
      RECT 466.500000 394.350000 499.500000 395.650000 ;
      RECT 457.500000 394.350000 458.500000 395.650000 ;
      RECT 416.500000 394.350000 449.500000 395.650000 ;
      RECT 407.500000 394.350000 408.500000 395.650000 ;
      RECT 366.500000 394.350000 399.500000 395.650000 ;
      RECT 357.500000 394.350000 358.500000 395.650000 ;
      RECT 316.500000 394.350000 349.500000 395.650000 ;
      RECT 307.500000 394.350000 308.500000 395.650000 ;
      RECT 266.500000 394.350000 299.500000 395.650000 ;
      RECT 257.500000 394.350000 258.500000 395.650000 ;
      RECT 216.500000 394.350000 249.500000 395.650000 ;
      RECT 207.500000 394.350000 208.500000 395.650000 ;
      RECT 166.500000 394.350000 199.500000 395.650000 ;
      RECT 157.500000 394.350000 158.500000 395.650000 ;
      RECT 116.500000 394.350000 149.500000 395.650000 ;
      RECT 107.500000 394.350000 108.500000 395.650000 ;
      RECT 66.500000 394.350000 99.500000 395.650000 ;
      RECT 57.500000 394.350000 58.500000 395.650000 ;
      RECT 29.500000 394.350000 49.500000 395.650000 ;
      RECT 15.500000 394.350000 16.500000 395.650000 ;
      RECT 1157.500000 393.650000 1170.500000 394.350000 ;
      RECT 1107.500000 393.650000 1149.500000 394.350000 ;
      RECT 1057.500000 393.650000 1099.500000 394.350000 ;
      RECT 1007.500000 393.650000 1049.500000 394.350000 ;
      RECT 957.500000 393.650000 999.500000 394.350000 ;
      RECT 907.500000 393.650000 949.500000 394.350000 ;
      RECT 857.500000 393.650000 899.500000 394.350000 ;
      RECT 807.500000 393.650000 849.500000 394.350000 ;
      RECT 757.500000 393.650000 799.500000 394.350000 ;
      RECT 707.500000 393.650000 749.500000 394.350000 ;
      RECT 657.500000 393.650000 699.500000 394.350000 ;
      RECT 607.500000 393.650000 649.500000 394.350000 ;
      RECT 557.500000 393.650000 599.500000 394.350000 ;
      RECT 507.500000 393.650000 549.500000 394.350000 ;
      RECT 457.500000 393.650000 499.500000 394.350000 ;
      RECT 407.500000 393.650000 449.500000 394.350000 ;
      RECT 357.500000 393.650000 399.500000 394.350000 ;
      RECT 307.500000 393.650000 349.500000 394.350000 ;
      RECT 257.500000 393.650000 299.500000 394.350000 ;
      RECT 207.500000 393.650000 249.500000 394.350000 ;
      RECT 157.500000 393.650000 199.500000 394.350000 ;
      RECT 107.500000 393.650000 149.500000 394.350000 ;
      RECT 57.500000 393.650000 99.500000 394.350000 ;
      RECT 15.500000 393.650000 49.500000 394.350000 ;
      RECT 1183.500000 393.485000 1186.000000 395.650000 ;
      RECT 1183.500000 392.350000 1183.980000 393.485000 ;
      RECT 1169.500000 392.350000 1170.500000 393.650000 ;
      RECT 1116.500000 392.350000 1149.500000 393.650000 ;
      RECT 1107.500000 392.350000 1108.500000 393.650000 ;
      RECT 1066.500000 392.350000 1099.500000 393.650000 ;
      RECT 1057.500000 392.350000 1058.500000 393.650000 ;
      RECT 1016.500000 392.350000 1049.500000 393.650000 ;
      RECT 1007.500000 392.350000 1008.500000 393.650000 ;
      RECT 966.500000 392.350000 999.500000 393.650000 ;
      RECT 957.500000 392.350000 958.500000 393.650000 ;
      RECT 916.500000 392.350000 949.500000 393.650000 ;
      RECT 907.500000 392.350000 908.500000 393.650000 ;
      RECT 866.500000 392.350000 899.500000 393.650000 ;
      RECT 857.500000 392.350000 858.500000 393.650000 ;
      RECT 816.500000 392.350000 849.500000 393.650000 ;
      RECT 807.500000 392.350000 808.500000 393.650000 ;
      RECT 766.500000 392.350000 799.500000 393.650000 ;
      RECT 757.500000 392.350000 758.500000 393.650000 ;
      RECT 716.500000 392.350000 749.500000 393.650000 ;
      RECT 707.500000 392.350000 708.500000 393.650000 ;
      RECT 666.500000 392.350000 699.500000 393.650000 ;
      RECT 657.500000 392.350000 658.500000 393.650000 ;
      RECT 616.500000 392.350000 649.500000 393.650000 ;
      RECT 607.500000 392.350000 608.500000 393.650000 ;
      RECT 566.500000 392.350000 599.500000 393.650000 ;
      RECT 557.500000 392.350000 558.500000 393.650000 ;
      RECT 516.500000 392.350000 549.500000 393.650000 ;
      RECT 507.500000 392.350000 508.500000 393.650000 ;
      RECT 466.500000 392.350000 499.500000 393.650000 ;
      RECT 457.500000 392.350000 458.500000 393.650000 ;
      RECT 416.500000 392.350000 449.500000 393.650000 ;
      RECT 407.500000 392.350000 408.500000 393.650000 ;
      RECT 366.500000 392.350000 399.500000 393.650000 ;
      RECT 357.500000 392.350000 358.500000 393.650000 ;
      RECT 316.500000 392.350000 349.500000 393.650000 ;
      RECT 307.500000 392.350000 308.500000 393.650000 ;
      RECT 266.500000 392.350000 299.500000 393.650000 ;
      RECT 257.500000 392.350000 258.500000 393.650000 ;
      RECT 216.500000 392.350000 249.500000 393.650000 ;
      RECT 207.500000 392.350000 208.500000 393.650000 ;
      RECT 166.500000 392.350000 199.500000 393.650000 ;
      RECT 157.500000 392.350000 158.500000 393.650000 ;
      RECT 116.500000 392.350000 149.500000 393.650000 ;
      RECT 107.500000 392.350000 108.500000 393.650000 ;
      RECT 66.500000 392.350000 99.500000 393.650000 ;
      RECT 57.500000 392.350000 58.500000 393.650000 ;
      RECT 29.500000 392.350000 49.500000 393.650000 ;
      RECT 15.500000 392.350000 16.500000 393.650000 ;
      RECT 0.000000 392.350000 2.500000 395.650000 ;
      RECT 1169.500000 391.650000 1183.980000 392.350000 ;
      RECT 1116.500000 391.650000 1156.500000 392.350000 ;
      RECT 1066.500000 391.650000 1108.500000 392.350000 ;
      RECT 1016.500000 391.650000 1058.500000 392.350000 ;
      RECT 966.500000 391.650000 1008.500000 392.350000 ;
      RECT 916.500000 391.650000 958.500000 392.350000 ;
      RECT 866.500000 391.650000 908.500000 392.350000 ;
      RECT 816.500000 391.650000 858.500000 392.350000 ;
      RECT 766.500000 391.650000 808.500000 392.350000 ;
      RECT 716.500000 391.650000 758.500000 392.350000 ;
      RECT 666.500000 391.650000 708.500000 392.350000 ;
      RECT 616.500000 391.650000 658.500000 392.350000 ;
      RECT 566.500000 391.650000 608.500000 392.350000 ;
      RECT 516.500000 391.650000 558.500000 392.350000 ;
      RECT 466.500000 391.650000 508.500000 392.350000 ;
      RECT 416.500000 391.650000 458.500000 392.350000 ;
      RECT 366.500000 391.650000 408.500000 392.350000 ;
      RECT 316.500000 391.650000 358.500000 392.350000 ;
      RECT 266.500000 391.650000 308.500000 392.350000 ;
      RECT 216.500000 391.650000 258.500000 392.350000 ;
      RECT 166.500000 391.650000 208.500000 392.350000 ;
      RECT 116.500000 391.650000 158.500000 392.350000 ;
      RECT 66.500000 391.650000 108.500000 392.350000 ;
      RECT 29.500000 391.650000 58.500000 392.350000 ;
      RECT 0.000000 391.650000 16.500000 392.350000 ;
      RECT 1183.500000 390.385000 1183.980000 391.650000 ;
      RECT 1169.500000 390.350000 1170.500000 391.650000 ;
      RECT 1116.500000 390.350000 1149.500000 391.650000 ;
      RECT 1107.500000 390.350000 1108.500000 391.650000 ;
      RECT 1066.500000 390.350000 1099.500000 391.650000 ;
      RECT 1057.500000 390.350000 1058.500000 391.650000 ;
      RECT 1016.500000 390.350000 1049.500000 391.650000 ;
      RECT 1007.500000 390.350000 1008.500000 391.650000 ;
      RECT 966.500000 390.350000 999.500000 391.650000 ;
      RECT 957.500000 390.350000 958.500000 391.650000 ;
      RECT 916.500000 390.350000 949.500000 391.650000 ;
      RECT 907.500000 390.350000 908.500000 391.650000 ;
      RECT 866.500000 390.350000 899.500000 391.650000 ;
      RECT 857.500000 390.350000 858.500000 391.650000 ;
      RECT 816.500000 390.350000 849.500000 391.650000 ;
      RECT 807.500000 390.350000 808.500000 391.650000 ;
      RECT 766.500000 390.350000 799.500000 391.650000 ;
      RECT 757.500000 390.350000 758.500000 391.650000 ;
      RECT 716.500000 390.350000 749.500000 391.650000 ;
      RECT 707.500000 390.350000 708.500000 391.650000 ;
      RECT 666.500000 390.350000 699.500000 391.650000 ;
      RECT 657.500000 390.350000 658.500000 391.650000 ;
      RECT 616.500000 390.350000 649.500000 391.650000 ;
      RECT 607.500000 390.350000 608.500000 391.650000 ;
      RECT 566.500000 390.350000 599.500000 391.650000 ;
      RECT 557.500000 390.350000 558.500000 391.650000 ;
      RECT 516.500000 390.350000 549.500000 391.650000 ;
      RECT 507.500000 390.350000 508.500000 391.650000 ;
      RECT 466.500000 390.350000 499.500000 391.650000 ;
      RECT 457.500000 390.350000 458.500000 391.650000 ;
      RECT 416.500000 390.350000 449.500000 391.650000 ;
      RECT 407.500000 390.350000 408.500000 391.650000 ;
      RECT 366.500000 390.350000 399.500000 391.650000 ;
      RECT 357.500000 390.350000 358.500000 391.650000 ;
      RECT 316.500000 390.350000 349.500000 391.650000 ;
      RECT 307.500000 390.350000 308.500000 391.650000 ;
      RECT 266.500000 390.350000 299.500000 391.650000 ;
      RECT 257.500000 390.350000 258.500000 391.650000 ;
      RECT 216.500000 390.350000 249.500000 391.650000 ;
      RECT 207.500000 390.350000 208.500000 391.650000 ;
      RECT 166.500000 390.350000 199.500000 391.650000 ;
      RECT 157.500000 390.350000 158.500000 391.650000 ;
      RECT 116.500000 390.350000 149.500000 391.650000 ;
      RECT 107.500000 390.350000 108.500000 391.650000 ;
      RECT 66.500000 390.350000 99.500000 391.650000 ;
      RECT 57.500000 390.350000 58.500000 391.650000 ;
      RECT 29.500000 390.350000 49.500000 391.650000 ;
      RECT 15.500000 390.350000 16.500000 391.650000 ;
      RECT 1157.500000 389.650000 1170.500000 390.350000 ;
      RECT 1107.500000 389.650000 1149.500000 390.350000 ;
      RECT 1057.500000 389.650000 1099.500000 390.350000 ;
      RECT 1007.500000 389.650000 1049.500000 390.350000 ;
      RECT 957.500000 389.650000 999.500000 390.350000 ;
      RECT 907.500000 389.650000 949.500000 390.350000 ;
      RECT 857.500000 389.650000 899.500000 390.350000 ;
      RECT 807.500000 389.650000 849.500000 390.350000 ;
      RECT 757.500000 389.650000 799.500000 390.350000 ;
      RECT 707.500000 389.650000 749.500000 390.350000 ;
      RECT 657.500000 389.650000 699.500000 390.350000 ;
      RECT 607.500000 389.650000 649.500000 390.350000 ;
      RECT 557.500000 389.650000 599.500000 390.350000 ;
      RECT 507.500000 389.650000 549.500000 390.350000 ;
      RECT 457.500000 389.650000 499.500000 390.350000 ;
      RECT 407.500000 389.650000 449.500000 390.350000 ;
      RECT 357.500000 389.650000 399.500000 390.350000 ;
      RECT 307.500000 389.650000 349.500000 390.350000 ;
      RECT 257.500000 389.650000 299.500000 390.350000 ;
      RECT 207.500000 389.650000 249.500000 390.350000 ;
      RECT 157.500000 389.650000 199.500000 390.350000 ;
      RECT 107.500000 389.650000 149.500000 390.350000 ;
      RECT 57.500000 389.650000 99.500000 390.350000 ;
      RECT 15.500000 389.650000 49.500000 390.350000 ;
      RECT 1183.500000 389.525000 1186.000000 390.385000 ;
      RECT 0.000000 388.575000 2.500000 391.650000 ;
      RECT 1183.500000 388.350000 1183.980000 389.525000 ;
      RECT 1169.500000 388.350000 1170.500000 389.650000 ;
      RECT 1116.500000 388.350000 1149.500000 389.650000 ;
      RECT 1107.500000 388.350000 1108.500000 389.650000 ;
      RECT 1066.500000 388.350000 1099.500000 389.650000 ;
      RECT 1057.500000 388.350000 1058.500000 389.650000 ;
      RECT 1016.500000 388.350000 1049.500000 389.650000 ;
      RECT 1007.500000 388.350000 1008.500000 389.650000 ;
      RECT 966.500000 388.350000 999.500000 389.650000 ;
      RECT 957.500000 388.350000 958.500000 389.650000 ;
      RECT 916.500000 388.350000 949.500000 389.650000 ;
      RECT 907.500000 388.350000 908.500000 389.650000 ;
      RECT 866.500000 388.350000 899.500000 389.650000 ;
      RECT 857.500000 388.350000 858.500000 389.650000 ;
      RECT 816.500000 388.350000 849.500000 389.650000 ;
      RECT 807.500000 388.350000 808.500000 389.650000 ;
      RECT 766.500000 388.350000 799.500000 389.650000 ;
      RECT 757.500000 388.350000 758.500000 389.650000 ;
      RECT 716.500000 388.350000 749.500000 389.650000 ;
      RECT 707.500000 388.350000 708.500000 389.650000 ;
      RECT 666.500000 388.350000 699.500000 389.650000 ;
      RECT 657.500000 388.350000 658.500000 389.650000 ;
      RECT 616.500000 388.350000 649.500000 389.650000 ;
      RECT 607.500000 388.350000 608.500000 389.650000 ;
      RECT 566.500000 388.350000 599.500000 389.650000 ;
      RECT 557.500000 388.350000 558.500000 389.650000 ;
      RECT 516.500000 388.350000 549.500000 389.650000 ;
      RECT 507.500000 388.350000 508.500000 389.650000 ;
      RECT 466.500000 388.350000 499.500000 389.650000 ;
      RECT 457.500000 388.350000 458.500000 389.650000 ;
      RECT 416.500000 388.350000 449.500000 389.650000 ;
      RECT 407.500000 388.350000 408.500000 389.650000 ;
      RECT 366.500000 388.350000 399.500000 389.650000 ;
      RECT 357.500000 388.350000 358.500000 389.650000 ;
      RECT 316.500000 388.350000 349.500000 389.650000 ;
      RECT 307.500000 388.350000 308.500000 389.650000 ;
      RECT 266.500000 388.350000 299.500000 389.650000 ;
      RECT 257.500000 388.350000 258.500000 389.650000 ;
      RECT 216.500000 388.350000 249.500000 389.650000 ;
      RECT 207.500000 388.350000 208.500000 389.650000 ;
      RECT 166.500000 388.350000 199.500000 389.650000 ;
      RECT 157.500000 388.350000 158.500000 389.650000 ;
      RECT 116.500000 388.350000 149.500000 389.650000 ;
      RECT 107.500000 388.350000 108.500000 389.650000 ;
      RECT 66.500000 388.350000 99.500000 389.650000 ;
      RECT 57.500000 388.350000 58.500000 389.650000 ;
      RECT 29.500000 388.350000 49.500000 389.650000 ;
      RECT 15.500000 388.350000 16.500000 389.650000 ;
      RECT 2.020000 388.350000 2.500000 388.575000 ;
      RECT 1169.500000 387.650000 1183.980000 388.350000 ;
      RECT 1116.500000 387.650000 1156.500000 388.350000 ;
      RECT 1066.500000 387.650000 1108.500000 388.350000 ;
      RECT 1016.500000 387.650000 1058.500000 388.350000 ;
      RECT 966.500000 387.650000 1008.500000 388.350000 ;
      RECT 916.500000 387.650000 958.500000 388.350000 ;
      RECT 866.500000 387.650000 908.500000 388.350000 ;
      RECT 816.500000 387.650000 858.500000 388.350000 ;
      RECT 766.500000 387.650000 808.500000 388.350000 ;
      RECT 716.500000 387.650000 758.500000 388.350000 ;
      RECT 666.500000 387.650000 708.500000 388.350000 ;
      RECT 616.500000 387.650000 658.500000 388.350000 ;
      RECT 566.500000 387.650000 608.500000 388.350000 ;
      RECT 516.500000 387.650000 558.500000 388.350000 ;
      RECT 466.500000 387.650000 508.500000 388.350000 ;
      RECT 416.500000 387.650000 458.500000 388.350000 ;
      RECT 366.500000 387.650000 408.500000 388.350000 ;
      RECT 316.500000 387.650000 358.500000 388.350000 ;
      RECT 266.500000 387.650000 308.500000 388.350000 ;
      RECT 216.500000 387.650000 258.500000 388.350000 ;
      RECT 166.500000 387.650000 208.500000 388.350000 ;
      RECT 116.500000 387.650000 158.500000 388.350000 ;
      RECT 66.500000 387.650000 108.500000 388.350000 ;
      RECT 29.500000 387.650000 58.500000 388.350000 ;
      RECT 2.020000 387.650000 16.500000 388.350000 ;
      RECT 1183.500000 386.425000 1183.980000 387.650000 ;
      RECT 1169.500000 386.350000 1170.500000 387.650000 ;
      RECT 1116.500000 386.350000 1149.500000 387.650000 ;
      RECT 1107.500000 386.350000 1108.500000 387.650000 ;
      RECT 1066.500000 386.350000 1099.500000 387.650000 ;
      RECT 1057.500000 386.350000 1058.500000 387.650000 ;
      RECT 1016.500000 386.350000 1049.500000 387.650000 ;
      RECT 1007.500000 386.350000 1008.500000 387.650000 ;
      RECT 966.500000 386.350000 999.500000 387.650000 ;
      RECT 957.500000 386.350000 958.500000 387.650000 ;
      RECT 916.500000 386.350000 949.500000 387.650000 ;
      RECT 907.500000 386.350000 908.500000 387.650000 ;
      RECT 866.500000 386.350000 899.500000 387.650000 ;
      RECT 857.500000 386.350000 858.500000 387.650000 ;
      RECT 816.500000 386.350000 849.500000 387.650000 ;
      RECT 807.500000 386.350000 808.500000 387.650000 ;
      RECT 766.500000 386.350000 799.500000 387.650000 ;
      RECT 757.500000 386.350000 758.500000 387.650000 ;
      RECT 716.500000 386.350000 749.500000 387.650000 ;
      RECT 707.500000 386.350000 708.500000 387.650000 ;
      RECT 666.500000 386.350000 699.500000 387.650000 ;
      RECT 657.500000 386.350000 658.500000 387.650000 ;
      RECT 616.500000 386.350000 649.500000 387.650000 ;
      RECT 607.500000 386.350000 608.500000 387.650000 ;
      RECT 566.500000 386.350000 599.500000 387.650000 ;
      RECT 557.500000 386.350000 558.500000 387.650000 ;
      RECT 516.500000 386.350000 549.500000 387.650000 ;
      RECT 507.500000 386.350000 508.500000 387.650000 ;
      RECT 466.500000 386.350000 499.500000 387.650000 ;
      RECT 457.500000 386.350000 458.500000 387.650000 ;
      RECT 416.500000 386.350000 449.500000 387.650000 ;
      RECT 407.500000 386.350000 408.500000 387.650000 ;
      RECT 366.500000 386.350000 399.500000 387.650000 ;
      RECT 357.500000 386.350000 358.500000 387.650000 ;
      RECT 316.500000 386.350000 349.500000 387.650000 ;
      RECT 307.500000 386.350000 308.500000 387.650000 ;
      RECT 266.500000 386.350000 299.500000 387.650000 ;
      RECT 257.500000 386.350000 258.500000 387.650000 ;
      RECT 216.500000 386.350000 249.500000 387.650000 ;
      RECT 207.500000 386.350000 208.500000 387.650000 ;
      RECT 166.500000 386.350000 199.500000 387.650000 ;
      RECT 157.500000 386.350000 158.500000 387.650000 ;
      RECT 116.500000 386.350000 149.500000 387.650000 ;
      RECT 107.500000 386.350000 108.500000 387.650000 ;
      RECT 66.500000 386.350000 99.500000 387.650000 ;
      RECT 57.500000 386.350000 58.500000 387.650000 ;
      RECT 29.500000 386.350000 49.500000 387.650000 ;
      RECT 15.500000 386.350000 16.500000 387.650000 ;
      RECT 1157.500000 385.650000 1170.500000 386.350000 ;
      RECT 1107.500000 385.650000 1149.500000 386.350000 ;
      RECT 1057.500000 385.650000 1099.500000 386.350000 ;
      RECT 1007.500000 385.650000 1049.500000 386.350000 ;
      RECT 957.500000 385.650000 999.500000 386.350000 ;
      RECT 907.500000 385.650000 949.500000 386.350000 ;
      RECT 857.500000 385.650000 899.500000 386.350000 ;
      RECT 807.500000 385.650000 849.500000 386.350000 ;
      RECT 757.500000 385.650000 799.500000 386.350000 ;
      RECT 707.500000 385.650000 749.500000 386.350000 ;
      RECT 657.500000 385.650000 699.500000 386.350000 ;
      RECT 607.500000 385.650000 649.500000 386.350000 ;
      RECT 557.500000 385.650000 599.500000 386.350000 ;
      RECT 507.500000 385.650000 549.500000 386.350000 ;
      RECT 457.500000 385.650000 499.500000 386.350000 ;
      RECT 407.500000 385.650000 449.500000 386.350000 ;
      RECT 357.500000 385.650000 399.500000 386.350000 ;
      RECT 307.500000 385.650000 349.500000 386.350000 ;
      RECT 257.500000 385.650000 299.500000 386.350000 ;
      RECT 207.500000 385.650000 249.500000 386.350000 ;
      RECT 157.500000 385.650000 199.500000 386.350000 ;
      RECT 107.500000 385.650000 149.500000 386.350000 ;
      RECT 57.500000 385.650000 99.500000 386.350000 ;
      RECT 15.500000 385.650000 49.500000 386.350000 ;
      RECT 2.020000 385.475000 2.500000 387.650000 ;
      RECT 0.000000 384.615000 2.500000 385.475000 ;
      RECT 1183.500000 384.350000 1186.000000 386.425000 ;
      RECT 1169.500000 384.350000 1170.500000 385.650000 ;
      RECT 1116.500000 384.350000 1149.500000 385.650000 ;
      RECT 1107.500000 384.350000 1108.500000 385.650000 ;
      RECT 1066.500000 384.350000 1099.500000 385.650000 ;
      RECT 1057.500000 384.350000 1058.500000 385.650000 ;
      RECT 1016.500000 384.350000 1049.500000 385.650000 ;
      RECT 1007.500000 384.350000 1008.500000 385.650000 ;
      RECT 966.500000 384.350000 999.500000 385.650000 ;
      RECT 957.500000 384.350000 958.500000 385.650000 ;
      RECT 916.500000 384.350000 949.500000 385.650000 ;
      RECT 907.500000 384.350000 908.500000 385.650000 ;
      RECT 866.500000 384.350000 899.500000 385.650000 ;
      RECT 857.500000 384.350000 858.500000 385.650000 ;
      RECT 816.500000 384.350000 849.500000 385.650000 ;
      RECT 807.500000 384.350000 808.500000 385.650000 ;
      RECT 766.500000 384.350000 799.500000 385.650000 ;
      RECT 757.500000 384.350000 758.500000 385.650000 ;
      RECT 716.500000 384.350000 749.500000 385.650000 ;
      RECT 707.500000 384.350000 708.500000 385.650000 ;
      RECT 666.500000 384.350000 699.500000 385.650000 ;
      RECT 657.500000 384.350000 658.500000 385.650000 ;
      RECT 616.500000 384.350000 649.500000 385.650000 ;
      RECT 607.500000 384.350000 608.500000 385.650000 ;
      RECT 566.500000 384.350000 599.500000 385.650000 ;
      RECT 557.500000 384.350000 558.500000 385.650000 ;
      RECT 516.500000 384.350000 549.500000 385.650000 ;
      RECT 507.500000 384.350000 508.500000 385.650000 ;
      RECT 466.500000 384.350000 499.500000 385.650000 ;
      RECT 457.500000 384.350000 458.500000 385.650000 ;
      RECT 416.500000 384.350000 449.500000 385.650000 ;
      RECT 407.500000 384.350000 408.500000 385.650000 ;
      RECT 366.500000 384.350000 399.500000 385.650000 ;
      RECT 357.500000 384.350000 358.500000 385.650000 ;
      RECT 316.500000 384.350000 349.500000 385.650000 ;
      RECT 307.500000 384.350000 308.500000 385.650000 ;
      RECT 266.500000 384.350000 299.500000 385.650000 ;
      RECT 257.500000 384.350000 258.500000 385.650000 ;
      RECT 216.500000 384.350000 249.500000 385.650000 ;
      RECT 207.500000 384.350000 208.500000 385.650000 ;
      RECT 166.500000 384.350000 199.500000 385.650000 ;
      RECT 157.500000 384.350000 158.500000 385.650000 ;
      RECT 116.500000 384.350000 149.500000 385.650000 ;
      RECT 107.500000 384.350000 108.500000 385.650000 ;
      RECT 66.500000 384.350000 99.500000 385.650000 ;
      RECT 57.500000 384.350000 58.500000 385.650000 ;
      RECT 29.500000 384.350000 49.500000 385.650000 ;
      RECT 15.500000 384.350000 16.500000 385.650000 ;
      RECT 2.020000 384.350000 2.500000 384.615000 ;
      RECT 1169.500000 383.650000 1186.000000 384.350000 ;
      RECT 1116.500000 383.650000 1156.500000 384.350000 ;
      RECT 1066.500000 383.650000 1108.500000 384.350000 ;
      RECT 1016.500000 383.650000 1058.500000 384.350000 ;
      RECT 966.500000 383.650000 1008.500000 384.350000 ;
      RECT 916.500000 383.650000 958.500000 384.350000 ;
      RECT 866.500000 383.650000 908.500000 384.350000 ;
      RECT 816.500000 383.650000 858.500000 384.350000 ;
      RECT 766.500000 383.650000 808.500000 384.350000 ;
      RECT 716.500000 383.650000 758.500000 384.350000 ;
      RECT 666.500000 383.650000 708.500000 384.350000 ;
      RECT 616.500000 383.650000 658.500000 384.350000 ;
      RECT 566.500000 383.650000 608.500000 384.350000 ;
      RECT 516.500000 383.650000 558.500000 384.350000 ;
      RECT 466.500000 383.650000 508.500000 384.350000 ;
      RECT 416.500000 383.650000 458.500000 384.350000 ;
      RECT 366.500000 383.650000 408.500000 384.350000 ;
      RECT 316.500000 383.650000 358.500000 384.350000 ;
      RECT 266.500000 383.650000 308.500000 384.350000 ;
      RECT 216.500000 383.650000 258.500000 384.350000 ;
      RECT 166.500000 383.650000 208.500000 384.350000 ;
      RECT 116.500000 383.650000 158.500000 384.350000 ;
      RECT 66.500000 383.650000 108.500000 384.350000 ;
      RECT 29.500000 383.650000 58.500000 384.350000 ;
      RECT 2.020000 383.650000 16.500000 384.350000 ;
      RECT 1169.500000 382.350000 1170.500000 383.650000 ;
      RECT 1116.500000 382.350000 1149.500000 383.650000 ;
      RECT 1107.500000 382.350000 1108.500000 383.650000 ;
      RECT 1066.500000 382.350000 1099.500000 383.650000 ;
      RECT 1057.500000 382.350000 1058.500000 383.650000 ;
      RECT 1016.500000 382.350000 1049.500000 383.650000 ;
      RECT 1007.500000 382.350000 1008.500000 383.650000 ;
      RECT 966.500000 382.350000 999.500000 383.650000 ;
      RECT 957.500000 382.350000 958.500000 383.650000 ;
      RECT 916.500000 382.350000 949.500000 383.650000 ;
      RECT 907.500000 382.350000 908.500000 383.650000 ;
      RECT 866.500000 382.350000 899.500000 383.650000 ;
      RECT 857.500000 382.350000 858.500000 383.650000 ;
      RECT 816.500000 382.350000 849.500000 383.650000 ;
      RECT 807.500000 382.350000 808.500000 383.650000 ;
      RECT 766.500000 382.350000 799.500000 383.650000 ;
      RECT 757.500000 382.350000 758.500000 383.650000 ;
      RECT 716.500000 382.350000 749.500000 383.650000 ;
      RECT 707.500000 382.350000 708.500000 383.650000 ;
      RECT 666.500000 382.350000 699.500000 383.650000 ;
      RECT 657.500000 382.350000 658.500000 383.650000 ;
      RECT 616.500000 382.350000 649.500000 383.650000 ;
      RECT 607.500000 382.350000 608.500000 383.650000 ;
      RECT 566.500000 382.350000 599.500000 383.650000 ;
      RECT 557.500000 382.350000 558.500000 383.650000 ;
      RECT 516.500000 382.350000 549.500000 383.650000 ;
      RECT 507.500000 382.350000 508.500000 383.650000 ;
      RECT 466.500000 382.350000 499.500000 383.650000 ;
      RECT 457.500000 382.350000 458.500000 383.650000 ;
      RECT 416.500000 382.350000 449.500000 383.650000 ;
      RECT 407.500000 382.350000 408.500000 383.650000 ;
      RECT 366.500000 382.350000 399.500000 383.650000 ;
      RECT 357.500000 382.350000 358.500000 383.650000 ;
      RECT 316.500000 382.350000 349.500000 383.650000 ;
      RECT 307.500000 382.350000 308.500000 383.650000 ;
      RECT 266.500000 382.350000 299.500000 383.650000 ;
      RECT 257.500000 382.350000 258.500000 383.650000 ;
      RECT 216.500000 382.350000 249.500000 383.650000 ;
      RECT 207.500000 382.350000 208.500000 383.650000 ;
      RECT 166.500000 382.350000 199.500000 383.650000 ;
      RECT 157.500000 382.350000 158.500000 383.650000 ;
      RECT 116.500000 382.350000 149.500000 383.650000 ;
      RECT 107.500000 382.350000 108.500000 383.650000 ;
      RECT 66.500000 382.350000 99.500000 383.650000 ;
      RECT 57.500000 382.350000 58.500000 383.650000 ;
      RECT 29.500000 382.350000 49.500000 383.650000 ;
      RECT 15.500000 382.350000 16.500000 383.650000 ;
      RECT 1157.500000 381.650000 1170.500000 382.350000 ;
      RECT 1107.500000 381.650000 1149.500000 382.350000 ;
      RECT 1057.500000 381.650000 1099.500000 382.350000 ;
      RECT 1007.500000 381.650000 1049.500000 382.350000 ;
      RECT 957.500000 381.650000 999.500000 382.350000 ;
      RECT 907.500000 381.650000 949.500000 382.350000 ;
      RECT 857.500000 381.650000 899.500000 382.350000 ;
      RECT 807.500000 381.650000 849.500000 382.350000 ;
      RECT 757.500000 381.650000 799.500000 382.350000 ;
      RECT 707.500000 381.650000 749.500000 382.350000 ;
      RECT 657.500000 381.650000 699.500000 382.350000 ;
      RECT 607.500000 381.650000 649.500000 382.350000 ;
      RECT 557.500000 381.650000 599.500000 382.350000 ;
      RECT 507.500000 381.650000 549.500000 382.350000 ;
      RECT 457.500000 381.650000 499.500000 382.350000 ;
      RECT 407.500000 381.650000 449.500000 382.350000 ;
      RECT 357.500000 381.650000 399.500000 382.350000 ;
      RECT 307.500000 381.650000 349.500000 382.350000 ;
      RECT 257.500000 381.650000 299.500000 382.350000 ;
      RECT 207.500000 381.650000 249.500000 382.350000 ;
      RECT 157.500000 381.650000 199.500000 382.350000 ;
      RECT 107.500000 381.650000 149.500000 382.350000 ;
      RECT 57.500000 381.650000 99.500000 382.350000 ;
      RECT 15.500000 381.650000 49.500000 382.350000 ;
      RECT 2.020000 381.515000 2.500000 383.650000 ;
      RECT 1183.500000 380.350000 1186.000000 383.650000 ;
      RECT 1169.500000 380.350000 1170.500000 381.650000 ;
      RECT 1116.500000 380.350000 1149.500000 381.650000 ;
      RECT 1107.500000 380.350000 1108.500000 381.650000 ;
      RECT 1066.500000 380.350000 1099.500000 381.650000 ;
      RECT 1057.500000 380.350000 1058.500000 381.650000 ;
      RECT 1016.500000 380.350000 1049.500000 381.650000 ;
      RECT 1007.500000 380.350000 1008.500000 381.650000 ;
      RECT 966.500000 380.350000 999.500000 381.650000 ;
      RECT 957.500000 380.350000 958.500000 381.650000 ;
      RECT 916.500000 380.350000 949.500000 381.650000 ;
      RECT 907.500000 380.350000 908.500000 381.650000 ;
      RECT 866.500000 380.350000 899.500000 381.650000 ;
      RECT 857.500000 380.350000 858.500000 381.650000 ;
      RECT 816.500000 380.350000 849.500000 381.650000 ;
      RECT 807.500000 380.350000 808.500000 381.650000 ;
      RECT 766.500000 380.350000 799.500000 381.650000 ;
      RECT 757.500000 380.350000 758.500000 381.650000 ;
      RECT 716.500000 380.350000 749.500000 381.650000 ;
      RECT 707.500000 380.350000 708.500000 381.650000 ;
      RECT 666.500000 380.350000 699.500000 381.650000 ;
      RECT 657.500000 380.350000 658.500000 381.650000 ;
      RECT 616.500000 380.350000 649.500000 381.650000 ;
      RECT 607.500000 380.350000 608.500000 381.650000 ;
      RECT 566.500000 380.350000 599.500000 381.650000 ;
      RECT 557.500000 380.350000 558.500000 381.650000 ;
      RECT 516.500000 380.350000 549.500000 381.650000 ;
      RECT 507.500000 380.350000 508.500000 381.650000 ;
      RECT 466.500000 380.350000 499.500000 381.650000 ;
      RECT 457.500000 380.350000 458.500000 381.650000 ;
      RECT 416.500000 380.350000 449.500000 381.650000 ;
      RECT 407.500000 380.350000 408.500000 381.650000 ;
      RECT 366.500000 380.350000 399.500000 381.650000 ;
      RECT 357.500000 380.350000 358.500000 381.650000 ;
      RECT 316.500000 380.350000 349.500000 381.650000 ;
      RECT 307.500000 380.350000 308.500000 381.650000 ;
      RECT 266.500000 380.350000 299.500000 381.650000 ;
      RECT 257.500000 380.350000 258.500000 381.650000 ;
      RECT 216.500000 380.350000 249.500000 381.650000 ;
      RECT 207.500000 380.350000 208.500000 381.650000 ;
      RECT 166.500000 380.350000 199.500000 381.650000 ;
      RECT 157.500000 380.350000 158.500000 381.650000 ;
      RECT 116.500000 380.350000 149.500000 381.650000 ;
      RECT 107.500000 380.350000 108.500000 381.650000 ;
      RECT 66.500000 380.350000 99.500000 381.650000 ;
      RECT 57.500000 380.350000 58.500000 381.650000 ;
      RECT 29.500000 380.350000 49.500000 381.650000 ;
      RECT 15.500000 380.350000 16.500000 381.650000 ;
      RECT 0.000000 380.350000 2.500000 381.515000 ;
      RECT 1169.500000 379.650000 1186.000000 380.350000 ;
      RECT 1116.500000 379.650000 1156.500000 380.350000 ;
      RECT 1066.500000 379.650000 1108.500000 380.350000 ;
      RECT 1016.500000 379.650000 1058.500000 380.350000 ;
      RECT 966.500000 379.650000 1008.500000 380.350000 ;
      RECT 916.500000 379.650000 958.500000 380.350000 ;
      RECT 866.500000 379.650000 908.500000 380.350000 ;
      RECT 816.500000 379.650000 858.500000 380.350000 ;
      RECT 766.500000 379.650000 808.500000 380.350000 ;
      RECT 716.500000 379.650000 758.500000 380.350000 ;
      RECT 666.500000 379.650000 708.500000 380.350000 ;
      RECT 616.500000 379.650000 658.500000 380.350000 ;
      RECT 566.500000 379.650000 608.500000 380.350000 ;
      RECT 516.500000 379.650000 558.500000 380.350000 ;
      RECT 466.500000 379.650000 508.500000 380.350000 ;
      RECT 416.500000 379.650000 458.500000 380.350000 ;
      RECT 366.500000 379.650000 408.500000 380.350000 ;
      RECT 316.500000 379.650000 358.500000 380.350000 ;
      RECT 266.500000 379.650000 308.500000 380.350000 ;
      RECT 216.500000 379.650000 258.500000 380.350000 ;
      RECT 166.500000 379.650000 208.500000 380.350000 ;
      RECT 116.500000 379.650000 158.500000 380.350000 ;
      RECT 66.500000 379.650000 108.500000 380.350000 ;
      RECT 29.500000 379.650000 58.500000 380.350000 ;
      RECT 0.000000 379.650000 16.500000 380.350000 ;
      RECT 0.000000 378.935000 2.500000 379.650000 ;
      RECT 1183.500000 378.930000 1186.000000 379.650000 ;
      RECT 1169.500000 378.350000 1170.500000 379.650000 ;
      RECT 1116.500000 378.350000 1149.500000 379.650000 ;
      RECT 1107.500000 378.350000 1108.500000 379.650000 ;
      RECT 1066.500000 378.350000 1099.500000 379.650000 ;
      RECT 1057.500000 378.350000 1058.500000 379.650000 ;
      RECT 1016.500000 378.350000 1049.500000 379.650000 ;
      RECT 1007.500000 378.350000 1008.500000 379.650000 ;
      RECT 966.500000 378.350000 999.500000 379.650000 ;
      RECT 957.500000 378.350000 958.500000 379.650000 ;
      RECT 916.500000 378.350000 949.500000 379.650000 ;
      RECT 907.500000 378.350000 908.500000 379.650000 ;
      RECT 866.500000 378.350000 899.500000 379.650000 ;
      RECT 857.500000 378.350000 858.500000 379.650000 ;
      RECT 816.500000 378.350000 849.500000 379.650000 ;
      RECT 807.500000 378.350000 808.500000 379.650000 ;
      RECT 766.500000 378.350000 799.500000 379.650000 ;
      RECT 757.500000 378.350000 758.500000 379.650000 ;
      RECT 716.500000 378.350000 749.500000 379.650000 ;
      RECT 707.500000 378.350000 708.500000 379.650000 ;
      RECT 666.500000 378.350000 699.500000 379.650000 ;
      RECT 657.500000 378.350000 658.500000 379.650000 ;
      RECT 616.500000 378.350000 649.500000 379.650000 ;
      RECT 607.500000 378.350000 608.500000 379.650000 ;
      RECT 566.500000 378.350000 599.500000 379.650000 ;
      RECT 557.500000 378.350000 558.500000 379.650000 ;
      RECT 516.500000 378.350000 549.500000 379.650000 ;
      RECT 507.500000 378.350000 508.500000 379.650000 ;
      RECT 466.500000 378.350000 499.500000 379.650000 ;
      RECT 457.500000 378.350000 458.500000 379.650000 ;
      RECT 416.500000 378.350000 449.500000 379.650000 ;
      RECT 407.500000 378.350000 408.500000 379.650000 ;
      RECT 366.500000 378.350000 399.500000 379.650000 ;
      RECT 357.500000 378.350000 358.500000 379.650000 ;
      RECT 316.500000 378.350000 349.500000 379.650000 ;
      RECT 307.500000 378.350000 308.500000 379.650000 ;
      RECT 266.500000 378.350000 299.500000 379.650000 ;
      RECT 257.500000 378.350000 258.500000 379.650000 ;
      RECT 216.500000 378.350000 249.500000 379.650000 ;
      RECT 207.500000 378.350000 208.500000 379.650000 ;
      RECT 166.500000 378.350000 199.500000 379.650000 ;
      RECT 157.500000 378.350000 158.500000 379.650000 ;
      RECT 116.500000 378.350000 149.500000 379.650000 ;
      RECT 107.500000 378.350000 108.500000 379.650000 ;
      RECT 66.500000 378.350000 99.500000 379.650000 ;
      RECT 57.500000 378.350000 58.500000 379.650000 ;
      RECT 29.500000 378.350000 49.500000 379.650000 ;
      RECT 15.500000 378.350000 16.500000 379.650000 ;
      RECT 1157.500000 377.650000 1170.500000 378.350000 ;
      RECT 1107.500000 377.650000 1149.500000 378.350000 ;
      RECT 1057.500000 377.650000 1099.500000 378.350000 ;
      RECT 1007.500000 377.650000 1049.500000 378.350000 ;
      RECT 957.500000 377.650000 999.500000 378.350000 ;
      RECT 907.500000 377.650000 949.500000 378.350000 ;
      RECT 857.500000 377.650000 899.500000 378.350000 ;
      RECT 807.500000 377.650000 849.500000 378.350000 ;
      RECT 757.500000 377.650000 799.500000 378.350000 ;
      RECT 707.500000 377.650000 749.500000 378.350000 ;
      RECT 657.500000 377.650000 699.500000 378.350000 ;
      RECT 607.500000 377.650000 649.500000 378.350000 ;
      RECT 557.500000 377.650000 599.500000 378.350000 ;
      RECT 507.500000 377.650000 549.500000 378.350000 ;
      RECT 457.500000 377.650000 499.500000 378.350000 ;
      RECT 407.500000 377.650000 449.500000 378.350000 ;
      RECT 357.500000 377.650000 399.500000 378.350000 ;
      RECT 307.500000 377.650000 349.500000 378.350000 ;
      RECT 257.500000 377.650000 299.500000 378.350000 ;
      RECT 207.500000 377.650000 249.500000 378.350000 ;
      RECT 157.500000 377.650000 199.500000 378.350000 ;
      RECT 107.500000 377.650000 149.500000 378.350000 ;
      RECT 57.500000 377.650000 99.500000 378.350000 ;
      RECT 15.500000 377.650000 49.500000 378.350000 ;
      RECT 1183.500000 376.350000 1183.980000 378.930000 ;
      RECT 1169.500000 376.350000 1170.500000 377.650000 ;
      RECT 1116.500000 376.350000 1149.500000 377.650000 ;
      RECT 1107.500000 376.350000 1108.500000 377.650000 ;
      RECT 1066.500000 376.350000 1099.500000 377.650000 ;
      RECT 1057.500000 376.350000 1058.500000 377.650000 ;
      RECT 1016.500000 376.350000 1049.500000 377.650000 ;
      RECT 1007.500000 376.350000 1008.500000 377.650000 ;
      RECT 966.500000 376.350000 999.500000 377.650000 ;
      RECT 957.500000 376.350000 958.500000 377.650000 ;
      RECT 916.500000 376.350000 949.500000 377.650000 ;
      RECT 907.500000 376.350000 908.500000 377.650000 ;
      RECT 866.500000 376.350000 899.500000 377.650000 ;
      RECT 857.500000 376.350000 858.500000 377.650000 ;
      RECT 816.500000 376.350000 849.500000 377.650000 ;
      RECT 807.500000 376.350000 808.500000 377.650000 ;
      RECT 766.500000 376.350000 799.500000 377.650000 ;
      RECT 757.500000 376.350000 758.500000 377.650000 ;
      RECT 716.500000 376.350000 749.500000 377.650000 ;
      RECT 707.500000 376.350000 708.500000 377.650000 ;
      RECT 666.500000 376.350000 699.500000 377.650000 ;
      RECT 657.500000 376.350000 658.500000 377.650000 ;
      RECT 616.500000 376.350000 649.500000 377.650000 ;
      RECT 607.500000 376.350000 608.500000 377.650000 ;
      RECT 566.500000 376.350000 599.500000 377.650000 ;
      RECT 557.500000 376.350000 558.500000 377.650000 ;
      RECT 516.500000 376.350000 549.500000 377.650000 ;
      RECT 507.500000 376.350000 508.500000 377.650000 ;
      RECT 466.500000 376.350000 499.500000 377.650000 ;
      RECT 457.500000 376.350000 458.500000 377.650000 ;
      RECT 416.500000 376.350000 449.500000 377.650000 ;
      RECT 407.500000 376.350000 408.500000 377.650000 ;
      RECT 366.500000 376.350000 399.500000 377.650000 ;
      RECT 357.500000 376.350000 358.500000 377.650000 ;
      RECT 316.500000 376.350000 349.500000 377.650000 ;
      RECT 307.500000 376.350000 308.500000 377.650000 ;
      RECT 266.500000 376.350000 299.500000 377.650000 ;
      RECT 257.500000 376.350000 258.500000 377.650000 ;
      RECT 216.500000 376.350000 249.500000 377.650000 ;
      RECT 207.500000 376.350000 208.500000 377.650000 ;
      RECT 166.500000 376.350000 199.500000 377.650000 ;
      RECT 157.500000 376.350000 158.500000 377.650000 ;
      RECT 116.500000 376.350000 149.500000 377.650000 ;
      RECT 107.500000 376.350000 108.500000 377.650000 ;
      RECT 66.500000 376.350000 99.500000 377.650000 ;
      RECT 57.500000 376.350000 58.500000 377.650000 ;
      RECT 29.500000 376.350000 49.500000 377.650000 ;
      RECT 15.500000 376.350000 16.500000 377.650000 ;
      RECT 2.020000 376.350000 2.500000 378.935000 ;
      RECT 2.020000 375.835000 16.500000 376.350000 ;
      RECT 1169.500000 375.830000 1183.980000 376.350000 ;
      RECT 1169.500000 375.650000 1186.000000 375.830000 ;
      RECT 1116.500000 375.650000 1156.500000 376.350000 ;
      RECT 1066.500000 375.650000 1108.500000 376.350000 ;
      RECT 1016.500000 375.650000 1058.500000 376.350000 ;
      RECT 966.500000 375.650000 1008.500000 376.350000 ;
      RECT 916.500000 375.650000 958.500000 376.350000 ;
      RECT 866.500000 375.650000 908.500000 376.350000 ;
      RECT 816.500000 375.650000 858.500000 376.350000 ;
      RECT 766.500000 375.650000 808.500000 376.350000 ;
      RECT 716.500000 375.650000 758.500000 376.350000 ;
      RECT 666.500000 375.650000 708.500000 376.350000 ;
      RECT 616.500000 375.650000 658.500000 376.350000 ;
      RECT 566.500000 375.650000 608.500000 376.350000 ;
      RECT 516.500000 375.650000 558.500000 376.350000 ;
      RECT 466.500000 375.650000 508.500000 376.350000 ;
      RECT 416.500000 375.650000 458.500000 376.350000 ;
      RECT 366.500000 375.650000 408.500000 376.350000 ;
      RECT 316.500000 375.650000 358.500000 376.350000 ;
      RECT 266.500000 375.650000 308.500000 376.350000 ;
      RECT 216.500000 375.650000 258.500000 376.350000 ;
      RECT 166.500000 375.650000 208.500000 376.350000 ;
      RECT 116.500000 375.650000 158.500000 376.350000 ;
      RECT 66.500000 375.650000 108.500000 376.350000 ;
      RECT 29.500000 375.650000 58.500000 376.350000 ;
      RECT 0.000000 375.650000 16.500000 375.835000 ;
      RECT 1169.500000 374.350000 1170.500000 375.650000 ;
      RECT 1116.500000 374.350000 1149.500000 375.650000 ;
      RECT 1107.500000 374.350000 1108.500000 375.650000 ;
      RECT 1066.500000 374.350000 1099.500000 375.650000 ;
      RECT 1057.500000 374.350000 1058.500000 375.650000 ;
      RECT 1016.500000 374.350000 1049.500000 375.650000 ;
      RECT 1007.500000 374.350000 1008.500000 375.650000 ;
      RECT 966.500000 374.350000 999.500000 375.650000 ;
      RECT 957.500000 374.350000 958.500000 375.650000 ;
      RECT 916.500000 374.350000 949.500000 375.650000 ;
      RECT 907.500000 374.350000 908.500000 375.650000 ;
      RECT 866.500000 374.350000 899.500000 375.650000 ;
      RECT 857.500000 374.350000 858.500000 375.650000 ;
      RECT 816.500000 374.350000 849.500000 375.650000 ;
      RECT 807.500000 374.350000 808.500000 375.650000 ;
      RECT 766.500000 374.350000 799.500000 375.650000 ;
      RECT 757.500000 374.350000 758.500000 375.650000 ;
      RECT 716.500000 374.350000 749.500000 375.650000 ;
      RECT 707.500000 374.350000 708.500000 375.650000 ;
      RECT 666.500000 374.350000 699.500000 375.650000 ;
      RECT 657.500000 374.350000 658.500000 375.650000 ;
      RECT 616.500000 374.350000 649.500000 375.650000 ;
      RECT 607.500000 374.350000 608.500000 375.650000 ;
      RECT 566.500000 374.350000 599.500000 375.650000 ;
      RECT 557.500000 374.350000 558.500000 375.650000 ;
      RECT 516.500000 374.350000 549.500000 375.650000 ;
      RECT 507.500000 374.350000 508.500000 375.650000 ;
      RECT 466.500000 374.350000 499.500000 375.650000 ;
      RECT 457.500000 374.350000 458.500000 375.650000 ;
      RECT 416.500000 374.350000 449.500000 375.650000 ;
      RECT 407.500000 374.350000 408.500000 375.650000 ;
      RECT 366.500000 374.350000 399.500000 375.650000 ;
      RECT 357.500000 374.350000 358.500000 375.650000 ;
      RECT 316.500000 374.350000 349.500000 375.650000 ;
      RECT 307.500000 374.350000 308.500000 375.650000 ;
      RECT 266.500000 374.350000 299.500000 375.650000 ;
      RECT 257.500000 374.350000 258.500000 375.650000 ;
      RECT 216.500000 374.350000 249.500000 375.650000 ;
      RECT 207.500000 374.350000 208.500000 375.650000 ;
      RECT 166.500000 374.350000 199.500000 375.650000 ;
      RECT 157.500000 374.350000 158.500000 375.650000 ;
      RECT 116.500000 374.350000 149.500000 375.650000 ;
      RECT 107.500000 374.350000 108.500000 375.650000 ;
      RECT 66.500000 374.350000 99.500000 375.650000 ;
      RECT 57.500000 374.350000 58.500000 375.650000 ;
      RECT 29.500000 374.350000 49.500000 375.650000 ;
      RECT 15.500000 374.350000 16.500000 375.650000 ;
      RECT 1157.500000 373.650000 1170.500000 374.350000 ;
      RECT 1107.500000 373.650000 1149.500000 374.350000 ;
      RECT 1057.500000 373.650000 1099.500000 374.350000 ;
      RECT 1007.500000 373.650000 1049.500000 374.350000 ;
      RECT 957.500000 373.650000 999.500000 374.350000 ;
      RECT 907.500000 373.650000 949.500000 374.350000 ;
      RECT 857.500000 373.650000 899.500000 374.350000 ;
      RECT 807.500000 373.650000 849.500000 374.350000 ;
      RECT 757.500000 373.650000 799.500000 374.350000 ;
      RECT 707.500000 373.650000 749.500000 374.350000 ;
      RECT 657.500000 373.650000 699.500000 374.350000 ;
      RECT 607.500000 373.650000 649.500000 374.350000 ;
      RECT 557.500000 373.650000 599.500000 374.350000 ;
      RECT 507.500000 373.650000 549.500000 374.350000 ;
      RECT 457.500000 373.650000 499.500000 374.350000 ;
      RECT 407.500000 373.650000 449.500000 374.350000 ;
      RECT 357.500000 373.650000 399.500000 374.350000 ;
      RECT 307.500000 373.650000 349.500000 374.350000 ;
      RECT 257.500000 373.650000 299.500000 374.350000 ;
      RECT 207.500000 373.650000 249.500000 374.350000 ;
      RECT 157.500000 373.650000 199.500000 374.350000 ;
      RECT 107.500000 373.650000 149.500000 374.350000 ;
      RECT 57.500000 373.650000 99.500000 374.350000 ;
      RECT 15.500000 373.650000 49.500000 374.350000 ;
      RECT 1183.500000 372.350000 1186.000000 375.650000 ;
      RECT 1169.500000 372.350000 1170.500000 373.650000 ;
      RECT 1116.500000 372.350000 1149.500000 373.650000 ;
      RECT 1107.500000 372.350000 1108.500000 373.650000 ;
      RECT 1066.500000 372.350000 1099.500000 373.650000 ;
      RECT 1057.500000 372.350000 1058.500000 373.650000 ;
      RECT 1016.500000 372.350000 1049.500000 373.650000 ;
      RECT 1007.500000 372.350000 1008.500000 373.650000 ;
      RECT 966.500000 372.350000 999.500000 373.650000 ;
      RECT 957.500000 372.350000 958.500000 373.650000 ;
      RECT 916.500000 372.350000 949.500000 373.650000 ;
      RECT 907.500000 372.350000 908.500000 373.650000 ;
      RECT 866.500000 372.350000 899.500000 373.650000 ;
      RECT 857.500000 372.350000 858.500000 373.650000 ;
      RECT 816.500000 372.350000 849.500000 373.650000 ;
      RECT 807.500000 372.350000 808.500000 373.650000 ;
      RECT 766.500000 372.350000 799.500000 373.650000 ;
      RECT 757.500000 372.350000 758.500000 373.650000 ;
      RECT 716.500000 372.350000 749.500000 373.650000 ;
      RECT 707.500000 372.350000 708.500000 373.650000 ;
      RECT 666.500000 372.350000 699.500000 373.650000 ;
      RECT 657.500000 372.350000 658.500000 373.650000 ;
      RECT 616.500000 372.350000 649.500000 373.650000 ;
      RECT 607.500000 372.350000 608.500000 373.650000 ;
      RECT 566.500000 372.350000 599.500000 373.650000 ;
      RECT 557.500000 372.350000 558.500000 373.650000 ;
      RECT 516.500000 372.350000 549.500000 373.650000 ;
      RECT 507.500000 372.350000 508.500000 373.650000 ;
      RECT 466.500000 372.350000 499.500000 373.650000 ;
      RECT 457.500000 372.350000 458.500000 373.650000 ;
      RECT 416.500000 372.350000 449.500000 373.650000 ;
      RECT 407.500000 372.350000 408.500000 373.650000 ;
      RECT 366.500000 372.350000 399.500000 373.650000 ;
      RECT 357.500000 372.350000 358.500000 373.650000 ;
      RECT 316.500000 372.350000 349.500000 373.650000 ;
      RECT 307.500000 372.350000 308.500000 373.650000 ;
      RECT 266.500000 372.350000 299.500000 373.650000 ;
      RECT 257.500000 372.350000 258.500000 373.650000 ;
      RECT 216.500000 372.350000 249.500000 373.650000 ;
      RECT 207.500000 372.350000 208.500000 373.650000 ;
      RECT 166.500000 372.350000 199.500000 373.650000 ;
      RECT 157.500000 372.350000 158.500000 373.650000 ;
      RECT 116.500000 372.350000 149.500000 373.650000 ;
      RECT 107.500000 372.350000 108.500000 373.650000 ;
      RECT 66.500000 372.350000 99.500000 373.650000 ;
      RECT 57.500000 372.350000 58.500000 373.650000 ;
      RECT 29.500000 372.350000 49.500000 373.650000 ;
      RECT 15.500000 372.350000 16.500000 373.650000 ;
      RECT 0.000000 372.350000 2.500000 375.650000 ;
      RECT 1169.500000 371.650000 1186.000000 372.350000 ;
      RECT 1116.500000 371.650000 1156.500000 372.350000 ;
      RECT 1066.500000 371.650000 1108.500000 372.350000 ;
      RECT 1016.500000 371.650000 1058.500000 372.350000 ;
      RECT 966.500000 371.650000 1008.500000 372.350000 ;
      RECT 916.500000 371.650000 958.500000 372.350000 ;
      RECT 866.500000 371.650000 908.500000 372.350000 ;
      RECT 816.500000 371.650000 858.500000 372.350000 ;
      RECT 766.500000 371.650000 808.500000 372.350000 ;
      RECT 716.500000 371.650000 758.500000 372.350000 ;
      RECT 666.500000 371.650000 708.500000 372.350000 ;
      RECT 616.500000 371.650000 658.500000 372.350000 ;
      RECT 566.500000 371.650000 608.500000 372.350000 ;
      RECT 516.500000 371.650000 558.500000 372.350000 ;
      RECT 466.500000 371.650000 508.500000 372.350000 ;
      RECT 416.500000 371.650000 458.500000 372.350000 ;
      RECT 366.500000 371.650000 408.500000 372.350000 ;
      RECT 316.500000 371.650000 358.500000 372.350000 ;
      RECT 266.500000 371.650000 308.500000 372.350000 ;
      RECT 216.500000 371.650000 258.500000 372.350000 ;
      RECT 166.500000 371.650000 208.500000 372.350000 ;
      RECT 116.500000 371.650000 158.500000 372.350000 ;
      RECT 66.500000 371.650000 108.500000 372.350000 ;
      RECT 29.500000 371.650000 58.500000 372.350000 ;
      RECT 0.000000 371.650000 16.500000 372.350000 ;
      RECT 1169.500000 370.350000 1170.500000 371.650000 ;
      RECT 1116.500000 370.350000 1149.500000 371.650000 ;
      RECT 1107.500000 370.350000 1108.500000 371.650000 ;
      RECT 1066.500000 370.350000 1099.500000 371.650000 ;
      RECT 1057.500000 370.350000 1058.500000 371.650000 ;
      RECT 1016.500000 370.350000 1049.500000 371.650000 ;
      RECT 1007.500000 370.350000 1008.500000 371.650000 ;
      RECT 966.500000 370.350000 999.500000 371.650000 ;
      RECT 957.500000 370.350000 958.500000 371.650000 ;
      RECT 916.500000 370.350000 949.500000 371.650000 ;
      RECT 907.500000 370.350000 908.500000 371.650000 ;
      RECT 866.500000 370.350000 899.500000 371.650000 ;
      RECT 857.500000 370.350000 858.500000 371.650000 ;
      RECT 816.500000 370.350000 849.500000 371.650000 ;
      RECT 807.500000 370.350000 808.500000 371.650000 ;
      RECT 766.500000 370.350000 799.500000 371.650000 ;
      RECT 757.500000 370.350000 758.500000 371.650000 ;
      RECT 716.500000 370.350000 749.500000 371.650000 ;
      RECT 707.500000 370.350000 708.500000 371.650000 ;
      RECT 666.500000 370.350000 699.500000 371.650000 ;
      RECT 657.500000 370.350000 658.500000 371.650000 ;
      RECT 616.500000 370.350000 649.500000 371.650000 ;
      RECT 607.500000 370.350000 608.500000 371.650000 ;
      RECT 566.500000 370.350000 599.500000 371.650000 ;
      RECT 557.500000 370.350000 558.500000 371.650000 ;
      RECT 516.500000 370.350000 549.500000 371.650000 ;
      RECT 507.500000 370.350000 508.500000 371.650000 ;
      RECT 466.500000 370.350000 499.500000 371.650000 ;
      RECT 457.500000 370.350000 458.500000 371.650000 ;
      RECT 416.500000 370.350000 449.500000 371.650000 ;
      RECT 407.500000 370.350000 408.500000 371.650000 ;
      RECT 366.500000 370.350000 399.500000 371.650000 ;
      RECT 357.500000 370.350000 358.500000 371.650000 ;
      RECT 316.500000 370.350000 349.500000 371.650000 ;
      RECT 307.500000 370.350000 308.500000 371.650000 ;
      RECT 266.500000 370.350000 299.500000 371.650000 ;
      RECT 257.500000 370.350000 258.500000 371.650000 ;
      RECT 216.500000 370.350000 249.500000 371.650000 ;
      RECT 207.500000 370.350000 208.500000 371.650000 ;
      RECT 166.500000 370.350000 199.500000 371.650000 ;
      RECT 157.500000 370.350000 158.500000 371.650000 ;
      RECT 116.500000 370.350000 149.500000 371.650000 ;
      RECT 107.500000 370.350000 108.500000 371.650000 ;
      RECT 66.500000 370.350000 99.500000 371.650000 ;
      RECT 57.500000 370.350000 58.500000 371.650000 ;
      RECT 29.500000 370.350000 49.500000 371.650000 ;
      RECT 15.500000 370.350000 16.500000 371.650000 ;
      RECT 1157.500000 369.650000 1170.500000 370.350000 ;
      RECT 1107.500000 369.650000 1149.500000 370.350000 ;
      RECT 1057.500000 369.650000 1099.500000 370.350000 ;
      RECT 1007.500000 369.650000 1049.500000 370.350000 ;
      RECT 957.500000 369.650000 999.500000 370.350000 ;
      RECT 907.500000 369.650000 949.500000 370.350000 ;
      RECT 857.500000 369.650000 899.500000 370.350000 ;
      RECT 807.500000 369.650000 849.500000 370.350000 ;
      RECT 757.500000 369.650000 799.500000 370.350000 ;
      RECT 707.500000 369.650000 749.500000 370.350000 ;
      RECT 657.500000 369.650000 699.500000 370.350000 ;
      RECT 607.500000 369.650000 649.500000 370.350000 ;
      RECT 557.500000 369.650000 599.500000 370.350000 ;
      RECT 507.500000 369.650000 549.500000 370.350000 ;
      RECT 407.500000 369.650000 449.500000 370.350000 ;
      RECT 357.500000 369.650000 399.500000 370.350000 ;
      RECT 307.500000 369.650000 349.500000 370.350000 ;
      RECT 257.500000 369.650000 299.500000 370.350000 ;
      RECT 207.500000 369.650000 249.500000 370.350000 ;
      RECT 157.500000 369.650000 199.500000 370.350000 ;
      RECT 107.500000 369.650000 149.500000 370.350000 ;
      RECT 57.500000 369.650000 99.500000 370.350000 ;
      RECT 15.500000 369.650000 49.500000 370.350000 ;
      RECT 1183.500000 368.350000 1186.000000 371.650000 ;
      RECT 1169.500000 368.350000 1170.500000 369.650000 ;
      RECT 1116.500000 368.350000 1149.500000 369.650000 ;
      RECT 1107.500000 368.350000 1108.500000 369.650000 ;
      RECT 1066.500000 368.350000 1099.500000 369.650000 ;
      RECT 1057.500000 368.350000 1058.500000 369.650000 ;
      RECT 1016.500000 368.350000 1049.500000 369.650000 ;
      RECT 1007.500000 368.350000 1008.500000 369.650000 ;
      RECT 966.500000 368.350000 999.500000 369.650000 ;
      RECT 957.500000 368.350000 958.500000 369.650000 ;
      RECT 916.500000 368.350000 949.500000 369.650000 ;
      RECT 907.500000 368.350000 908.500000 369.650000 ;
      RECT 866.500000 368.350000 899.500000 369.650000 ;
      RECT 857.500000 368.350000 858.500000 369.650000 ;
      RECT 816.500000 368.350000 849.500000 369.650000 ;
      RECT 807.500000 368.350000 808.500000 369.650000 ;
      RECT 766.500000 368.350000 799.500000 369.650000 ;
      RECT 757.500000 368.350000 758.500000 369.650000 ;
      RECT 716.500000 368.350000 749.500000 369.650000 ;
      RECT 707.500000 368.350000 708.500000 369.650000 ;
      RECT 666.500000 368.350000 699.500000 369.650000 ;
      RECT 657.500000 368.350000 658.500000 369.650000 ;
      RECT 616.500000 368.350000 649.500000 369.650000 ;
      RECT 607.500000 368.350000 608.500000 369.650000 ;
      RECT 566.500000 368.350000 599.500000 369.650000 ;
      RECT 557.500000 368.350000 558.500000 369.650000 ;
      RECT 516.500000 368.350000 549.500000 369.650000 ;
      RECT 507.500000 368.350000 508.500000 369.650000 ;
      RECT 457.500000 368.350000 499.500000 370.350000 ;
      RECT 416.500000 368.350000 449.500000 369.650000 ;
      RECT 407.500000 368.350000 408.500000 369.650000 ;
      RECT 366.500000 368.350000 399.500000 369.650000 ;
      RECT 357.500000 368.350000 358.500000 369.650000 ;
      RECT 316.500000 368.350000 349.500000 369.650000 ;
      RECT 307.500000 368.350000 308.500000 369.650000 ;
      RECT 266.500000 368.350000 299.500000 369.650000 ;
      RECT 257.500000 368.350000 258.500000 369.650000 ;
      RECT 216.500000 368.350000 249.500000 369.650000 ;
      RECT 207.500000 368.350000 208.500000 369.650000 ;
      RECT 166.500000 368.350000 199.500000 369.650000 ;
      RECT 157.500000 368.350000 158.500000 369.650000 ;
      RECT 116.500000 368.350000 149.500000 369.650000 ;
      RECT 107.500000 368.350000 108.500000 369.650000 ;
      RECT 66.500000 368.350000 99.500000 369.650000 ;
      RECT 57.500000 368.350000 58.500000 369.650000 ;
      RECT 29.500000 368.350000 49.500000 369.650000 ;
      RECT 15.500000 368.350000 16.500000 369.650000 ;
      RECT 0.000000 368.350000 2.500000 371.650000 ;
      RECT 1169.500000 367.650000 1186.000000 368.350000 ;
      RECT 1116.500000 367.650000 1156.500000 368.350000 ;
      RECT 1066.500000 367.650000 1108.500000 368.350000 ;
      RECT 1016.500000 367.650000 1058.500000 368.350000 ;
      RECT 966.500000 367.650000 1008.500000 368.350000 ;
      RECT 916.500000 367.650000 958.500000 368.350000 ;
      RECT 866.500000 367.650000 908.500000 368.350000 ;
      RECT 816.500000 367.650000 858.500000 368.350000 ;
      RECT 766.500000 367.650000 808.500000 368.350000 ;
      RECT 716.500000 367.650000 758.500000 368.350000 ;
      RECT 666.500000 367.650000 708.500000 368.350000 ;
      RECT 616.500000 367.650000 658.500000 368.350000 ;
      RECT 566.500000 367.650000 608.500000 368.350000 ;
      RECT 516.500000 367.650000 558.500000 368.350000 ;
      RECT 416.500000 367.650000 508.500000 368.350000 ;
      RECT 366.500000 367.650000 408.500000 368.350000 ;
      RECT 316.500000 367.650000 358.500000 368.350000 ;
      RECT 266.500000 367.650000 308.500000 368.350000 ;
      RECT 216.500000 367.650000 258.500000 368.350000 ;
      RECT 166.500000 367.650000 208.500000 368.350000 ;
      RECT 116.500000 367.650000 158.500000 368.350000 ;
      RECT 66.500000 367.650000 108.500000 368.350000 ;
      RECT 29.500000 367.650000 58.500000 368.350000 ;
      RECT 0.000000 367.650000 16.500000 368.350000 ;
      RECT 1169.500000 366.350000 1170.500000 367.650000 ;
      RECT 1116.500000 366.350000 1149.500000 367.650000 ;
      RECT 1107.500000 366.350000 1108.500000 367.650000 ;
      RECT 1066.500000 366.350000 1099.500000 367.650000 ;
      RECT 1057.500000 366.350000 1058.500000 367.650000 ;
      RECT 1016.500000 366.350000 1049.500000 367.650000 ;
      RECT 1007.500000 366.350000 1008.500000 367.650000 ;
      RECT 966.500000 366.350000 999.500000 367.650000 ;
      RECT 957.500000 366.350000 958.500000 367.650000 ;
      RECT 916.500000 366.350000 949.500000 367.650000 ;
      RECT 907.500000 366.350000 908.500000 367.650000 ;
      RECT 866.500000 366.350000 899.500000 367.650000 ;
      RECT 857.500000 366.350000 858.500000 367.650000 ;
      RECT 816.500000 366.350000 849.500000 367.650000 ;
      RECT 807.500000 366.350000 808.500000 367.650000 ;
      RECT 766.500000 366.350000 799.500000 367.650000 ;
      RECT 757.500000 366.350000 758.500000 367.650000 ;
      RECT 716.500000 366.350000 749.500000 367.650000 ;
      RECT 707.500000 366.350000 708.500000 367.650000 ;
      RECT 666.500000 366.350000 699.500000 367.650000 ;
      RECT 657.500000 366.350000 658.500000 367.650000 ;
      RECT 616.500000 366.350000 649.500000 367.650000 ;
      RECT 607.500000 366.350000 608.500000 367.650000 ;
      RECT 566.500000 366.350000 599.500000 367.650000 ;
      RECT 557.500000 366.350000 558.500000 367.650000 ;
      RECT 516.500000 366.350000 549.500000 367.650000 ;
      RECT 507.500000 366.350000 508.500000 367.650000 ;
      RECT 416.500000 366.350000 499.500000 367.650000 ;
      RECT 407.500000 366.350000 408.500000 367.650000 ;
      RECT 366.500000 366.350000 399.500000 367.650000 ;
      RECT 357.500000 366.350000 358.500000 367.650000 ;
      RECT 316.500000 366.350000 349.500000 367.650000 ;
      RECT 307.500000 366.350000 308.500000 367.650000 ;
      RECT 266.500000 366.350000 299.500000 367.650000 ;
      RECT 257.500000 366.350000 258.500000 367.650000 ;
      RECT 216.500000 366.350000 249.500000 367.650000 ;
      RECT 207.500000 366.350000 208.500000 367.650000 ;
      RECT 166.500000 366.350000 199.500000 367.650000 ;
      RECT 157.500000 366.350000 158.500000 367.650000 ;
      RECT 116.500000 366.350000 149.500000 367.650000 ;
      RECT 107.500000 366.350000 108.500000 367.650000 ;
      RECT 66.500000 366.350000 99.500000 367.650000 ;
      RECT 57.500000 366.350000 58.500000 367.650000 ;
      RECT 29.500000 366.350000 49.500000 367.650000 ;
      RECT 15.500000 366.350000 16.500000 367.650000 ;
      RECT 1157.500000 365.650000 1170.500000 366.350000 ;
      RECT 1107.500000 365.650000 1149.500000 366.350000 ;
      RECT 1057.500000 365.650000 1099.500000 366.350000 ;
      RECT 1007.500000 365.650000 1049.500000 366.350000 ;
      RECT 957.500000 365.650000 999.500000 366.350000 ;
      RECT 907.500000 365.650000 949.500000 366.350000 ;
      RECT 857.500000 365.650000 899.500000 366.350000 ;
      RECT 807.500000 365.650000 849.500000 366.350000 ;
      RECT 757.500000 365.650000 799.500000 366.350000 ;
      RECT 707.500000 365.650000 749.500000 366.350000 ;
      RECT 657.500000 365.650000 699.500000 366.350000 ;
      RECT 607.500000 365.650000 649.500000 366.350000 ;
      RECT 557.500000 365.650000 599.500000 366.350000 ;
      RECT 507.500000 365.650000 549.500000 366.350000 ;
      RECT 407.500000 365.650000 499.500000 366.350000 ;
      RECT 357.500000 365.650000 399.500000 366.350000 ;
      RECT 307.500000 365.650000 349.500000 366.350000 ;
      RECT 257.500000 365.650000 299.500000 366.350000 ;
      RECT 207.500000 365.650000 249.500000 366.350000 ;
      RECT 157.500000 365.650000 199.500000 366.350000 ;
      RECT 107.500000 365.650000 149.500000 366.350000 ;
      RECT 57.500000 365.650000 99.500000 366.350000 ;
      RECT 15.500000 365.650000 49.500000 366.350000 ;
      RECT 1183.500000 364.350000 1186.000000 367.650000 ;
      RECT 1169.500000 364.350000 1170.500000 365.650000 ;
      RECT 1116.500000 364.350000 1149.500000 365.650000 ;
      RECT 1107.500000 364.350000 1108.500000 365.650000 ;
      RECT 1066.500000 364.350000 1099.500000 365.650000 ;
      RECT 1057.500000 364.350000 1058.500000 365.650000 ;
      RECT 1016.500000 364.350000 1049.500000 365.650000 ;
      RECT 1007.500000 364.350000 1008.500000 365.650000 ;
      RECT 966.500000 364.350000 999.500000 365.650000 ;
      RECT 957.500000 364.350000 958.500000 365.650000 ;
      RECT 916.500000 364.350000 949.500000 365.650000 ;
      RECT 907.500000 364.350000 908.500000 365.650000 ;
      RECT 866.500000 364.350000 899.500000 365.650000 ;
      RECT 857.500000 364.350000 858.500000 365.650000 ;
      RECT 816.500000 364.350000 849.500000 365.650000 ;
      RECT 807.500000 364.350000 808.500000 365.650000 ;
      RECT 766.500000 364.350000 799.500000 365.650000 ;
      RECT 757.500000 364.350000 758.500000 365.650000 ;
      RECT 716.500000 364.350000 749.500000 365.650000 ;
      RECT 707.500000 364.350000 708.500000 365.650000 ;
      RECT 666.500000 364.350000 699.500000 365.650000 ;
      RECT 657.500000 364.350000 658.500000 365.650000 ;
      RECT 616.500000 364.350000 649.500000 365.650000 ;
      RECT 607.500000 364.350000 608.500000 365.650000 ;
      RECT 566.500000 364.350000 599.500000 365.650000 ;
      RECT 557.500000 364.350000 558.500000 365.650000 ;
      RECT 516.500000 364.350000 549.500000 365.650000 ;
      RECT 507.500000 364.350000 508.500000 365.650000 ;
      RECT 416.500000 364.350000 499.500000 365.650000 ;
      RECT 407.500000 364.350000 408.500000 365.650000 ;
      RECT 366.500000 364.350000 399.500000 365.650000 ;
      RECT 357.500000 364.350000 358.500000 365.650000 ;
      RECT 316.500000 364.350000 349.500000 365.650000 ;
      RECT 307.500000 364.350000 308.500000 365.650000 ;
      RECT 266.500000 364.350000 299.500000 365.650000 ;
      RECT 257.500000 364.350000 258.500000 365.650000 ;
      RECT 216.500000 364.350000 249.500000 365.650000 ;
      RECT 207.500000 364.350000 208.500000 365.650000 ;
      RECT 166.500000 364.350000 199.500000 365.650000 ;
      RECT 157.500000 364.350000 158.500000 365.650000 ;
      RECT 116.500000 364.350000 149.500000 365.650000 ;
      RECT 107.500000 364.350000 108.500000 365.650000 ;
      RECT 66.500000 364.350000 99.500000 365.650000 ;
      RECT 57.500000 364.350000 58.500000 365.650000 ;
      RECT 29.500000 364.350000 49.500000 365.650000 ;
      RECT 15.500000 364.350000 16.500000 365.650000 ;
      RECT 0.000000 364.350000 2.500000 367.650000 ;
      RECT 1169.500000 363.650000 1186.000000 364.350000 ;
      RECT 1116.500000 363.650000 1156.500000 364.350000 ;
      RECT 1066.500000 363.650000 1108.500000 364.350000 ;
      RECT 1016.500000 363.650000 1058.500000 364.350000 ;
      RECT 966.500000 363.650000 1008.500000 364.350000 ;
      RECT 916.500000 363.650000 958.500000 364.350000 ;
      RECT 866.500000 363.650000 908.500000 364.350000 ;
      RECT 816.500000 363.650000 858.500000 364.350000 ;
      RECT 766.500000 363.650000 808.500000 364.350000 ;
      RECT 716.500000 363.650000 758.500000 364.350000 ;
      RECT 666.500000 363.650000 708.500000 364.350000 ;
      RECT 616.500000 363.650000 658.500000 364.350000 ;
      RECT 566.500000 363.650000 608.500000 364.350000 ;
      RECT 516.500000 363.650000 558.500000 364.350000 ;
      RECT 416.500000 363.650000 508.500000 364.350000 ;
      RECT 366.500000 363.650000 408.500000 364.350000 ;
      RECT 316.500000 363.650000 358.500000 364.350000 ;
      RECT 266.500000 363.650000 308.500000 364.350000 ;
      RECT 216.500000 363.650000 258.500000 364.350000 ;
      RECT 166.500000 363.650000 208.500000 364.350000 ;
      RECT 116.500000 363.650000 158.500000 364.350000 ;
      RECT 66.500000 363.650000 108.500000 364.350000 ;
      RECT 29.500000 363.650000 58.500000 364.350000 ;
      RECT 0.000000 363.650000 16.500000 364.350000 ;
      RECT 1169.500000 362.350000 1170.500000 363.650000 ;
      RECT 1116.500000 362.350000 1149.500000 363.650000 ;
      RECT 1107.500000 362.350000 1108.500000 363.650000 ;
      RECT 1066.500000 362.350000 1099.500000 363.650000 ;
      RECT 1057.500000 362.350000 1058.500000 363.650000 ;
      RECT 1016.500000 362.350000 1049.500000 363.650000 ;
      RECT 1007.500000 362.350000 1008.500000 363.650000 ;
      RECT 966.500000 362.350000 999.500000 363.650000 ;
      RECT 957.500000 362.350000 958.500000 363.650000 ;
      RECT 916.500000 362.350000 949.500000 363.650000 ;
      RECT 907.500000 362.350000 908.500000 363.650000 ;
      RECT 866.500000 362.350000 899.500000 363.650000 ;
      RECT 857.500000 362.350000 858.500000 363.650000 ;
      RECT 816.500000 362.350000 849.500000 363.650000 ;
      RECT 807.500000 362.350000 808.500000 363.650000 ;
      RECT 766.500000 362.350000 799.500000 363.650000 ;
      RECT 757.500000 362.350000 758.500000 363.650000 ;
      RECT 716.500000 362.350000 749.500000 363.650000 ;
      RECT 707.500000 362.350000 708.500000 363.650000 ;
      RECT 666.500000 362.350000 699.500000 363.650000 ;
      RECT 657.500000 362.350000 658.500000 363.650000 ;
      RECT 616.500000 362.350000 649.500000 363.650000 ;
      RECT 607.500000 362.350000 608.500000 363.650000 ;
      RECT 566.500000 362.350000 599.500000 363.650000 ;
      RECT 557.500000 362.350000 558.500000 363.650000 ;
      RECT 516.500000 362.350000 549.500000 363.650000 ;
      RECT 507.500000 362.350000 508.500000 363.650000 ;
      RECT 416.500000 362.350000 499.500000 363.650000 ;
      RECT 407.500000 362.350000 408.500000 363.650000 ;
      RECT 366.500000 362.350000 399.500000 363.650000 ;
      RECT 357.500000 362.350000 358.500000 363.650000 ;
      RECT 316.500000 362.350000 349.500000 363.650000 ;
      RECT 307.500000 362.350000 308.500000 363.650000 ;
      RECT 266.500000 362.350000 299.500000 363.650000 ;
      RECT 257.500000 362.350000 258.500000 363.650000 ;
      RECT 216.500000 362.350000 249.500000 363.650000 ;
      RECT 207.500000 362.350000 208.500000 363.650000 ;
      RECT 166.500000 362.350000 199.500000 363.650000 ;
      RECT 157.500000 362.350000 158.500000 363.650000 ;
      RECT 116.500000 362.350000 149.500000 363.650000 ;
      RECT 107.500000 362.350000 108.500000 363.650000 ;
      RECT 66.500000 362.350000 99.500000 363.650000 ;
      RECT 57.500000 362.350000 58.500000 363.650000 ;
      RECT 29.500000 362.350000 49.500000 363.650000 ;
      RECT 15.500000 362.350000 16.500000 363.650000 ;
      RECT 1157.500000 361.650000 1170.500000 362.350000 ;
      RECT 1107.500000 361.650000 1149.500000 362.350000 ;
      RECT 1057.500000 361.650000 1099.500000 362.350000 ;
      RECT 1007.500000 361.650000 1049.500000 362.350000 ;
      RECT 957.500000 361.650000 999.500000 362.350000 ;
      RECT 907.500000 361.650000 949.500000 362.350000 ;
      RECT 857.500000 361.650000 899.500000 362.350000 ;
      RECT 807.500000 361.650000 849.500000 362.350000 ;
      RECT 757.500000 361.650000 799.500000 362.350000 ;
      RECT 707.500000 361.650000 749.500000 362.350000 ;
      RECT 657.500000 361.650000 699.500000 362.350000 ;
      RECT 607.500000 361.650000 649.500000 362.350000 ;
      RECT 557.500000 361.650000 599.500000 362.350000 ;
      RECT 507.500000 361.650000 549.500000 362.350000 ;
      RECT 407.500000 361.650000 499.500000 362.350000 ;
      RECT 357.500000 361.650000 399.500000 362.350000 ;
      RECT 307.500000 361.650000 349.500000 362.350000 ;
      RECT 257.500000 361.650000 299.500000 362.350000 ;
      RECT 207.500000 361.650000 249.500000 362.350000 ;
      RECT 157.500000 361.650000 199.500000 362.350000 ;
      RECT 107.500000 361.650000 149.500000 362.350000 ;
      RECT 15.500000 361.650000 49.500000 362.350000 ;
      RECT 1183.500000 360.350000 1186.000000 363.650000 ;
      RECT 1169.500000 360.350000 1170.500000 361.650000 ;
      RECT 1116.500000 360.350000 1149.500000 361.650000 ;
      RECT 1107.500000 360.350000 1108.500000 361.650000 ;
      RECT 1066.500000 360.350000 1099.500000 361.650000 ;
      RECT 1057.500000 360.350000 1058.500000 361.650000 ;
      RECT 1016.500000 360.350000 1049.500000 361.650000 ;
      RECT 1007.500000 360.350000 1008.500000 361.650000 ;
      RECT 966.500000 360.350000 999.500000 361.650000 ;
      RECT 957.500000 360.350000 958.500000 361.650000 ;
      RECT 916.500000 360.350000 949.500000 361.650000 ;
      RECT 907.500000 360.350000 908.500000 361.650000 ;
      RECT 866.500000 360.350000 899.500000 361.650000 ;
      RECT 857.500000 360.350000 858.500000 361.650000 ;
      RECT 816.500000 360.350000 849.500000 361.650000 ;
      RECT 807.500000 360.350000 808.500000 361.650000 ;
      RECT 766.500000 360.350000 799.500000 361.650000 ;
      RECT 757.500000 360.350000 758.500000 361.650000 ;
      RECT 716.500000 360.350000 749.500000 361.650000 ;
      RECT 707.500000 360.350000 708.500000 361.650000 ;
      RECT 666.500000 360.350000 699.500000 361.650000 ;
      RECT 657.500000 360.350000 658.500000 361.650000 ;
      RECT 616.500000 360.350000 649.500000 361.650000 ;
      RECT 607.500000 360.350000 608.500000 361.650000 ;
      RECT 566.500000 360.350000 599.500000 361.650000 ;
      RECT 557.500000 360.350000 558.500000 361.650000 ;
      RECT 516.500000 360.350000 549.500000 361.650000 ;
      RECT 507.500000 360.350000 508.500000 361.650000 ;
      RECT 416.500000 360.350000 499.500000 361.650000 ;
      RECT 407.500000 360.350000 408.500000 361.650000 ;
      RECT 366.500000 360.350000 399.500000 361.650000 ;
      RECT 357.500000 360.350000 358.500000 361.650000 ;
      RECT 316.500000 360.350000 349.500000 361.650000 ;
      RECT 307.500000 360.350000 308.500000 361.650000 ;
      RECT 266.500000 360.350000 299.500000 361.650000 ;
      RECT 257.500000 360.350000 258.500000 361.650000 ;
      RECT 216.500000 360.350000 249.500000 361.650000 ;
      RECT 207.500000 360.350000 208.500000 361.650000 ;
      RECT 166.500000 360.350000 199.500000 361.650000 ;
      RECT 157.500000 360.350000 158.500000 361.650000 ;
      RECT 116.500000 360.350000 149.500000 361.650000 ;
      RECT 107.500000 360.350000 108.500000 361.650000 ;
      RECT 57.500000 360.350000 99.500000 362.350000 ;
      RECT 29.500000 360.350000 49.500000 361.650000 ;
      RECT 15.500000 360.350000 16.500000 361.650000 ;
      RECT 0.000000 360.350000 2.500000 363.650000 ;
      RECT 1169.500000 359.650000 1186.000000 360.350000 ;
      RECT 1116.500000 359.650000 1156.500000 360.350000 ;
      RECT 1066.500000 359.650000 1108.500000 360.350000 ;
      RECT 1016.500000 359.650000 1058.500000 360.350000 ;
      RECT 966.500000 359.650000 1008.500000 360.350000 ;
      RECT 916.500000 359.650000 958.500000 360.350000 ;
      RECT 866.500000 359.650000 908.500000 360.350000 ;
      RECT 816.500000 359.650000 858.500000 360.350000 ;
      RECT 766.500000 359.650000 808.500000 360.350000 ;
      RECT 716.500000 359.650000 758.500000 360.350000 ;
      RECT 666.500000 359.650000 708.500000 360.350000 ;
      RECT 616.500000 359.650000 658.500000 360.350000 ;
      RECT 566.500000 359.650000 608.500000 360.350000 ;
      RECT 516.500000 359.650000 558.500000 360.350000 ;
      RECT 416.500000 359.650000 508.500000 360.350000 ;
      RECT 366.500000 359.650000 408.500000 360.350000 ;
      RECT 316.500000 359.650000 358.500000 360.350000 ;
      RECT 266.500000 359.650000 308.500000 360.350000 ;
      RECT 216.500000 359.650000 258.500000 360.350000 ;
      RECT 166.500000 359.650000 208.500000 360.350000 ;
      RECT 116.500000 359.650000 158.500000 360.350000 ;
      RECT 29.500000 359.650000 108.500000 360.350000 ;
      RECT 0.000000 359.650000 16.500000 360.350000 ;
      RECT 1169.500000 358.350000 1170.500000 359.650000 ;
      RECT 1116.500000 358.350000 1149.500000 359.650000 ;
      RECT 1107.500000 358.350000 1108.500000 359.650000 ;
      RECT 1066.500000 358.350000 1099.500000 359.650000 ;
      RECT 1057.500000 358.350000 1058.500000 359.650000 ;
      RECT 1016.500000 358.350000 1049.500000 359.650000 ;
      RECT 1007.500000 358.350000 1008.500000 359.650000 ;
      RECT 966.500000 358.350000 999.500000 359.650000 ;
      RECT 957.500000 358.350000 958.500000 359.650000 ;
      RECT 916.500000 358.350000 949.500000 359.650000 ;
      RECT 907.500000 358.350000 908.500000 359.650000 ;
      RECT 866.500000 358.350000 899.500000 359.650000 ;
      RECT 857.500000 358.350000 858.500000 359.650000 ;
      RECT 816.500000 358.350000 849.500000 359.650000 ;
      RECT 807.500000 358.350000 808.500000 359.650000 ;
      RECT 766.500000 358.350000 799.500000 359.650000 ;
      RECT 757.500000 358.350000 758.500000 359.650000 ;
      RECT 716.500000 358.350000 749.500000 359.650000 ;
      RECT 707.500000 358.350000 708.500000 359.650000 ;
      RECT 666.500000 358.350000 699.500000 359.650000 ;
      RECT 657.500000 358.350000 658.500000 359.650000 ;
      RECT 616.500000 358.350000 649.500000 359.650000 ;
      RECT 607.500000 358.350000 608.500000 359.650000 ;
      RECT 566.500000 358.350000 599.500000 359.650000 ;
      RECT 557.500000 358.350000 558.500000 359.650000 ;
      RECT 516.500000 358.350000 549.500000 359.650000 ;
      RECT 507.500000 358.350000 508.500000 359.650000 ;
      RECT 416.500000 358.350000 499.500000 359.650000 ;
      RECT 407.500000 358.350000 408.500000 359.650000 ;
      RECT 366.500000 358.350000 399.500000 359.650000 ;
      RECT 357.500000 358.350000 358.500000 359.650000 ;
      RECT 316.500000 358.350000 349.500000 359.650000 ;
      RECT 307.500000 358.350000 308.500000 359.650000 ;
      RECT 266.500000 358.350000 299.500000 359.650000 ;
      RECT 257.500000 358.350000 258.500000 359.650000 ;
      RECT 216.500000 358.350000 249.500000 359.650000 ;
      RECT 207.500000 358.350000 208.500000 359.650000 ;
      RECT 166.500000 358.350000 199.500000 359.650000 ;
      RECT 157.500000 358.350000 158.500000 359.650000 ;
      RECT 116.500000 358.350000 149.500000 359.650000 ;
      RECT 107.500000 358.350000 108.500000 359.650000 ;
      RECT 29.500000 358.350000 99.500000 359.650000 ;
      RECT 15.500000 358.350000 16.500000 359.650000 ;
      RECT 1157.500000 357.650000 1170.500000 358.350000 ;
      RECT 1107.500000 357.650000 1149.500000 358.350000 ;
      RECT 1057.500000 357.650000 1099.500000 358.350000 ;
      RECT 1007.500000 357.650000 1049.500000 358.350000 ;
      RECT 957.500000 357.650000 999.500000 358.350000 ;
      RECT 907.500000 357.650000 949.500000 358.350000 ;
      RECT 857.500000 357.650000 899.500000 358.350000 ;
      RECT 807.500000 357.650000 849.500000 358.350000 ;
      RECT 757.500000 357.650000 799.500000 358.350000 ;
      RECT 707.500000 357.650000 749.500000 358.350000 ;
      RECT 657.500000 357.650000 699.500000 358.350000 ;
      RECT 607.500000 357.650000 649.500000 358.350000 ;
      RECT 557.500000 357.650000 599.500000 358.350000 ;
      RECT 507.500000 357.650000 549.500000 358.350000 ;
      RECT 407.500000 357.650000 499.500000 358.350000 ;
      RECT 357.500000 357.650000 399.500000 358.350000 ;
      RECT 307.500000 357.650000 349.500000 358.350000 ;
      RECT 257.500000 357.650000 299.500000 358.350000 ;
      RECT 207.500000 357.650000 249.500000 358.350000 ;
      RECT 157.500000 357.650000 199.500000 358.350000 ;
      RECT 107.500000 357.650000 149.500000 358.350000 ;
      RECT 15.500000 357.650000 99.500000 358.350000 ;
      RECT 1183.500000 356.350000 1186.000000 359.650000 ;
      RECT 1169.500000 356.350000 1170.500000 357.650000 ;
      RECT 1116.500000 356.350000 1149.500000 357.650000 ;
      RECT 1107.500000 356.350000 1108.500000 357.650000 ;
      RECT 1066.500000 356.350000 1099.500000 357.650000 ;
      RECT 1057.500000 356.350000 1058.500000 357.650000 ;
      RECT 1016.500000 356.350000 1049.500000 357.650000 ;
      RECT 1007.500000 356.350000 1008.500000 357.650000 ;
      RECT 966.500000 356.350000 999.500000 357.650000 ;
      RECT 957.500000 356.350000 958.500000 357.650000 ;
      RECT 916.500000 356.350000 949.500000 357.650000 ;
      RECT 907.500000 356.350000 908.500000 357.650000 ;
      RECT 866.500000 356.350000 899.500000 357.650000 ;
      RECT 857.500000 356.350000 858.500000 357.650000 ;
      RECT 816.500000 356.350000 849.500000 357.650000 ;
      RECT 807.500000 356.350000 808.500000 357.650000 ;
      RECT 766.500000 356.350000 799.500000 357.650000 ;
      RECT 757.500000 356.350000 758.500000 357.650000 ;
      RECT 716.500000 356.350000 749.500000 357.650000 ;
      RECT 707.500000 356.350000 708.500000 357.650000 ;
      RECT 666.500000 356.350000 699.500000 357.650000 ;
      RECT 657.500000 356.350000 658.500000 357.650000 ;
      RECT 616.500000 356.350000 649.500000 357.650000 ;
      RECT 607.500000 356.350000 608.500000 357.650000 ;
      RECT 566.500000 356.350000 599.500000 357.650000 ;
      RECT 557.500000 356.350000 558.500000 357.650000 ;
      RECT 516.500000 356.350000 549.500000 357.650000 ;
      RECT 507.500000 356.350000 508.500000 357.650000 ;
      RECT 416.500000 356.350000 499.500000 357.650000 ;
      RECT 407.500000 356.350000 408.500000 357.650000 ;
      RECT 366.500000 356.350000 399.500000 357.650000 ;
      RECT 357.500000 356.350000 358.500000 357.650000 ;
      RECT 316.500000 356.350000 349.500000 357.650000 ;
      RECT 307.500000 356.350000 308.500000 357.650000 ;
      RECT 266.500000 356.350000 299.500000 357.650000 ;
      RECT 257.500000 356.350000 258.500000 357.650000 ;
      RECT 216.500000 356.350000 249.500000 357.650000 ;
      RECT 207.500000 356.350000 208.500000 357.650000 ;
      RECT 166.500000 356.350000 199.500000 357.650000 ;
      RECT 157.500000 356.350000 158.500000 357.650000 ;
      RECT 116.500000 356.350000 149.500000 357.650000 ;
      RECT 107.500000 356.350000 108.500000 357.650000 ;
      RECT 29.500000 356.350000 99.500000 357.650000 ;
      RECT 15.500000 356.350000 16.500000 357.650000 ;
      RECT 0.000000 356.350000 2.500000 359.650000 ;
      RECT 1169.500000 355.650000 1186.000000 356.350000 ;
      RECT 1116.500000 355.650000 1156.500000 356.350000 ;
      RECT 1066.500000 355.650000 1108.500000 356.350000 ;
      RECT 1016.500000 355.650000 1058.500000 356.350000 ;
      RECT 966.500000 355.650000 1008.500000 356.350000 ;
      RECT 916.500000 355.650000 958.500000 356.350000 ;
      RECT 866.500000 355.650000 908.500000 356.350000 ;
      RECT 816.500000 355.650000 858.500000 356.350000 ;
      RECT 766.500000 355.650000 808.500000 356.350000 ;
      RECT 716.500000 355.650000 758.500000 356.350000 ;
      RECT 666.500000 355.650000 708.500000 356.350000 ;
      RECT 616.500000 355.650000 658.500000 356.350000 ;
      RECT 566.500000 355.650000 608.500000 356.350000 ;
      RECT 516.500000 355.650000 558.500000 356.350000 ;
      RECT 416.500000 355.650000 508.500000 356.350000 ;
      RECT 366.500000 355.650000 408.500000 356.350000 ;
      RECT 316.500000 355.650000 358.500000 356.350000 ;
      RECT 266.500000 355.650000 308.500000 356.350000 ;
      RECT 216.500000 355.650000 258.500000 356.350000 ;
      RECT 166.500000 355.650000 208.500000 356.350000 ;
      RECT 116.500000 355.650000 158.500000 356.350000 ;
      RECT 29.500000 355.650000 108.500000 356.350000 ;
      RECT 0.000000 355.650000 16.500000 356.350000 ;
      RECT 1169.500000 354.350000 1170.500000 355.650000 ;
      RECT 1116.500000 354.350000 1149.500000 355.650000 ;
      RECT 1107.500000 354.350000 1108.500000 355.650000 ;
      RECT 1066.500000 354.350000 1099.500000 355.650000 ;
      RECT 1057.500000 354.350000 1058.500000 355.650000 ;
      RECT 1016.500000 354.350000 1049.500000 355.650000 ;
      RECT 1007.500000 354.350000 1008.500000 355.650000 ;
      RECT 966.500000 354.350000 999.500000 355.650000 ;
      RECT 957.500000 354.350000 958.500000 355.650000 ;
      RECT 916.500000 354.350000 949.500000 355.650000 ;
      RECT 907.500000 354.350000 908.500000 355.650000 ;
      RECT 866.500000 354.350000 899.500000 355.650000 ;
      RECT 857.500000 354.350000 858.500000 355.650000 ;
      RECT 816.500000 354.350000 849.500000 355.650000 ;
      RECT 807.500000 354.350000 808.500000 355.650000 ;
      RECT 766.500000 354.350000 799.500000 355.650000 ;
      RECT 757.500000 354.350000 758.500000 355.650000 ;
      RECT 716.500000 354.350000 749.500000 355.650000 ;
      RECT 707.500000 354.350000 708.500000 355.650000 ;
      RECT 666.500000 354.350000 699.500000 355.650000 ;
      RECT 657.500000 354.350000 658.500000 355.650000 ;
      RECT 616.500000 354.350000 649.500000 355.650000 ;
      RECT 607.500000 354.350000 608.500000 355.650000 ;
      RECT 566.500000 354.350000 599.500000 355.650000 ;
      RECT 557.500000 354.350000 558.500000 355.650000 ;
      RECT 516.500000 354.350000 549.500000 355.650000 ;
      RECT 507.500000 354.350000 508.500000 355.650000 ;
      RECT 416.500000 354.350000 499.500000 355.650000 ;
      RECT 407.500000 354.350000 408.500000 355.650000 ;
      RECT 366.500000 354.350000 399.500000 355.650000 ;
      RECT 357.500000 354.350000 358.500000 355.650000 ;
      RECT 316.500000 354.350000 349.500000 355.650000 ;
      RECT 307.500000 354.350000 308.500000 355.650000 ;
      RECT 266.500000 354.350000 299.500000 355.650000 ;
      RECT 257.500000 354.350000 258.500000 355.650000 ;
      RECT 216.500000 354.350000 249.500000 355.650000 ;
      RECT 207.500000 354.350000 208.500000 355.650000 ;
      RECT 166.500000 354.350000 199.500000 355.650000 ;
      RECT 157.500000 354.350000 158.500000 355.650000 ;
      RECT 116.500000 354.350000 149.500000 355.650000 ;
      RECT 107.500000 354.350000 108.500000 355.650000 ;
      RECT 29.500000 354.350000 99.500000 355.650000 ;
      RECT 15.500000 354.350000 16.500000 355.650000 ;
      RECT 1157.500000 353.650000 1170.500000 354.350000 ;
      RECT 1107.500000 353.650000 1149.500000 354.350000 ;
      RECT 1057.500000 353.650000 1099.500000 354.350000 ;
      RECT 1007.500000 353.650000 1049.500000 354.350000 ;
      RECT 957.500000 353.650000 999.500000 354.350000 ;
      RECT 907.500000 353.650000 949.500000 354.350000 ;
      RECT 857.500000 353.650000 899.500000 354.350000 ;
      RECT 807.500000 353.650000 849.500000 354.350000 ;
      RECT 757.500000 353.650000 799.500000 354.350000 ;
      RECT 707.500000 353.650000 749.500000 354.350000 ;
      RECT 657.500000 353.650000 699.500000 354.350000 ;
      RECT 607.500000 353.650000 649.500000 354.350000 ;
      RECT 557.500000 353.650000 599.500000 354.350000 ;
      RECT 507.500000 353.650000 549.500000 354.350000 ;
      RECT 407.500000 353.650000 499.500000 354.350000 ;
      RECT 357.500000 353.650000 399.500000 354.350000 ;
      RECT 307.500000 353.650000 349.500000 354.350000 ;
      RECT 257.500000 353.650000 299.500000 354.350000 ;
      RECT 207.500000 353.650000 249.500000 354.350000 ;
      RECT 157.500000 353.650000 199.500000 354.350000 ;
      RECT 107.500000 353.650000 149.500000 354.350000 ;
      RECT 15.500000 353.650000 99.500000 354.350000 ;
      RECT 1183.500000 352.350000 1186.000000 355.650000 ;
      RECT 1169.500000 352.350000 1170.500000 353.650000 ;
      RECT 1116.500000 352.350000 1149.500000 353.650000 ;
      RECT 1107.500000 352.350000 1108.500000 353.650000 ;
      RECT 1066.500000 352.350000 1099.500000 353.650000 ;
      RECT 1057.500000 352.350000 1058.500000 353.650000 ;
      RECT 1016.500000 352.350000 1049.500000 353.650000 ;
      RECT 1007.500000 352.350000 1008.500000 353.650000 ;
      RECT 966.500000 352.350000 999.500000 353.650000 ;
      RECT 957.500000 352.350000 958.500000 353.650000 ;
      RECT 916.500000 352.350000 949.500000 353.650000 ;
      RECT 907.500000 352.350000 908.500000 353.650000 ;
      RECT 866.500000 352.350000 899.500000 353.650000 ;
      RECT 857.500000 352.350000 858.500000 353.650000 ;
      RECT 816.500000 352.350000 849.500000 353.650000 ;
      RECT 807.500000 352.350000 808.500000 353.650000 ;
      RECT 766.500000 352.350000 799.500000 353.650000 ;
      RECT 757.500000 352.350000 758.500000 353.650000 ;
      RECT 716.500000 352.350000 749.500000 353.650000 ;
      RECT 707.500000 352.350000 708.500000 353.650000 ;
      RECT 666.500000 352.350000 699.500000 353.650000 ;
      RECT 657.500000 352.350000 658.500000 353.650000 ;
      RECT 616.500000 352.350000 649.500000 353.650000 ;
      RECT 607.500000 352.350000 608.500000 353.650000 ;
      RECT 566.500000 352.350000 599.500000 353.650000 ;
      RECT 557.500000 352.350000 558.500000 353.650000 ;
      RECT 516.500000 352.350000 549.500000 353.650000 ;
      RECT 507.500000 352.350000 508.500000 353.650000 ;
      RECT 416.500000 352.350000 499.500000 353.650000 ;
      RECT 407.500000 352.350000 408.500000 353.650000 ;
      RECT 366.500000 352.350000 399.500000 353.650000 ;
      RECT 357.500000 352.350000 358.500000 353.650000 ;
      RECT 316.500000 352.350000 349.500000 353.650000 ;
      RECT 307.500000 352.350000 308.500000 353.650000 ;
      RECT 266.500000 352.350000 299.500000 353.650000 ;
      RECT 257.500000 352.350000 258.500000 353.650000 ;
      RECT 216.500000 352.350000 249.500000 353.650000 ;
      RECT 207.500000 352.350000 208.500000 353.650000 ;
      RECT 166.500000 352.350000 199.500000 353.650000 ;
      RECT 157.500000 352.350000 158.500000 353.650000 ;
      RECT 116.500000 352.350000 149.500000 353.650000 ;
      RECT 107.500000 352.350000 108.500000 353.650000 ;
      RECT 29.500000 352.350000 99.500000 353.650000 ;
      RECT 15.500000 352.350000 16.500000 353.650000 ;
      RECT 0.000000 352.350000 2.500000 355.650000 ;
      RECT 1169.500000 351.650000 1186.000000 352.350000 ;
      RECT 1116.500000 351.650000 1156.500000 352.350000 ;
      RECT 1066.500000 351.650000 1108.500000 352.350000 ;
      RECT 1016.500000 351.650000 1058.500000 352.350000 ;
      RECT 966.500000 351.650000 1008.500000 352.350000 ;
      RECT 916.500000 351.650000 958.500000 352.350000 ;
      RECT 866.500000 351.650000 908.500000 352.350000 ;
      RECT 816.500000 351.650000 858.500000 352.350000 ;
      RECT 766.500000 351.650000 808.500000 352.350000 ;
      RECT 716.500000 351.650000 758.500000 352.350000 ;
      RECT 666.500000 351.650000 708.500000 352.350000 ;
      RECT 616.500000 351.650000 658.500000 352.350000 ;
      RECT 566.500000 351.650000 608.500000 352.350000 ;
      RECT 516.500000 351.650000 558.500000 352.350000 ;
      RECT 416.500000 351.650000 508.500000 352.350000 ;
      RECT 366.500000 351.650000 408.500000 352.350000 ;
      RECT 316.500000 351.650000 358.500000 352.350000 ;
      RECT 266.500000 351.650000 308.500000 352.350000 ;
      RECT 216.500000 351.650000 258.500000 352.350000 ;
      RECT 166.500000 351.650000 208.500000 352.350000 ;
      RECT 116.500000 351.650000 158.500000 352.350000 ;
      RECT 29.500000 351.650000 108.500000 352.350000 ;
      RECT 0.000000 351.650000 16.500000 352.350000 ;
      RECT 1169.500000 350.350000 1170.500000 351.650000 ;
      RECT 1116.500000 350.350000 1149.500000 351.650000 ;
      RECT 1107.500000 350.350000 1108.500000 351.650000 ;
      RECT 1066.500000 350.350000 1099.500000 351.650000 ;
      RECT 1057.500000 350.350000 1058.500000 351.650000 ;
      RECT 1016.500000 350.350000 1049.500000 351.650000 ;
      RECT 1007.500000 350.350000 1008.500000 351.650000 ;
      RECT 966.500000 350.350000 999.500000 351.650000 ;
      RECT 957.500000 350.350000 958.500000 351.650000 ;
      RECT 916.500000 350.350000 949.500000 351.650000 ;
      RECT 907.500000 350.350000 908.500000 351.650000 ;
      RECT 866.500000 350.350000 899.500000 351.650000 ;
      RECT 857.500000 350.350000 858.500000 351.650000 ;
      RECT 816.500000 350.350000 849.500000 351.650000 ;
      RECT 807.500000 350.350000 808.500000 351.650000 ;
      RECT 766.500000 350.350000 799.500000 351.650000 ;
      RECT 757.500000 350.350000 758.500000 351.650000 ;
      RECT 716.500000 350.350000 749.500000 351.650000 ;
      RECT 707.500000 350.350000 708.500000 351.650000 ;
      RECT 666.500000 350.350000 699.500000 351.650000 ;
      RECT 657.500000 350.350000 658.500000 351.650000 ;
      RECT 616.500000 350.350000 649.500000 351.650000 ;
      RECT 607.500000 350.350000 608.500000 351.650000 ;
      RECT 566.500000 350.350000 599.500000 351.650000 ;
      RECT 557.500000 350.350000 558.500000 351.650000 ;
      RECT 516.500000 350.350000 549.500000 351.650000 ;
      RECT 507.500000 350.350000 508.500000 351.650000 ;
      RECT 416.500000 350.350000 499.500000 351.650000 ;
      RECT 407.500000 350.350000 408.500000 351.650000 ;
      RECT 366.500000 350.350000 399.500000 351.650000 ;
      RECT 357.500000 350.350000 358.500000 351.650000 ;
      RECT 316.500000 350.350000 349.500000 351.650000 ;
      RECT 307.500000 350.350000 308.500000 351.650000 ;
      RECT 266.500000 350.350000 299.500000 351.650000 ;
      RECT 257.500000 350.350000 258.500000 351.650000 ;
      RECT 216.500000 350.350000 249.500000 351.650000 ;
      RECT 207.500000 350.350000 208.500000 351.650000 ;
      RECT 166.500000 350.350000 199.500000 351.650000 ;
      RECT 157.500000 350.350000 158.500000 351.650000 ;
      RECT 116.500000 350.350000 149.500000 351.650000 ;
      RECT 107.500000 350.350000 108.500000 351.650000 ;
      RECT 29.500000 350.350000 99.500000 351.650000 ;
      RECT 15.500000 350.350000 16.500000 351.650000 ;
      RECT 1157.500000 349.650000 1170.500000 350.350000 ;
      RECT 1107.500000 349.650000 1149.500000 350.350000 ;
      RECT 1057.500000 349.650000 1099.500000 350.350000 ;
      RECT 1007.500000 349.650000 1049.500000 350.350000 ;
      RECT 957.500000 349.650000 999.500000 350.350000 ;
      RECT 907.500000 349.650000 949.500000 350.350000 ;
      RECT 857.500000 349.650000 899.500000 350.350000 ;
      RECT 807.500000 349.650000 849.500000 350.350000 ;
      RECT 757.500000 349.650000 799.500000 350.350000 ;
      RECT 707.500000 349.650000 749.500000 350.350000 ;
      RECT 657.500000 349.650000 699.500000 350.350000 ;
      RECT 607.500000 349.650000 649.500000 350.350000 ;
      RECT 557.500000 349.650000 599.500000 350.350000 ;
      RECT 507.500000 349.650000 549.500000 350.350000 ;
      RECT 407.500000 349.650000 499.500000 350.350000 ;
      RECT 357.500000 349.650000 399.500000 350.350000 ;
      RECT 307.500000 349.650000 349.500000 350.350000 ;
      RECT 257.500000 349.650000 299.500000 350.350000 ;
      RECT 207.500000 349.650000 249.500000 350.350000 ;
      RECT 157.500000 349.650000 199.500000 350.350000 ;
      RECT 107.500000 349.650000 149.500000 350.350000 ;
      RECT 15.500000 349.650000 99.500000 350.350000 ;
      RECT 1183.500000 348.350000 1186.000000 351.650000 ;
      RECT 1169.500000 348.350000 1170.500000 349.650000 ;
      RECT 1116.500000 348.350000 1149.500000 349.650000 ;
      RECT 1107.500000 348.350000 1108.500000 349.650000 ;
      RECT 1066.500000 348.350000 1099.500000 349.650000 ;
      RECT 1057.500000 348.350000 1058.500000 349.650000 ;
      RECT 1016.500000 348.350000 1049.500000 349.650000 ;
      RECT 1007.500000 348.350000 1008.500000 349.650000 ;
      RECT 966.500000 348.350000 999.500000 349.650000 ;
      RECT 957.500000 348.350000 958.500000 349.650000 ;
      RECT 916.500000 348.350000 949.500000 349.650000 ;
      RECT 907.500000 348.350000 908.500000 349.650000 ;
      RECT 866.500000 348.350000 899.500000 349.650000 ;
      RECT 857.500000 348.350000 858.500000 349.650000 ;
      RECT 816.500000 348.350000 849.500000 349.650000 ;
      RECT 807.500000 348.350000 808.500000 349.650000 ;
      RECT 766.500000 348.350000 799.500000 349.650000 ;
      RECT 757.500000 348.350000 758.500000 349.650000 ;
      RECT 716.500000 348.350000 749.500000 349.650000 ;
      RECT 707.500000 348.350000 708.500000 349.650000 ;
      RECT 666.500000 348.350000 699.500000 349.650000 ;
      RECT 657.500000 348.350000 658.500000 349.650000 ;
      RECT 616.500000 348.350000 649.500000 349.650000 ;
      RECT 607.500000 348.350000 608.500000 349.650000 ;
      RECT 566.500000 348.350000 599.500000 349.650000 ;
      RECT 557.500000 348.350000 558.500000 349.650000 ;
      RECT 516.500000 348.350000 549.500000 349.650000 ;
      RECT 507.500000 348.350000 508.500000 349.650000 ;
      RECT 466.500000 348.350000 499.500000 349.650000 ;
      RECT 407.500000 348.350000 408.500000 349.650000 ;
      RECT 366.500000 348.350000 399.500000 349.650000 ;
      RECT 357.500000 348.350000 358.500000 349.650000 ;
      RECT 316.500000 348.350000 349.500000 349.650000 ;
      RECT 307.500000 348.350000 308.500000 349.650000 ;
      RECT 266.500000 348.350000 299.500000 349.650000 ;
      RECT 257.500000 348.350000 258.500000 349.650000 ;
      RECT 216.500000 348.350000 249.500000 349.650000 ;
      RECT 207.500000 348.350000 208.500000 349.650000 ;
      RECT 166.500000 348.350000 199.500000 349.650000 ;
      RECT 157.500000 348.350000 158.500000 349.650000 ;
      RECT 116.500000 348.350000 149.500000 349.650000 ;
      RECT 107.500000 348.350000 108.500000 349.650000 ;
      RECT 66.500000 348.350000 99.500000 349.650000 ;
      RECT 15.500000 348.350000 16.500000 349.650000 ;
      RECT 0.000000 348.350000 2.500000 351.650000 ;
      RECT 1169.500000 347.650000 1186.000000 348.350000 ;
      RECT 1116.500000 347.650000 1156.500000 348.350000 ;
      RECT 1066.500000 347.650000 1108.500000 348.350000 ;
      RECT 1016.500000 347.650000 1058.500000 348.350000 ;
      RECT 966.500000 347.650000 1008.500000 348.350000 ;
      RECT 916.500000 347.650000 958.500000 348.350000 ;
      RECT 866.500000 347.650000 908.500000 348.350000 ;
      RECT 816.500000 347.650000 858.500000 348.350000 ;
      RECT 766.500000 347.650000 808.500000 348.350000 ;
      RECT 716.500000 347.650000 758.500000 348.350000 ;
      RECT 666.500000 347.650000 708.500000 348.350000 ;
      RECT 616.500000 347.650000 658.500000 348.350000 ;
      RECT 566.500000 347.650000 608.500000 348.350000 ;
      RECT 516.500000 347.650000 558.500000 348.350000 ;
      RECT 466.500000 347.650000 508.500000 348.350000 ;
      RECT 416.500000 347.650000 458.500000 349.650000 ;
      RECT 366.500000 347.650000 408.500000 348.350000 ;
      RECT 316.500000 347.650000 358.500000 348.350000 ;
      RECT 266.500000 347.650000 308.500000 348.350000 ;
      RECT 216.500000 347.650000 258.500000 348.350000 ;
      RECT 166.500000 347.650000 208.500000 348.350000 ;
      RECT 116.500000 347.650000 158.500000 348.350000 ;
      RECT 66.500000 347.650000 108.500000 348.350000 ;
      RECT 29.500000 347.650000 58.500000 349.650000 ;
      RECT 0.000000 347.650000 16.500000 348.350000 ;
      RECT 1169.500000 346.350000 1170.500000 347.650000 ;
      RECT 1116.500000 346.350000 1149.500000 347.650000 ;
      RECT 1107.500000 346.350000 1108.500000 347.650000 ;
      RECT 1066.500000 346.350000 1099.500000 347.650000 ;
      RECT 1057.500000 346.350000 1058.500000 347.650000 ;
      RECT 1016.500000 346.350000 1049.500000 347.650000 ;
      RECT 1007.500000 346.350000 1008.500000 347.650000 ;
      RECT 966.500000 346.350000 999.500000 347.650000 ;
      RECT 957.500000 346.350000 958.500000 347.650000 ;
      RECT 916.500000 346.350000 949.500000 347.650000 ;
      RECT 907.500000 346.350000 908.500000 347.650000 ;
      RECT 866.500000 346.350000 899.500000 347.650000 ;
      RECT 857.500000 346.350000 858.500000 347.650000 ;
      RECT 816.500000 346.350000 849.500000 347.650000 ;
      RECT 807.500000 346.350000 808.500000 347.650000 ;
      RECT 766.500000 346.350000 799.500000 347.650000 ;
      RECT 757.500000 346.350000 758.500000 347.650000 ;
      RECT 716.500000 346.350000 749.500000 347.650000 ;
      RECT 707.500000 346.350000 708.500000 347.650000 ;
      RECT 666.500000 346.350000 699.500000 347.650000 ;
      RECT 657.500000 346.350000 658.500000 347.650000 ;
      RECT 616.500000 346.350000 649.500000 347.650000 ;
      RECT 607.500000 346.350000 608.500000 347.650000 ;
      RECT 566.500000 346.350000 599.500000 347.650000 ;
      RECT 557.500000 346.350000 558.500000 347.650000 ;
      RECT 516.500000 346.350000 549.500000 347.650000 ;
      RECT 507.500000 346.350000 508.500000 347.650000 ;
      RECT 466.500000 346.350000 499.500000 347.650000 ;
      RECT 457.500000 346.350000 458.500000 347.650000 ;
      RECT 416.500000 346.350000 449.500000 347.650000 ;
      RECT 407.500000 346.350000 408.500000 347.650000 ;
      RECT 366.500000 346.350000 399.500000 347.650000 ;
      RECT 357.500000 346.350000 358.500000 347.650000 ;
      RECT 316.500000 346.350000 349.500000 347.650000 ;
      RECT 307.500000 346.350000 308.500000 347.650000 ;
      RECT 266.500000 346.350000 299.500000 347.650000 ;
      RECT 257.500000 346.350000 258.500000 347.650000 ;
      RECT 216.500000 346.350000 249.500000 347.650000 ;
      RECT 207.500000 346.350000 208.500000 347.650000 ;
      RECT 166.500000 346.350000 199.500000 347.650000 ;
      RECT 157.500000 346.350000 158.500000 347.650000 ;
      RECT 116.500000 346.350000 149.500000 347.650000 ;
      RECT 107.500000 346.350000 108.500000 347.650000 ;
      RECT 66.500000 346.350000 99.500000 347.650000 ;
      RECT 57.500000 346.350000 58.500000 347.650000 ;
      RECT 29.500000 346.350000 49.500000 347.650000 ;
      RECT 15.500000 346.350000 16.500000 347.650000 ;
      RECT 1157.500000 345.650000 1170.500000 346.350000 ;
      RECT 1107.500000 345.650000 1149.500000 346.350000 ;
      RECT 1057.500000 345.650000 1099.500000 346.350000 ;
      RECT 1007.500000 345.650000 1049.500000 346.350000 ;
      RECT 957.500000 345.650000 999.500000 346.350000 ;
      RECT 907.500000 345.650000 949.500000 346.350000 ;
      RECT 857.500000 345.650000 899.500000 346.350000 ;
      RECT 807.500000 345.650000 849.500000 346.350000 ;
      RECT 757.500000 345.650000 799.500000 346.350000 ;
      RECT 707.500000 345.650000 749.500000 346.350000 ;
      RECT 657.500000 345.650000 699.500000 346.350000 ;
      RECT 607.500000 345.650000 649.500000 346.350000 ;
      RECT 557.500000 345.650000 599.500000 346.350000 ;
      RECT 507.500000 345.650000 549.500000 346.350000 ;
      RECT 457.500000 345.650000 499.500000 346.350000 ;
      RECT 407.500000 345.650000 449.500000 346.350000 ;
      RECT 357.500000 345.650000 399.500000 346.350000 ;
      RECT 307.500000 345.650000 349.500000 346.350000 ;
      RECT 257.500000 345.650000 299.500000 346.350000 ;
      RECT 207.500000 345.650000 249.500000 346.350000 ;
      RECT 157.500000 345.650000 199.500000 346.350000 ;
      RECT 107.500000 345.650000 149.500000 346.350000 ;
      RECT 57.500000 345.650000 99.500000 346.350000 ;
      RECT 15.500000 345.650000 49.500000 346.350000 ;
      RECT 1183.500000 344.350000 1186.000000 347.650000 ;
      RECT 1169.500000 344.350000 1170.500000 345.650000 ;
      RECT 1116.500000 344.350000 1149.500000 345.650000 ;
      RECT 1107.500000 344.350000 1108.500000 345.650000 ;
      RECT 1066.500000 344.350000 1099.500000 345.650000 ;
      RECT 1057.500000 344.350000 1058.500000 345.650000 ;
      RECT 1016.500000 344.350000 1049.500000 345.650000 ;
      RECT 1007.500000 344.350000 1008.500000 345.650000 ;
      RECT 966.500000 344.350000 999.500000 345.650000 ;
      RECT 957.500000 344.350000 958.500000 345.650000 ;
      RECT 916.500000 344.350000 949.500000 345.650000 ;
      RECT 907.500000 344.350000 908.500000 345.650000 ;
      RECT 866.500000 344.350000 899.500000 345.650000 ;
      RECT 857.500000 344.350000 858.500000 345.650000 ;
      RECT 816.500000 344.350000 849.500000 345.650000 ;
      RECT 807.500000 344.350000 808.500000 345.650000 ;
      RECT 766.500000 344.350000 799.500000 345.650000 ;
      RECT 757.500000 344.350000 758.500000 345.650000 ;
      RECT 716.500000 344.350000 749.500000 345.650000 ;
      RECT 707.500000 344.350000 708.500000 345.650000 ;
      RECT 666.500000 344.350000 699.500000 345.650000 ;
      RECT 657.500000 344.350000 658.500000 345.650000 ;
      RECT 616.500000 344.350000 649.500000 345.650000 ;
      RECT 607.500000 344.350000 608.500000 345.650000 ;
      RECT 566.500000 344.350000 599.500000 345.650000 ;
      RECT 557.500000 344.350000 558.500000 345.650000 ;
      RECT 516.500000 344.350000 549.500000 345.650000 ;
      RECT 507.500000 344.350000 508.500000 345.650000 ;
      RECT 466.500000 344.350000 499.500000 345.650000 ;
      RECT 457.500000 344.350000 458.500000 345.650000 ;
      RECT 416.500000 344.350000 449.500000 345.650000 ;
      RECT 407.500000 344.350000 408.500000 345.650000 ;
      RECT 366.500000 344.350000 399.500000 345.650000 ;
      RECT 357.500000 344.350000 358.500000 345.650000 ;
      RECT 316.500000 344.350000 349.500000 345.650000 ;
      RECT 307.500000 344.350000 308.500000 345.650000 ;
      RECT 266.500000 344.350000 299.500000 345.650000 ;
      RECT 257.500000 344.350000 258.500000 345.650000 ;
      RECT 216.500000 344.350000 249.500000 345.650000 ;
      RECT 207.500000 344.350000 208.500000 345.650000 ;
      RECT 166.500000 344.350000 199.500000 345.650000 ;
      RECT 157.500000 344.350000 158.500000 345.650000 ;
      RECT 116.500000 344.350000 149.500000 345.650000 ;
      RECT 107.500000 344.350000 108.500000 345.650000 ;
      RECT 66.500000 344.350000 99.500000 345.650000 ;
      RECT 57.500000 344.350000 58.500000 345.650000 ;
      RECT 29.500000 344.350000 49.500000 345.650000 ;
      RECT 15.500000 344.350000 16.500000 345.650000 ;
      RECT 0.000000 344.350000 2.500000 347.650000 ;
      RECT 1169.500000 343.650000 1186.000000 344.350000 ;
      RECT 1116.500000 343.650000 1156.500000 344.350000 ;
      RECT 1066.500000 343.650000 1108.500000 344.350000 ;
      RECT 1016.500000 343.650000 1058.500000 344.350000 ;
      RECT 966.500000 343.650000 1008.500000 344.350000 ;
      RECT 916.500000 343.650000 958.500000 344.350000 ;
      RECT 866.500000 343.650000 908.500000 344.350000 ;
      RECT 816.500000 343.650000 858.500000 344.350000 ;
      RECT 766.500000 343.650000 808.500000 344.350000 ;
      RECT 716.500000 343.650000 758.500000 344.350000 ;
      RECT 666.500000 343.650000 708.500000 344.350000 ;
      RECT 616.500000 343.650000 658.500000 344.350000 ;
      RECT 566.500000 343.650000 608.500000 344.350000 ;
      RECT 516.500000 343.650000 558.500000 344.350000 ;
      RECT 466.500000 343.650000 508.500000 344.350000 ;
      RECT 416.500000 343.650000 458.500000 344.350000 ;
      RECT 366.500000 343.650000 408.500000 344.350000 ;
      RECT 316.500000 343.650000 358.500000 344.350000 ;
      RECT 266.500000 343.650000 308.500000 344.350000 ;
      RECT 216.500000 343.650000 258.500000 344.350000 ;
      RECT 166.500000 343.650000 208.500000 344.350000 ;
      RECT 116.500000 343.650000 158.500000 344.350000 ;
      RECT 66.500000 343.650000 108.500000 344.350000 ;
      RECT 29.500000 343.650000 58.500000 344.350000 ;
      RECT 0.000000 343.650000 16.500000 344.350000 ;
      RECT 1169.500000 342.350000 1170.500000 343.650000 ;
      RECT 1116.500000 342.350000 1149.500000 343.650000 ;
      RECT 1107.500000 342.350000 1108.500000 343.650000 ;
      RECT 1066.500000 342.350000 1099.500000 343.650000 ;
      RECT 1057.500000 342.350000 1058.500000 343.650000 ;
      RECT 1016.500000 342.350000 1049.500000 343.650000 ;
      RECT 1007.500000 342.350000 1008.500000 343.650000 ;
      RECT 966.500000 342.350000 999.500000 343.650000 ;
      RECT 957.500000 342.350000 958.500000 343.650000 ;
      RECT 916.500000 342.350000 949.500000 343.650000 ;
      RECT 907.500000 342.350000 908.500000 343.650000 ;
      RECT 866.500000 342.350000 899.500000 343.650000 ;
      RECT 857.500000 342.350000 858.500000 343.650000 ;
      RECT 816.500000 342.350000 849.500000 343.650000 ;
      RECT 807.500000 342.350000 808.500000 343.650000 ;
      RECT 766.500000 342.350000 799.500000 343.650000 ;
      RECT 757.500000 342.350000 758.500000 343.650000 ;
      RECT 716.500000 342.350000 749.500000 343.650000 ;
      RECT 707.500000 342.350000 708.500000 343.650000 ;
      RECT 666.500000 342.350000 699.500000 343.650000 ;
      RECT 657.500000 342.350000 658.500000 343.650000 ;
      RECT 616.500000 342.350000 649.500000 343.650000 ;
      RECT 607.500000 342.350000 608.500000 343.650000 ;
      RECT 566.500000 342.350000 599.500000 343.650000 ;
      RECT 557.500000 342.350000 558.500000 343.650000 ;
      RECT 516.500000 342.350000 549.500000 343.650000 ;
      RECT 507.500000 342.350000 508.500000 343.650000 ;
      RECT 466.500000 342.350000 499.500000 343.650000 ;
      RECT 457.500000 342.350000 458.500000 343.650000 ;
      RECT 416.500000 342.350000 449.500000 343.650000 ;
      RECT 407.500000 342.350000 408.500000 343.650000 ;
      RECT 366.500000 342.350000 399.500000 343.650000 ;
      RECT 357.500000 342.350000 358.500000 343.650000 ;
      RECT 316.500000 342.350000 349.500000 343.650000 ;
      RECT 307.500000 342.350000 308.500000 343.650000 ;
      RECT 266.500000 342.350000 299.500000 343.650000 ;
      RECT 257.500000 342.350000 258.500000 343.650000 ;
      RECT 216.500000 342.350000 249.500000 343.650000 ;
      RECT 207.500000 342.350000 208.500000 343.650000 ;
      RECT 166.500000 342.350000 199.500000 343.650000 ;
      RECT 157.500000 342.350000 158.500000 343.650000 ;
      RECT 116.500000 342.350000 149.500000 343.650000 ;
      RECT 107.500000 342.350000 108.500000 343.650000 ;
      RECT 66.500000 342.350000 99.500000 343.650000 ;
      RECT 57.500000 342.350000 58.500000 343.650000 ;
      RECT 29.500000 342.350000 49.500000 343.650000 ;
      RECT 15.500000 342.350000 16.500000 343.650000 ;
      RECT 1157.500000 341.650000 1170.500000 342.350000 ;
      RECT 1107.500000 341.650000 1149.500000 342.350000 ;
      RECT 1057.500000 341.650000 1099.500000 342.350000 ;
      RECT 1007.500000 341.650000 1049.500000 342.350000 ;
      RECT 957.500000 341.650000 999.500000 342.350000 ;
      RECT 907.500000 341.650000 949.500000 342.350000 ;
      RECT 857.500000 341.650000 899.500000 342.350000 ;
      RECT 807.500000 341.650000 849.500000 342.350000 ;
      RECT 757.500000 341.650000 799.500000 342.350000 ;
      RECT 707.500000 341.650000 749.500000 342.350000 ;
      RECT 657.500000 341.650000 699.500000 342.350000 ;
      RECT 607.500000 341.650000 649.500000 342.350000 ;
      RECT 557.500000 341.650000 599.500000 342.350000 ;
      RECT 507.500000 341.650000 549.500000 342.350000 ;
      RECT 457.500000 341.650000 499.500000 342.350000 ;
      RECT 407.500000 341.650000 449.500000 342.350000 ;
      RECT 357.500000 341.650000 399.500000 342.350000 ;
      RECT 307.500000 341.650000 349.500000 342.350000 ;
      RECT 257.500000 341.650000 299.500000 342.350000 ;
      RECT 207.500000 341.650000 249.500000 342.350000 ;
      RECT 157.500000 341.650000 199.500000 342.350000 ;
      RECT 107.500000 341.650000 149.500000 342.350000 ;
      RECT 57.500000 341.650000 99.500000 342.350000 ;
      RECT 15.500000 341.650000 49.500000 342.350000 ;
      RECT 1183.500000 340.350000 1186.000000 343.650000 ;
      RECT 1169.500000 340.350000 1170.500000 341.650000 ;
      RECT 1116.500000 340.350000 1149.500000 341.650000 ;
      RECT 1107.500000 340.350000 1108.500000 341.650000 ;
      RECT 1066.500000 340.350000 1099.500000 341.650000 ;
      RECT 1057.500000 340.350000 1058.500000 341.650000 ;
      RECT 1016.500000 340.350000 1049.500000 341.650000 ;
      RECT 1007.500000 340.350000 1008.500000 341.650000 ;
      RECT 966.500000 340.350000 999.500000 341.650000 ;
      RECT 957.500000 340.350000 958.500000 341.650000 ;
      RECT 916.500000 340.350000 949.500000 341.650000 ;
      RECT 907.500000 340.350000 908.500000 341.650000 ;
      RECT 866.500000 340.350000 899.500000 341.650000 ;
      RECT 857.500000 340.350000 858.500000 341.650000 ;
      RECT 816.500000 340.350000 849.500000 341.650000 ;
      RECT 807.500000 340.350000 808.500000 341.650000 ;
      RECT 766.500000 340.350000 799.500000 341.650000 ;
      RECT 757.500000 340.350000 758.500000 341.650000 ;
      RECT 716.500000 340.350000 749.500000 341.650000 ;
      RECT 707.500000 340.350000 708.500000 341.650000 ;
      RECT 666.500000 340.350000 699.500000 341.650000 ;
      RECT 657.500000 340.350000 658.500000 341.650000 ;
      RECT 616.500000 340.350000 649.500000 341.650000 ;
      RECT 607.500000 340.350000 608.500000 341.650000 ;
      RECT 566.500000 340.350000 599.500000 341.650000 ;
      RECT 557.500000 340.350000 558.500000 341.650000 ;
      RECT 516.500000 340.350000 549.500000 341.650000 ;
      RECT 507.500000 340.350000 508.500000 341.650000 ;
      RECT 466.500000 340.350000 499.500000 341.650000 ;
      RECT 457.500000 340.350000 458.500000 341.650000 ;
      RECT 416.500000 340.350000 449.500000 341.650000 ;
      RECT 407.500000 340.350000 408.500000 341.650000 ;
      RECT 366.500000 340.350000 399.500000 341.650000 ;
      RECT 357.500000 340.350000 358.500000 341.650000 ;
      RECT 316.500000 340.350000 349.500000 341.650000 ;
      RECT 307.500000 340.350000 308.500000 341.650000 ;
      RECT 266.500000 340.350000 299.500000 341.650000 ;
      RECT 257.500000 340.350000 258.500000 341.650000 ;
      RECT 216.500000 340.350000 249.500000 341.650000 ;
      RECT 207.500000 340.350000 208.500000 341.650000 ;
      RECT 166.500000 340.350000 199.500000 341.650000 ;
      RECT 157.500000 340.350000 158.500000 341.650000 ;
      RECT 116.500000 340.350000 149.500000 341.650000 ;
      RECT 107.500000 340.350000 108.500000 341.650000 ;
      RECT 66.500000 340.350000 99.500000 341.650000 ;
      RECT 57.500000 340.350000 58.500000 341.650000 ;
      RECT 29.500000 340.350000 49.500000 341.650000 ;
      RECT 15.500000 340.350000 16.500000 341.650000 ;
      RECT 0.000000 340.350000 2.500000 343.650000 ;
      RECT 1169.500000 339.650000 1186.000000 340.350000 ;
      RECT 1116.500000 339.650000 1156.500000 340.350000 ;
      RECT 1066.500000 339.650000 1108.500000 340.350000 ;
      RECT 1016.500000 339.650000 1058.500000 340.350000 ;
      RECT 966.500000 339.650000 1008.500000 340.350000 ;
      RECT 916.500000 339.650000 958.500000 340.350000 ;
      RECT 866.500000 339.650000 908.500000 340.350000 ;
      RECT 816.500000 339.650000 858.500000 340.350000 ;
      RECT 766.500000 339.650000 808.500000 340.350000 ;
      RECT 716.500000 339.650000 758.500000 340.350000 ;
      RECT 666.500000 339.650000 708.500000 340.350000 ;
      RECT 616.500000 339.650000 658.500000 340.350000 ;
      RECT 566.500000 339.650000 608.500000 340.350000 ;
      RECT 516.500000 339.650000 558.500000 340.350000 ;
      RECT 466.500000 339.650000 508.500000 340.350000 ;
      RECT 416.500000 339.650000 458.500000 340.350000 ;
      RECT 366.500000 339.650000 408.500000 340.350000 ;
      RECT 316.500000 339.650000 358.500000 340.350000 ;
      RECT 266.500000 339.650000 308.500000 340.350000 ;
      RECT 216.500000 339.650000 258.500000 340.350000 ;
      RECT 166.500000 339.650000 208.500000 340.350000 ;
      RECT 116.500000 339.650000 158.500000 340.350000 ;
      RECT 66.500000 339.650000 108.500000 340.350000 ;
      RECT 29.500000 339.650000 58.500000 340.350000 ;
      RECT 0.000000 339.650000 16.500000 340.350000 ;
      RECT 1169.500000 338.350000 1170.500000 339.650000 ;
      RECT 1116.500000 338.350000 1149.500000 339.650000 ;
      RECT 1107.500000 338.350000 1108.500000 339.650000 ;
      RECT 1066.500000 338.350000 1099.500000 339.650000 ;
      RECT 1057.500000 338.350000 1058.500000 339.650000 ;
      RECT 1016.500000 338.350000 1049.500000 339.650000 ;
      RECT 1007.500000 338.350000 1008.500000 339.650000 ;
      RECT 966.500000 338.350000 999.500000 339.650000 ;
      RECT 957.500000 338.350000 958.500000 339.650000 ;
      RECT 916.500000 338.350000 949.500000 339.650000 ;
      RECT 907.500000 338.350000 908.500000 339.650000 ;
      RECT 866.500000 338.350000 899.500000 339.650000 ;
      RECT 857.500000 338.350000 858.500000 339.650000 ;
      RECT 816.500000 338.350000 849.500000 339.650000 ;
      RECT 807.500000 338.350000 808.500000 339.650000 ;
      RECT 766.500000 338.350000 799.500000 339.650000 ;
      RECT 757.500000 338.350000 758.500000 339.650000 ;
      RECT 716.500000 338.350000 749.500000 339.650000 ;
      RECT 707.500000 338.350000 708.500000 339.650000 ;
      RECT 666.500000 338.350000 699.500000 339.650000 ;
      RECT 657.500000 338.350000 658.500000 339.650000 ;
      RECT 616.500000 338.350000 649.500000 339.650000 ;
      RECT 607.500000 338.350000 608.500000 339.650000 ;
      RECT 566.500000 338.350000 599.500000 339.650000 ;
      RECT 557.500000 338.350000 558.500000 339.650000 ;
      RECT 516.500000 338.350000 549.500000 339.650000 ;
      RECT 507.500000 338.350000 508.500000 339.650000 ;
      RECT 466.500000 338.350000 499.500000 339.650000 ;
      RECT 457.500000 338.350000 458.500000 339.650000 ;
      RECT 416.500000 338.350000 449.500000 339.650000 ;
      RECT 407.500000 338.350000 408.500000 339.650000 ;
      RECT 366.500000 338.350000 399.500000 339.650000 ;
      RECT 357.500000 338.350000 358.500000 339.650000 ;
      RECT 316.500000 338.350000 349.500000 339.650000 ;
      RECT 307.500000 338.350000 308.500000 339.650000 ;
      RECT 266.500000 338.350000 299.500000 339.650000 ;
      RECT 257.500000 338.350000 258.500000 339.650000 ;
      RECT 216.500000 338.350000 249.500000 339.650000 ;
      RECT 207.500000 338.350000 208.500000 339.650000 ;
      RECT 166.500000 338.350000 199.500000 339.650000 ;
      RECT 157.500000 338.350000 158.500000 339.650000 ;
      RECT 116.500000 338.350000 149.500000 339.650000 ;
      RECT 107.500000 338.350000 108.500000 339.650000 ;
      RECT 66.500000 338.350000 99.500000 339.650000 ;
      RECT 57.500000 338.350000 58.500000 339.650000 ;
      RECT 29.500000 338.350000 49.500000 339.650000 ;
      RECT 15.500000 338.350000 16.500000 339.650000 ;
      RECT 1157.500000 337.650000 1170.500000 338.350000 ;
      RECT 1107.500000 337.650000 1149.500000 338.350000 ;
      RECT 1057.500000 337.650000 1099.500000 338.350000 ;
      RECT 1007.500000 337.650000 1049.500000 338.350000 ;
      RECT 957.500000 337.650000 999.500000 338.350000 ;
      RECT 907.500000 337.650000 949.500000 338.350000 ;
      RECT 857.500000 337.650000 899.500000 338.350000 ;
      RECT 807.500000 337.650000 849.500000 338.350000 ;
      RECT 757.500000 337.650000 799.500000 338.350000 ;
      RECT 707.500000 337.650000 749.500000 338.350000 ;
      RECT 657.500000 337.650000 699.500000 338.350000 ;
      RECT 607.500000 337.650000 649.500000 338.350000 ;
      RECT 557.500000 337.650000 599.500000 338.350000 ;
      RECT 507.500000 337.650000 549.500000 338.350000 ;
      RECT 457.500000 337.650000 499.500000 338.350000 ;
      RECT 407.500000 337.650000 449.500000 338.350000 ;
      RECT 357.500000 337.650000 399.500000 338.350000 ;
      RECT 307.500000 337.650000 349.500000 338.350000 ;
      RECT 257.500000 337.650000 299.500000 338.350000 ;
      RECT 207.500000 337.650000 249.500000 338.350000 ;
      RECT 157.500000 337.650000 199.500000 338.350000 ;
      RECT 107.500000 337.650000 149.500000 338.350000 ;
      RECT 57.500000 337.650000 99.500000 338.350000 ;
      RECT 15.500000 337.650000 49.500000 338.350000 ;
      RECT 1183.500000 336.350000 1186.000000 339.650000 ;
      RECT 1169.500000 336.350000 1170.500000 337.650000 ;
      RECT 1116.500000 336.350000 1149.500000 337.650000 ;
      RECT 1107.500000 336.350000 1108.500000 337.650000 ;
      RECT 1066.500000 336.350000 1099.500000 337.650000 ;
      RECT 1057.500000 336.350000 1058.500000 337.650000 ;
      RECT 1016.500000 336.350000 1049.500000 337.650000 ;
      RECT 1007.500000 336.350000 1008.500000 337.650000 ;
      RECT 966.500000 336.350000 999.500000 337.650000 ;
      RECT 957.500000 336.350000 958.500000 337.650000 ;
      RECT 916.500000 336.350000 949.500000 337.650000 ;
      RECT 907.500000 336.350000 908.500000 337.650000 ;
      RECT 866.500000 336.350000 899.500000 337.650000 ;
      RECT 857.500000 336.350000 858.500000 337.650000 ;
      RECT 816.500000 336.350000 849.500000 337.650000 ;
      RECT 807.500000 336.350000 808.500000 337.650000 ;
      RECT 766.500000 336.350000 799.500000 337.650000 ;
      RECT 757.500000 336.350000 758.500000 337.650000 ;
      RECT 716.500000 336.350000 749.500000 337.650000 ;
      RECT 707.500000 336.350000 708.500000 337.650000 ;
      RECT 666.500000 336.350000 699.500000 337.650000 ;
      RECT 657.500000 336.350000 658.500000 337.650000 ;
      RECT 616.500000 336.350000 649.500000 337.650000 ;
      RECT 607.500000 336.350000 608.500000 337.650000 ;
      RECT 566.500000 336.350000 599.500000 337.650000 ;
      RECT 557.500000 336.350000 558.500000 337.650000 ;
      RECT 516.500000 336.350000 549.500000 337.650000 ;
      RECT 507.500000 336.350000 508.500000 337.650000 ;
      RECT 466.500000 336.350000 499.500000 337.650000 ;
      RECT 457.500000 336.350000 458.500000 337.650000 ;
      RECT 416.500000 336.350000 449.500000 337.650000 ;
      RECT 407.500000 336.350000 408.500000 337.650000 ;
      RECT 366.500000 336.350000 399.500000 337.650000 ;
      RECT 357.500000 336.350000 358.500000 337.650000 ;
      RECT 316.500000 336.350000 349.500000 337.650000 ;
      RECT 307.500000 336.350000 308.500000 337.650000 ;
      RECT 266.500000 336.350000 299.500000 337.650000 ;
      RECT 257.500000 336.350000 258.500000 337.650000 ;
      RECT 216.500000 336.350000 249.500000 337.650000 ;
      RECT 207.500000 336.350000 208.500000 337.650000 ;
      RECT 166.500000 336.350000 199.500000 337.650000 ;
      RECT 157.500000 336.350000 158.500000 337.650000 ;
      RECT 116.500000 336.350000 149.500000 337.650000 ;
      RECT 107.500000 336.350000 108.500000 337.650000 ;
      RECT 66.500000 336.350000 99.500000 337.650000 ;
      RECT 57.500000 336.350000 58.500000 337.650000 ;
      RECT 29.500000 336.350000 49.500000 337.650000 ;
      RECT 15.500000 336.350000 16.500000 337.650000 ;
      RECT 0.000000 336.350000 2.500000 339.650000 ;
      RECT 1169.500000 335.650000 1186.000000 336.350000 ;
      RECT 1116.500000 335.650000 1156.500000 336.350000 ;
      RECT 1066.500000 335.650000 1108.500000 336.350000 ;
      RECT 1016.500000 335.650000 1058.500000 336.350000 ;
      RECT 966.500000 335.650000 1008.500000 336.350000 ;
      RECT 916.500000 335.650000 958.500000 336.350000 ;
      RECT 866.500000 335.650000 908.500000 336.350000 ;
      RECT 816.500000 335.650000 858.500000 336.350000 ;
      RECT 766.500000 335.650000 808.500000 336.350000 ;
      RECT 716.500000 335.650000 758.500000 336.350000 ;
      RECT 666.500000 335.650000 708.500000 336.350000 ;
      RECT 616.500000 335.650000 658.500000 336.350000 ;
      RECT 566.500000 335.650000 608.500000 336.350000 ;
      RECT 516.500000 335.650000 558.500000 336.350000 ;
      RECT 466.500000 335.650000 508.500000 336.350000 ;
      RECT 416.500000 335.650000 458.500000 336.350000 ;
      RECT 366.500000 335.650000 408.500000 336.350000 ;
      RECT 316.500000 335.650000 358.500000 336.350000 ;
      RECT 266.500000 335.650000 308.500000 336.350000 ;
      RECT 216.500000 335.650000 258.500000 336.350000 ;
      RECT 166.500000 335.650000 208.500000 336.350000 ;
      RECT 116.500000 335.650000 158.500000 336.350000 ;
      RECT 66.500000 335.650000 108.500000 336.350000 ;
      RECT 29.500000 335.650000 58.500000 336.350000 ;
      RECT 0.000000 335.650000 16.500000 336.350000 ;
      RECT 1169.500000 334.350000 1170.500000 335.650000 ;
      RECT 1116.500000 334.350000 1149.500000 335.650000 ;
      RECT 1107.500000 334.350000 1108.500000 335.650000 ;
      RECT 1066.500000 334.350000 1099.500000 335.650000 ;
      RECT 1057.500000 334.350000 1058.500000 335.650000 ;
      RECT 1016.500000 334.350000 1049.500000 335.650000 ;
      RECT 1007.500000 334.350000 1008.500000 335.650000 ;
      RECT 966.500000 334.350000 999.500000 335.650000 ;
      RECT 957.500000 334.350000 958.500000 335.650000 ;
      RECT 916.500000 334.350000 949.500000 335.650000 ;
      RECT 907.500000 334.350000 908.500000 335.650000 ;
      RECT 866.500000 334.350000 899.500000 335.650000 ;
      RECT 857.500000 334.350000 858.500000 335.650000 ;
      RECT 816.500000 334.350000 849.500000 335.650000 ;
      RECT 807.500000 334.350000 808.500000 335.650000 ;
      RECT 766.500000 334.350000 799.500000 335.650000 ;
      RECT 757.500000 334.350000 758.500000 335.650000 ;
      RECT 716.500000 334.350000 749.500000 335.650000 ;
      RECT 707.500000 334.350000 708.500000 335.650000 ;
      RECT 666.500000 334.350000 699.500000 335.650000 ;
      RECT 657.500000 334.350000 658.500000 335.650000 ;
      RECT 616.500000 334.350000 649.500000 335.650000 ;
      RECT 607.500000 334.350000 608.500000 335.650000 ;
      RECT 566.500000 334.350000 599.500000 335.650000 ;
      RECT 557.500000 334.350000 558.500000 335.650000 ;
      RECT 516.500000 334.350000 549.500000 335.650000 ;
      RECT 507.500000 334.350000 508.500000 335.650000 ;
      RECT 466.500000 334.350000 499.500000 335.650000 ;
      RECT 457.500000 334.350000 458.500000 335.650000 ;
      RECT 416.500000 334.350000 449.500000 335.650000 ;
      RECT 407.500000 334.350000 408.500000 335.650000 ;
      RECT 366.500000 334.350000 399.500000 335.650000 ;
      RECT 357.500000 334.350000 358.500000 335.650000 ;
      RECT 316.500000 334.350000 349.500000 335.650000 ;
      RECT 307.500000 334.350000 308.500000 335.650000 ;
      RECT 266.500000 334.350000 299.500000 335.650000 ;
      RECT 257.500000 334.350000 258.500000 335.650000 ;
      RECT 216.500000 334.350000 249.500000 335.650000 ;
      RECT 207.500000 334.350000 208.500000 335.650000 ;
      RECT 166.500000 334.350000 199.500000 335.650000 ;
      RECT 157.500000 334.350000 158.500000 335.650000 ;
      RECT 116.500000 334.350000 149.500000 335.650000 ;
      RECT 107.500000 334.350000 108.500000 335.650000 ;
      RECT 66.500000 334.350000 99.500000 335.650000 ;
      RECT 57.500000 334.350000 58.500000 335.650000 ;
      RECT 29.500000 334.350000 49.500000 335.650000 ;
      RECT 15.500000 334.350000 16.500000 335.650000 ;
      RECT 1157.500000 333.650000 1170.500000 334.350000 ;
      RECT 1107.500000 333.650000 1149.500000 334.350000 ;
      RECT 1057.500000 333.650000 1099.500000 334.350000 ;
      RECT 1007.500000 333.650000 1049.500000 334.350000 ;
      RECT 957.500000 333.650000 999.500000 334.350000 ;
      RECT 907.500000 333.650000 949.500000 334.350000 ;
      RECT 857.500000 333.650000 899.500000 334.350000 ;
      RECT 807.500000 333.650000 849.500000 334.350000 ;
      RECT 757.500000 333.650000 799.500000 334.350000 ;
      RECT 707.500000 333.650000 749.500000 334.350000 ;
      RECT 657.500000 333.650000 699.500000 334.350000 ;
      RECT 607.500000 333.650000 649.500000 334.350000 ;
      RECT 557.500000 333.650000 599.500000 334.350000 ;
      RECT 507.500000 333.650000 549.500000 334.350000 ;
      RECT 457.500000 333.650000 499.500000 334.350000 ;
      RECT 407.500000 333.650000 449.500000 334.350000 ;
      RECT 357.500000 333.650000 399.500000 334.350000 ;
      RECT 307.500000 333.650000 349.500000 334.350000 ;
      RECT 257.500000 333.650000 299.500000 334.350000 ;
      RECT 207.500000 333.650000 249.500000 334.350000 ;
      RECT 157.500000 333.650000 199.500000 334.350000 ;
      RECT 107.500000 333.650000 149.500000 334.350000 ;
      RECT 57.500000 333.650000 99.500000 334.350000 ;
      RECT 15.500000 333.650000 49.500000 334.350000 ;
      RECT 1183.500000 332.350000 1186.000000 335.650000 ;
      RECT 1169.500000 332.350000 1170.500000 333.650000 ;
      RECT 1116.500000 332.350000 1149.500000 333.650000 ;
      RECT 1107.500000 332.350000 1108.500000 333.650000 ;
      RECT 1066.500000 332.350000 1099.500000 333.650000 ;
      RECT 1057.500000 332.350000 1058.500000 333.650000 ;
      RECT 1016.500000 332.350000 1049.500000 333.650000 ;
      RECT 1007.500000 332.350000 1008.500000 333.650000 ;
      RECT 966.500000 332.350000 999.500000 333.650000 ;
      RECT 957.500000 332.350000 958.500000 333.650000 ;
      RECT 916.500000 332.350000 949.500000 333.650000 ;
      RECT 907.500000 332.350000 908.500000 333.650000 ;
      RECT 866.500000 332.350000 899.500000 333.650000 ;
      RECT 857.500000 332.350000 858.500000 333.650000 ;
      RECT 816.500000 332.350000 849.500000 333.650000 ;
      RECT 807.500000 332.350000 808.500000 333.650000 ;
      RECT 766.500000 332.350000 799.500000 333.650000 ;
      RECT 757.500000 332.350000 758.500000 333.650000 ;
      RECT 716.500000 332.350000 749.500000 333.650000 ;
      RECT 707.500000 332.350000 708.500000 333.650000 ;
      RECT 666.500000 332.350000 699.500000 333.650000 ;
      RECT 657.500000 332.350000 658.500000 333.650000 ;
      RECT 616.500000 332.350000 649.500000 333.650000 ;
      RECT 607.500000 332.350000 608.500000 333.650000 ;
      RECT 566.500000 332.350000 599.500000 333.650000 ;
      RECT 557.500000 332.350000 558.500000 333.650000 ;
      RECT 516.500000 332.350000 549.500000 333.650000 ;
      RECT 507.500000 332.350000 508.500000 333.650000 ;
      RECT 466.500000 332.350000 499.500000 333.650000 ;
      RECT 457.500000 332.350000 458.500000 333.650000 ;
      RECT 416.500000 332.350000 449.500000 333.650000 ;
      RECT 407.500000 332.350000 408.500000 333.650000 ;
      RECT 366.500000 332.350000 399.500000 333.650000 ;
      RECT 357.500000 332.350000 358.500000 333.650000 ;
      RECT 316.500000 332.350000 349.500000 333.650000 ;
      RECT 307.500000 332.350000 308.500000 333.650000 ;
      RECT 266.500000 332.350000 299.500000 333.650000 ;
      RECT 257.500000 332.350000 258.500000 333.650000 ;
      RECT 216.500000 332.350000 249.500000 333.650000 ;
      RECT 207.500000 332.350000 208.500000 333.650000 ;
      RECT 166.500000 332.350000 199.500000 333.650000 ;
      RECT 157.500000 332.350000 158.500000 333.650000 ;
      RECT 116.500000 332.350000 149.500000 333.650000 ;
      RECT 107.500000 332.350000 108.500000 333.650000 ;
      RECT 66.500000 332.350000 99.500000 333.650000 ;
      RECT 57.500000 332.350000 58.500000 333.650000 ;
      RECT 29.500000 332.350000 49.500000 333.650000 ;
      RECT 15.500000 332.350000 16.500000 333.650000 ;
      RECT 0.000000 332.350000 2.500000 335.650000 ;
      RECT 1169.500000 331.650000 1186.000000 332.350000 ;
      RECT 1116.500000 331.650000 1156.500000 332.350000 ;
      RECT 1066.500000 331.650000 1108.500000 332.350000 ;
      RECT 1016.500000 331.650000 1058.500000 332.350000 ;
      RECT 966.500000 331.650000 1008.500000 332.350000 ;
      RECT 916.500000 331.650000 958.500000 332.350000 ;
      RECT 866.500000 331.650000 908.500000 332.350000 ;
      RECT 816.500000 331.650000 858.500000 332.350000 ;
      RECT 766.500000 331.650000 808.500000 332.350000 ;
      RECT 716.500000 331.650000 758.500000 332.350000 ;
      RECT 666.500000 331.650000 708.500000 332.350000 ;
      RECT 616.500000 331.650000 658.500000 332.350000 ;
      RECT 566.500000 331.650000 608.500000 332.350000 ;
      RECT 516.500000 331.650000 558.500000 332.350000 ;
      RECT 466.500000 331.650000 508.500000 332.350000 ;
      RECT 416.500000 331.650000 458.500000 332.350000 ;
      RECT 366.500000 331.650000 408.500000 332.350000 ;
      RECT 316.500000 331.650000 358.500000 332.350000 ;
      RECT 266.500000 331.650000 308.500000 332.350000 ;
      RECT 216.500000 331.650000 258.500000 332.350000 ;
      RECT 166.500000 331.650000 208.500000 332.350000 ;
      RECT 116.500000 331.650000 158.500000 332.350000 ;
      RECT 66.500000 331.650000 108.500000 332.350000 ;
      RECT 29.500000 331.650000 58.500000 332.350000 ;
      RECT 0.000000 331.650000 16.500000 332.350000 ;
      RECT 1169.500000 330.350000 1170.500000 331.650000 ;
      RECT 1116.500000 330.350000 1149.500000 331.650000 ;
      RECT 1107.500000 330.350000 1108.500000 331.650000 ;
      RECT 1066.500000 330.350000 1099.500000 331.650000 ;
      RECT 1057.500000 330.350000 1058.500000 331.650000 ;
      RECT 1016.500000 330.350000 1049.500000 331.650000 ;
      RECT 1007.500000 330.350000 1008.500000 331.650000 ;
      RECT 966.500000 330.350000 999.500000 331.650000 ;
      RECT 957.500000 330.350000 958.500000 331.650000 ;
      RECT 916.500000 330.350000 949.500000 331.650000 ;
      RECT 907.500000 330.350000 908.500000 331.650000 ;
      RECT 866.500000 330.350000 899.500000 331.650000 ;
      RECT 857.500000 330.350000 858.500000 331.650000 ;
      RECT 816.500000 330.350000 849.500000 331.650000 ;
      RECT 807.500000 330.350000 808.500000 331.650000 ;
      RECT 766.500000 330.350000 799.500000 331.650000 ;
      RECT 757.500000 330.350000 758.500000 331.650000 ;
      RECT 716.500000 330.350000 749.500000 331.650000 ;
      RECT 707.500000 330.350000 708.500000 331.650000 ;
      RECT 666.500000 330.350000 699.500000 331.650000 ;
      RECT 657.500000 330.350000 658.500000 331.650000 ;
      RECT 616.500000 330.350000 649.500000 331.650000 ;
      RECT 607.500000 330.350000 608.500000 331.650000 ;
      RECT 566.500000 330.350000 599.500000 331.650000 ;
      RECT 557.500000 330.350000 558.500000 331.650000 ;
      RECT 516.500000 330.350000 549.500000 331.650000 ;
      RECT 507.500000 330.350000 508.500000 331.650000 ;
      RECT 466.500000 330.350000 499.500000 331.650000 ;
      RECT 457.500000 330.350000 458.500000 331.650000 ;
      RECT 416.500000 330.350000 449.500000 331.650000 ;
      RECT 407.500000 330.350000 408.500000 331.650000 ;
      RECT 366.500000 330.350000 399.500000 331.650000 ;
      RECT 357.500000 330.350000 358.500000 331.650000 ;
      RECT 316.500000 330.350000 349.500000 331.650000 ;
      RECT 307.500000 330.350000 308.500000 331.650000 ;
      RECT 266.500000 330.350000 299.500000 331.650000 ;
      RECT 257.500000 330.350000 258.500000 331.650000 ;
      RECT 216.500000 330.350000 249.500000 331.650000 ;
      RECT 207.500000 330.350000 208.500000 331.650000 ;
      RECT 166.500000 330.350000 199.500000 331.650000 ;
      RECT 157.500000 330.350000 158.500000 331.650000 ;
      RECT 116.500000 330.350000 149.500000 331.650000 ;
      RECT 107.500000 330.350000 108.500000 331.650000 ;
      RECT 66.500000 330.350000 99.500000 331.650000 ;
      RECT 57.500000 330.350000 58.500000 331.650000 ;
      RECT 29.500000 330.350000 49.500000 331.650000 ;
      RECT 15.500000 330.350000 16.500000 331.650000 ;
      RECT 1157.500000 329.650000 1170.500000 330.350000 ;
      RECT 1107.500000 329.650000 1149.500000 330.350000 ;
      RECT 1057.500000 329.650000 1099.500000 330.350000 ;
      RECT 1007.500000 329.650000 1049.500000 330.350000 ;
      RECT 957.500000 329.650000 999.500000 330.350000 ;
      RECT 907.500000 329.650000 949.500000 330.350000 ;
      RECT 857.500000 329.650000 899.500000 330.350000 ;
      RECT 807.500000 329.650000 849.500000 330.350000 ;
      RECT 757.500000 329.650000 799.500000 330.350000 ;
      RECT 707.500000 329.650000 749.500000 330.350000 ;
      RECT 657.500000 329.650000 699.500000 330.350000 ;
      RECT 607.500000 329.650000 649.500000 330.350000 ;
      RECT 557.500000 329.650000 599.500000 330.350000 ;
      RECT 507.500000 329.650000 549.500000 330.350000 ;
      RECT 457.500000 329.650000 499.500000 330.350000 ;
      RECT 407.500000 329.650000 449.500000 330.350000 ;
      RECT 357.500000 329.650000 399.500000 330.350000 ;
      RECT 307.500000 329.650000 349.500000 330.350000 ;
      RECT 257.500000 329.650000 299.500000 330.350000 ;
      RECT 207.500000 329.650000 249.500000 330.350000 ;
      RECT 157.500000 329.650000 199.500000 330.350000 ;
      RECT 107.500000 329.650000 149.500000 330.350000 ;
      RECT 57.500000 329.650000 99.500000 330.350000 ;
      RECT 15.500000 329.650000 49.500000 330.350000 ;
      RECT 1183.500000 328.350000 1186.000000 331.650000 ;
      RECT 1169.500000 328.350000 1170.500000 329.650000 ;
      RECT 1116.500000 328.350000 1149.500000 329.650000 ;
      RECT 1107.500000 328.350000 1108.500000 329.650000 ;
      RECT 1066.500000 328.350000 1099.500000 329.650000 ;
      RECT 1057.500000 328.350000 1058.500000 329.650000 ;
      RECT 1016.500000 328.350000 1049.500000 329.650000 ;
      RECT 1007.500000 328.350000 1008.500000 329.650000 ;
      RECT 966.500000 328.350000 999.500000 329.650000 ;
      RECT 957.500000 328.350000 958.500000 329.650000 ;
      RECT 916.500000 328.350000 949.500000 329.650000 ;
      RECT 907.500000 328.350000 908.500000 329.650000 ;
      RECT 866.500000 328.350000 899.500000 329.650000 ;
      RECT 857.500000 328.350000 858.500000 329.650000 ;
      RECT 816.500000 328.350000 849.500000 329.650000 ;
      RECT 807.500000 328.350000 808.500000 329.650000 ;
      RECT 766.500000 328.350000 799.500000 329.650000 ;
      RECT 757.500000 328.350000 758.500000 329.650000 ;
      RECT 716.500000 328.350000 749.500000 329.650000 ;
      RECT 707.500000 328.350000 708.500000 329.650000 ;
      RECT 666.500000 328.350000 699.500000 329.650000 ;
      RECT 657.500000 328.350000 658.500000 329.650000 ;
      RECT 616.500000 328.350000 649.500000 329.650000 ;
      RECT 607.500000 328.350000 608.500000 329.650000 ;
      RECT 566.500000 328.350000 599.500000 329.650000 ;
      RECT 557.500000 328.350000 558.500000 329.650000 ;
      RECT 516.500000 328.350000 549.500000 329.650000 ;
      RECT 507.500000 328.350000 508.500000 329.650000 ;
      RECT 466.500000 328.350000 499.500000 329.650000 ;
      RECT 457.500000 328.350000 458.500000 329.650000 ;
      RECT 416.500000 328.350000 449.500000 329.650000 ;
      RECT 407.500000 328.350000 408.500000 329.650000 ;
      RECT 366.500000 328.350000 399.500000 329.650000 ;
      RECT 357.500000 328.350000 358.500000 329.650000 ;
      RECT 316.500000 328.350000 349.500000 329.650000 ;
      RECT 307.500000 328.350000 308.500000 329.650000 ;
      RECT 266.500000 328.350000 299.500000 329.650000 ;
      RECT 257.500000 328.350000 258.500000 329.650000 ;
      RECT 216.500000 328.350000 249.500000 329.650000 ;
      RECT 207.500000 328.350000 208.500000 329.650000 ;
      RECT 166.500000 328.350000 199.500000 329.650000 ;
      RECT 157.500000 328.350000 158.500000 329.650000 ;
      RECT 116.500000 328.350000 149.500000 329.650000 ;
      RECT 107.500000 328.350000 108.500000 329.650000 ;
      RECT 66.500000 328.350000 99.500000 329.650000 ;
      RECT 57.500000 328.350000 58.500000 329.650000 ;
      RECT 29.500000 328.350000 49.500000 329.650000 ;
      RECT 15.500000 328.350000 16.500000 329.650000 ;
      RECT 0.000000 328.350000 2.500000 331.650000 ;
      RECT 1169.500000 327.650000 1186.000000 328.350000 ;
      RECT 1116.500000 327.650000 1156.500000 328.350000 ;
      RECT 1066.500000 327.650000 1108.500000 328.350000 ;
      RECT 1016.500000 327.650000 1058.500000 328.350000 ;
      RECT 966.500000 327.650000 1008.500000 328.350000 ;
      RECT 916.500000 327.650000 958.500000 328.350000 ;
      RECT 866.500000 327.650000 908.500000 328.350000 ;
      RECT 816.500000 327.650000 858.500000 328.350000 ;
      RECT 766.500000 327.650000 808.500000 328.350000 ;
      RECT 716.500000 327.650000 758.500000 328.350000 ;
      RECT 666.500000 327.650000 708.500000 328.350000 ;
      RECT 616.500000 327.650000 658.500000 328.350000 ;
      RECT 566.500000 327.650000 608.500000 328.350000 ;
      RECT 516.500000 327.650000 558.500000 328.350000 ;
      RECT 466.500000 327.650000 508.500000 328.350000 ;
      RECT 416.500000 327.650000 458.500000 328.350000 ;
      RECT 366.500000 327.650000 408.500000 328.350000 ;
      RECT 316.500000 327.650000 358.500000 328.350000 ;
      RECT 266.500000 327.650000 308.500000 328.350000 ;
      RECT 216.500000 327.650000 258.500000 328.350000 ;
      RECT 166.500000 327.650000 208.500000 328.350000 ;
      RECT 116.500000 327.650000 158.500000 328.350000 ;
      RECT 66.500000 327.650000 108.500000 328.350000 ;
      RECT 29.500000 327.650000 58.500000 328.350000 ;
      RECT 0.000000 327.650000 16.500000 328.350000 ;
      RECT 1169.500000 326.350000 1170.500000 327.650000 ;
      RECT 1116.500000 326.350000 1149.500000 327.650000 ;
      RECT 1107.500000 326.350000 1108.500000 327.650000 ;
      RECT 1066.500000 326.350000 1099.500000 327.650000 ;
      RECT 1057.500000 326.350000 1058.500000 327.650000 ;
      RECT 1016.500000 326.350000 1049.500000 327.650000 ;
      RECT 1007.500000 326.350000 1008.500000 327.650000 ;
      RECT 966.500000 326.350000 999.500000 327.650000 ;
      RECT 957.500000 326.350000 958.500000 327.650000 ;
      RECT 916.500000 326.350000 949.500000 327.650000 ;
      RECT 907.500000 326.350000 908.500000 327.650000 ;
      RECT 866.500000 326.350000 899.500000 327.650000 ;
      RECT 857.500000 326.350000 858.500000 327.650000 ;
      RECT 816.500000 326.350000 849.500000 327.650000 ;
      RECT 807.500000 326.350000 808.500000 327.650000 ;
      RECT 766.500000 326.350000 799.500000 327.650000 ;
      RECT 757.500000 326.350000 758.500000 327.650000 ;
      RECT 716.500000 326.350000 749.500000 327.650000 ;
      RECT 707.500000 326.350000 708.500000 327.650000 ;
      RECT 666.500000 326.350000 699.500000 327.650000 ;
      RECT 657.500000 326.350000 658.500000 327.650000 ;
      RECT 616.500000 326.350000 649.500000 327.650000 ;
      RECT 607.500000 326.350000 608.500000 327.650000 ;
      RECT 566.500000 326.350000 599.500000 327.650000 ;
      RECT 557.500000 326.350000 558.500000 327.650000 ;
      RECT 516.500000 326.350000 549.500000 327.650000 ;
      RECT 507.500000 326.350000 508.500000 327.650000 ;
      RECT 466.500000 326.350000 499.500000 327.650000 ;
      RECT 457.500000 326.350000 458.500000 327.650000 ;
      RECT 416.500000 326.350000 449.500000 327.650000 ;
      RECT 407.500000 326.350000 408.500000 327.650000 ;
      RECT 366.500000 326.350000 399.500000 327.650000 ;
      RECT 357.500000 326.350000 358.500000 327.650000 ;
      RECT 316.500000 326.350000 349.500000 327.650000 ;
      RECT 307.500000 326.350000 308.500000 327.650000 ;
      RECT 266.500000 326.350000 299.500000 327.650000 ;
      RECT 257.500000 326.350000 258.500000 327.650000 ;
      RECT 216.500000 326.350000 249.500000 327.650000 ;
      RECT 207.500000 326.350000 208.500000 327.650000 ;
      RECT 166.500000 326.350000 199.500000 327.650000 ;
      RECT 157.500000 326.350000 158.500000 327.650000 ;
      RECT 116.500000 326.350000 149.500000 327.650000 ;
      RECT 107.500000 326.350000 108.500000 327.650000 ;
      RECT 66.500000 326.350000 99.500000 327.650000 ;
      RECT 57.500000 326.350000 58.500000 327.650000 ;
      RECT 29.500000 326.350000 49.500000 327.650000 ;
      RECT 15.500000 326.350000 16.500000 327.650000 ;
      RECT 1157.500000 325.650000 1170.500000 326.350000 ;
      RECT 1107.500000 325.650000 1149.500000 326.350000 ;
      RECT 1057.500000 325.650000 1099.500000 326.350000 ;
      RECT 1007.500000 325.650000 1049.500000 326.350000 ;
      RECT 957.500000 325.650000 999.500000 326.350000 ;
      RECT 907.500000 325.650000 949.500000 326.350000 ;
      RECT 857.500000 325.650000 899.500000 326.350000 ;
      RECT 807.500000 325.650000 849.500000 326.350000 ;
      RECT 757.500000 325.650000 799.500000 326.350000 ;
      RECT 707.500000 325.650000 749.500000 326.350000 ;
      RECT 657.500000 325.650000 699.500000 326.350000 ;
      RECT 607.500000 325.650000 649.500000 326.350000 ;
      RECT 557.500000 325.650000 599.500000 326.350000 ;
      RECT 507.500000 325.650000 549.500000 326.350000 ;
      RECT 457.500000 325.650000 499.500000 326.350000 ;
      RECT 407.500000 325.650000 449.500000 326.350000 ;
      RECT 357.500000 325.650000 399.500000 326.350000 ;
      RECT 307.500000 325.650000 349.500000 326.350000 ;
      RECT 257.500000 325.650000 299.500000 326.350000 ;
      RECT 207.500000 325.650000 249.500000 326.350000 ;
      RECT 157.500000 325.650000 199.500000 326.350000 ;
      RECT 107.500000 325.650000 149.500000 326.350000 ;
      RECT 57.500000 325.650000 99.500000 326.350000 ;
      RECT 15.500000 325.650000 49.500000 326.350000 ;
      RECT 1183.500000 324.350000 1186.000000 327.650000 ;
      RECT 1169.500000 324.350000 1170.500000 325.650000 ;
      RECT 1116.500000 324.350000 1149.500000 325.650000 ;
      RECT 1107.500000 324.350000 1108.500000 325.650000 ;
      RECT 1066.500000 324.350000 1099.500000 325.650000 ;
      RECT 1057.500000 324.350000 1058.500000 325.650000 ;
      RECT 1016.500000 324.350000 1049.500000 325.650000 ;
      RECT 1007.500000 324.350000 1008.500000 325.650000 ;
      RECT 966.500000 324.350000 999.500000 325.650000 ;
      RECT 957.500000 324.350000 958.500000 325.650000 ;
      RECT 916.500000 324.350000 949.500000 325.650000 ;
      RECT 907.500000 324.350000 908.500000 325.650000 ;
      RECT 866.500000 324.350000 899.500000 325.650000 ;
      RECT 857.500000 324.350000 858.500000 325.650000 ;
      RECT 816.500000 324.350000 849.500000 325.650000 ;
      RECT 807.500000 324.350000 808.500000 325.650000 ;
      RECT 766.500000 324.350000 799.500000 325.650000 ;
      RECT 757.500000 324.350000 758.500000 325.650000 ;
      RECT 716.500000 324.350000 749.500000 325.650000 ;
      RECT 707.500000 324.350000 708.500000 325.650000 ;
      RECT 666.500000 324.350000 699.500000 325.650000 ;
      RECT 657.500000 324.350000 658.500000 325.650000 ;
      RECT 616.500000 324.350000 649.500000 325.650000 ;
      RECT 607.500000 324.350000 608.500000 325.650000 ;
      RECT 566.500000 324.350000 599.500000 325.650000 ;
      RECT 557.500000 324.350000 558.500000 325.650000 ;
      RECT 516.500000 324.350000 549.500000 325.650000 ;
      RECT 507.500000 324.350000 508.500000 325.650000 ;
      RECT 466.500000 324.350000 499.500000 325.650000 ;
      RECT 457.500000 324.350000 458.500000 325.650000 ;
      RECT 416.500000 324.350000 449.500000 325.650000 ;
      RECT 407.500000 324.350000 408.500000 325.650000 ;
      RECT 366.500000 324.350000 399.500000 325.650000 ;
      RECT 357.500000 324.350000 358.500000 325.650000 ;
      RECT 316.500000 324.350000 349.500000 325.650000 ;
      RECT 307.500000 324.350000 308.500000 325.650000 ;
      RECT 266.500000 324.350000 299.500000 325.650000 ;
      RECT 257.500000 324.350000 258.500000 325.650000 ;
      RECT 216.500000 324.350000 249.500000 325.650000 ;
      RECT 207.500000 324.350000 208.500000 325.650000 ;
      RECT 166.500000 324.350000 199.500000 325.650000 ;
      RECT 157.500000 324.350000 158.500000 325.650000 ;
      RECT 116.500000 324.350000 149.500000 325.650000 ;
      RECT 107.500000 324.350000 108.500000 325.650000 ;
      RECT 66.500000 324.350000 99.500000 325.650000 ;
      RECT 57.500000 324.350000 58.500000 325.650000 ;
      RECT 29.500000 324.350000 49.500000 325.650000 ;
      RECT 15.500000 324.350000 16.500000 325.650000 ;
      RECT 0.000000 324.350000 2.500000 327.650000 ;
      RECT 1169.500000 323.650000 1186.000000 324.350000 ;
      RECT 1116.500000 323.650000 1156.500000 324.350000 ;
      RECT 1066.500000 323.650000 1108.500000 324.350000 ;
      RECT 1016.500000 323.650000 1058.500000 324.350000 ;
      RECT 966.500000 323.650000 1008.500000 324.350000 ;
      RECT 916.500000 323.650000 958.500000 324.350000 ;
      RECT 866.500000 323.650000 908.500000 324.350000 ;
      RECT 816.500000 323.650000 858.500000 324.350000 ;
      RECT 766.500000 323.650000 808.500000 324.350000 ;
      RECT 716.500000 323.650000 758.500000 324.350000 ;
      RECT 666.500000 323.650000 708.500000 324.350000 ;
      RECT 616.500000 323.650000 658.500000 324.350000 ;
      RECT 566.500000 323.650000 608.500000 324.350000 ;
      RECT 516.500000 323.650000 558.500000 324.350000 ;
      RECT 466.500000 323.650000 508.500000 324.350000 ;
      RECT 416.500000 323.650000 458.500000 324.350000 ;
      RECT 366.500000 323.650000 408.500000 324.350000 ;
      RECT 316.500000 323.650000 358.500000 324.350000 ;
      RECT 266.500000 323.650000 308.500000 324.350000 ;
      RECT 216.500000 323.650000 258.500000 324.350000 ;
      RECT 166.500000 323.650000 208.500000 324.350000 ;
      RECT 116.500000 323.650000 158.500000 324.350000 ;
      RECT 66.500000 323.650000 108.500000 324.350000 ;
      RECT 29.500000 323.650000 58.500000 324.350000 ;
      RECT 0.000000 323.650000 16.500000 324.350000 ;
      RECT 1169.500000 322.350000 1170.500000 323.650000 ;
      RECT 1116.500000 322.350000 1149.500000 323.650000 ;
      RECT 1107.500000 322.350000 1108.500000 323.650000 ;
      RECT 1066.500000 322.350000 1099.500000 323.650000 ;
      RECT 1057.500000 322.350000 1058.500000 323.650000 ;
      RECT 1016.500000 322.350000 1049.500000 323.650000 ;
      RECT 1007.500000 322.350000 1008.500000 323.650000 ;
      RECT 966.500000 322.350000 999.500000 323.650000 ;
      RECT 957.500000 322.350000 958.500000 323.650000 ;
      RECT 916.500000 322.350000 949.500000 323.650000 ;
      RECT 907.500000 322.350000 908.500000 323.650000 ;
      RECT 866.500000 322.350000 899.500000 323.650000 ;
      RECT 857.500000 322.350000 858.500000 323.650000 ;
      RECT 816.500000 322.350000 849.500000 323.650000 ;
      RECT 807.500000 322.350000 808.500000 323.650000 ;
      RECT 766.500000 322.350000 799.500000 323.650000 ;
      RECT 757.500000 322.350000 758.500000 323.650000 ;
      RECT 716.500000 322.350000 749.500000 323.650000 ;
      RECT 707.500000 322.350000 708.500000 323.650000 ;
      RECT 666.500000 322.350000 699.500000 323.650000 ;
      RECT 657.500000 322.350000 658.500000 323.650000 ;
      RECT 616.500000 322.350000 649.500000 323.650000 ;
      RECT 607.500000 322.350000 608.500000 323.650000 ;
      RECT 566.500000 322.350000 599.500000 323.650000 ;
      RECT 557.500000 322.350000 558.500000 323.650000 ;
      RECT 516.500000 322.350000 549.500000 323.650000 ;
      RECT 507.500000 322.350000 508.500000 323.650000 ;
      RECT 466.500000 322.350000 499.500000 323.650000 ;
      RECT 457.500000 322.350000 458.500000 323.650000 ;
      RECT 416.500000 322.350000 449.500000 323.650000 ;
      RECT 407.500000 322.350000 408.500000 323.650000 ;
      RECT 366.500000 322.350000 399.500000 323.650000 ;
      RECT 357.500000 322.350000 358.500000 323.650000 ;
      RECT 316.500000 322.350000 349.500000 323.650000 ;
      RECT 307.500000 322.350000 308.500000 323.650000 ;
      RECT 266.500000 322.350000 299.500000 323.650000 ;
      RECT 257.500000 322.350000 258.500000 323.650000 ;
      RECT 216.500000 322.350000 249.500000 323.650000 ;
      RECT 207.500000 322.350000 208.500000 323.650000 ;
      RECT 166.500000 322.350000 199.500000 323.650000 ;
      RECT 157.500000 322.350000 158.500000 323.650000 ;
      RECT 116.500000 322.350000 149.500000 323.650000 ;
      RECT 107.500000 322.350000 108.500000 323.650000 ;
      RECT 66.500000 322.350000 99.500000 323.650000 ;
      RECT 57.500000 322.350000 58.500000 323.650000 ;
      RECT 29.500000 322.350000 49.500000 323.650000 ;
      RECT 15.500000 322.350000 16.500000 323.650000 ;
      RECT 1157.500000 321.650000 1170.500000 322.350000 ;
      RECT 1107.500000 321.650000 1149.500000 322.350000 ;
      RECT 1057.500000 321.650000 1099.500000 322.350000 ;
      RECT 1007.500000 321.650000 1049.500000 322.350000 ;
      RECT 957.500000 321.650000 999.500000 322.350000 ;
      RECT 907.500000 321.650000 949.500000 322.350000 ;
      RECT 857.500000 321.650000 899.500000 322.350000 ;
      RECT 807.500000 321.650000 849.500000 322.350000 ;
      RECT 757.500000 321.650000 799.500000 322.350000 ;
      RECT 707.500000 321.650000 749.500000 322.350000 ;
      RECT 657.500000 321.650000 699.500000 322.350000 ;
      RECT 607.500000 321.650000 649.500000 322.350000 ;
      RECT 557.500000 321.650000 599.500000 322.350000 ;
      RECT 507.500000 321.650000 549.500000 322.350000 ;
      RECT 457.500000 321.650000 499.500000 322.350000 ;
      RECT 407.500000 321.650000 449.500000 322.350000 ;
      RECT 357.500000 321.650000 399.500000 322.350000 ;
      RECT 307.500000 321.650000 349.500000 322.350000 ;
      RECT 257.500000 321.650000 299.500000 322.350000 ;
      RECT 207.500000 321.650000 249.500000 322.350000 ;
      RECT 157.500000 321.650000 199.500000 322.350000 ;
      RECT 107.500000 321.650000 149.500000 322.350000 ;
      RECT 57.500000 321.650000 99.500000 322.350000 ;
      RECT 15.500000 321.650000 49.500000 322.350000 ;
      RECT 1183.500000 320.350000 1186.000000 323.650000 ;
      RECT 1169.500000 320.350000 1170.500000 321.650000 ;
      RECT 1116.500000 320.350000 1149.500000 321.650000 ;
      RECT 1107.500000 320.350000 1108.500000 321.650000 ;
      RECT 1066.500000 320.350000 1099.500000 321.650000 ;
      RECT 1057.500000 320.350000 1058.500000 321.650000 ;
      RECT 1016.500000 320.350000 1049.500000 321.650000 ;
      RECT 1007.500000 320.350000 1008.500000 321.650000 ;
      RECT 966.500000 320.350000 999.500000 321.650000 ;
      RECT 957.500000 320.350000 958.500000 321.650000 ;
      RECT 916.500000 320.350000 949.500000 321.650000 ;
      RECT 907.500000 320.350000 908.500000 321.650000 ;
      RECT 866.500000 320.350000 899.500000 321.650000 ;
      RECT 857.500000 320.350000 858.500000 321.650000 ;
      RECT 816.500000 320.350000 849.500000 321.650000 ;
      RECT 807.500000 320.350000 808.500000 321.650000 ;
      RECT 766.500000 320.350000 799.500000 321.650000 ;
      RECT 757.500000 320.350000 758.500000 321.650000 ;
      RECT 716.500000 320.350000 749.500000 321.650000 ;
      RECT 707.500000 320.350000 708.500000 321.650000 ;
      RECT 666.500000 320.350000 699.500000 321.650000 ;
      RECT 657.500000 320.350000 658.500000 321.650000 ;
      RECT 616.500000 320.350000 649.500000 321.650000 ;
      RECT 607.500000 320.350000 608.500000 321.650000 ;
      RECT 566.500000 320.350000 599.500000 321.650000 ;
      RECT 557.500000 320.350000 558.500000 321.650000 ;
      RECT 516.500000 320.350000 549.500000 321.650000 ;
      RECT 507.500000 320.350000 508.500000 321.650000 ;
      RECT 466.500000 320.350000 499.500000 321.650000 ;
      RECT 457.500000 320.350000 458.500000 321.650000 ;
      RECT 416.500000 320.350000 449.500000 321.650000 ;
      RECT 407.500000 320.350000 408.500000 321.650000 ;
      RECT 366.500000 320.350000 399.500000 321.650000 ;
      RECT 357.500000 320.350000 358.500000 321.650000 ;
      RECT 316.500000 320.350000 349.500000 321.650000 ;
      RECT 307.500000 320.350000 308.500000 321.650000 ;
      RECT 266.500000 320.350000 299.500000 321.650000 ;
      RECT 257.500000 320.350000 258.500000 321.650000 ;
      RECT 216.500000 320.350000 249.500000 321.650000 ;
      RECT 207.500000 320.350000 208.500000 321.650000 ;
      RECT 166.500000 320.350000 199.500000 321.650000 ;
      RECT 157.500000 320.350000 158.500000 321.650000 ;
      RECT 116.500000 320.350000 149.500000 321.650000 ;
      RECT 107.500000 320.350000 108.500000 321.650000 ;
      RECT 66.500000 320.350000 99.500000 321.650000 ;
      RECT 57.500000 320.350000 58.500000 321.650000 ;
      RECT 29.500000 320.350000 49.500000 321.650000 ;
      RECT 15.500000 320.350000 16.500000 321.650000 ;
      RECT 0.000000 320.350000 2.500000 323.650000 ;
      RECT 1169.500000 319.650000 1186.000000 320.350000 ;
      RECT 1116.500000 319.650000 1156.500000 320.350000 ;
      RECT 1066.500000 319.650000 1108.500000 320.350000 ;
      RECT 1016.500000 319.650000 1058.500000 320.350000 ;
      RECT 966.500000 319.650000 1008.500000 320.350000 ;
      RECT 916.500000 319.650000 958.500000 320.350000 ;
      RECT 866.500000 319.650000 908.500000 320.350000 ;
      RECT 816.500000 319.650000 858.500000 320.350000 ;
      RECT 766.500000 319.650000 808.500000 320.350000 ;
      RECT 716.500000 319.650000 758.500000 320.350000 ;
      RECT 666.500000 319.650000 708.500000 320.350000 ;
      RECT 616.500000 319.650000 658.500000 320.350000 ;
      RECT 566.500000 319.650000 608.500000 320.350000 ;
      RECT 516.500000 319.650000 558.500000 320.350000 ;
      RECT 466.500000 319.650000 508.500000 320.350000 ;
      RECT 366.500000 319.650000 408.500000 320.350000 ;
      RECT 316.500000 319.650000 358.500000 320.350000 ;
      RECT 266.500000 319.650000 308.500000 320.350000 ;
      RECT 216.500000 319.650000 258.500000 320.350000 ;
      RECT 166.500000 319.650000 208.500000 320.350000 ;
      RECT 116.500000 319.650000 158.500000 320.350000 ;
      RECT 66.500000 319.650000 108.500000 320.350000 ;
      RECT 29.500000 319.650000 58.500000 320.350000 ;
      RECT 0.000000 319.650000 16.500000 320.350000 ;
      RECT 1169.500000 318.350000 1170.500000 319.650000 ;
      RECT 1116.500000 318.350000 1149.500000 319.650000 ;
      RECT 1107.500000 318.350000 1108.500000 319.650000 ;
      RECT 1066.500000 318.350000 1099.500000 319.650000 ;
      RECT 1057.500000 318.350000 1058.500000 319.650000 ;
      RECT 1016.500000 318.350000 1049.500000 319.650000 ;
      RECT 1007.500000 318.350000 1008.500000 319.650000 ;
      RECT 966.500000 318.350000 999.500000 319.650000 ;
      RECT 957.500000 318.350000 958.500000 319.650000 ;
      RECT 916.500000 318.350000 949.500000 319.650000 ;
      RECT 907.500000 318.350000 908.500000 319.650000 ;
      RECT 866.500000 318.350000 899.500000 319.650000 ;
      RECT 857.500000 318.350000 858.500000 319.650000 ;
      RECT 816.500000 318.350000 849.500000 319.650000 ;
      RECT 807.500000 318.350000 808.500000 319.650000 ;
      RECT 766.500000 318.350000 799.500000 319.650000 ;
      RECT 757.500000 318.350000 758.500000 319.650000 ;
      RECT 716.500000 318.350000 749.500000 319.650000 ;
      RECT 707.500000 318.350000 708.500000 319.650000 ;
      RECT 666.500000 318.350000 699.500000 319.650000 ;
      RECT 657.500000 318.350000 658.500000 319.650000 ;
      RECT 616.500000 318.350000 649.500000 319.650000 ;
      RECT 607.500000 318.350000 608.500000 319.650000 ;
      RECT 566.500000 318.350000 599.500000 319.650000 ;
      RECT 557.500000 318.350000 558.500000 319.650000 ;
      RECT 516.500000 318.350000 549.500000 319.650000 ;
      RECT 507.500000 318.350000 508.500000 319.650000 ;
      RECT 466.500000 318.350000 499.500000 319.650000 ;
      RECT 416.500000 318.350000 458.500000 320.350000 ;
      RECT 407.500000 318.350000 408.500000 319.650000 ;
      RECT 366.500000 318.350000 399.500000 319.650000 ;
      RECT 357.500000 318.350000 358.500000 319.650000 ;
      RECT 316.500000 318.350000 349.500000 319.650000 ;
      RECT 307.500000 318.350000 308.500000 319.650000 ;
      RECT 266.500000 318.350000 299.500000 319.650000 ;
      RECT 257.500000 318.350000 258.500000 319.650000 ;
      RECT 216.500000 318.350000 249.500000 319.650000 ;
      RECT 207.500000 318.350000 208.500000 319.650000 ;
      RECT 166.500000 318.350000 199.500000 319.650000 ;
      RECT 157.500000 318.350000 158.500000 319.650000 ;
      RECT 116.500000 318.350000 149.500000 319.650000 ;
      RECT 107.500000 318.350000 108.500000 319.650000 ;
      RECT 66.500000 318.350000 99.500000 319.650000 ;
      RECT 57.500000 318.350000 58.500000 319.650000 ;
      RECT 29.500000 318.350000 49.500000 319.650000 ;
      RECT 15.500000 318.350000 16.500000 319.650000 ;
      RECT 1157.500000 317.650000 1170.500000 318.350000 ;
      RECT 1107.500000 317.650000 1149.500000 318.350000 ;
      RECT 1057.500000 317.650000 1099.500000 318.350000 ;
      RECT 1007.500000 317.650000 1049.500000 318.350000 ;
      RECT 957.500000 317.650000 999.500000 318.350000 ;
      RECT 907.500000 317.650000 949.500000 318.350000 ;
      RECT 857.500000 317.650000 899.500000 318.350000 ;
      RECT 807.500000 317.650000 849.500000 318.350000 ;
      RECT 757.500000 317.650000 799.500000 318.350000 ;
      RECT 707.500000 317.650000 749.500000 318.350000 ;
      RECT 657.500000 317.650000 699.500000 318.350000 ;
      RECT 607.500000 317.650000 649.500000 318.350000 ;
      RECT 557.500000 317.650000 599.500000 318.350000 ;
      RECT 507.500000 317.650000 549.500000 318.350000 ;
      RECT 407.500000 317.650000 499.500000 318.350000 ;
      RECT 357.500000 317.650000 399.500000 318.350000 ;
      RECT 307.500000 317.650000 349.500000 318.350000 ;
      RECT 257.500000 317.650000 299.500000 318.350000 ;
      RECT 207.500000 317.650000 249.500000 318.350000 ;
      RECT 157.500000 317.650000 199.500000 318.350000 ;
      RECT 107.500000 317.650000 149.500000 318.350000 ;
      RECT 57.500000 317.650000 99.500000 318.350000 ;
      RECT 15.500000 317.650000 49.500000 318.350000 ;
      RECT 1183.500000 316.350000 1186.000000 319.650000 ;
      RECT 1169.500000 316.350000 1170.500000 317.650000 ;
      RECT 1116.500000 316.350000 1149.500000 317.650000 ;
      RECT 1107.500000 316.350000 1108.500000 317.650000 ;
      RECT 1066.500000 316.350000 1099.500000 317.650000 ;
      RECT 1057.500000 316.350000 1058.500000 317.650000 ;
      RECT 1016.500000 316.350000 1049.500000 317.650000 ;
      RECT 1007.500000 316.350000 1008.500000 317.650000 ;
      RECT 966.500000 316.350000 999.500000 317.650000 ;
      RECT 957.500000 316.350000 958.500000 317.650000 ;
      RECT 916.500000 316.350000 949.500000 317.650000 ;
      RECT 907.500000 316.350000 908.500000 317.650000 ;
      RECT 866.500000 316.350000 899.500000 317.650000 ;
      RECT 857.500000 316.350000 858.500000 317.650000 ;
      RECT 816.500000 316.350000 849.500000 317.650000 ;
      RECT 807.500000 316.350000 808.500000 317.650000 ;
      RECT 766.500000 316.350000 799.500000 317.650000 ;
      RECT 757.500000 316.350000 758.500000 317.650000 ;
      RECT 716.500000 316.350000 749.500000 317.650000 ;
      RECT 707.500000 316.350000 708.500000 317.650000 ;
      RECT 666.500000 316.350000 699.500000 317.650000 ;
      RECT 657.500000 316.350000 658.500000 317.650000 ;
      RECT 616.500000 316.350000 649.500000 317.650000 ;
      RECT 607.500000 316.350000 608.500000 317.650000 ;
      RECT 566.500000 316.350000 599.500000 317.650000 ;
      RECT 557.500000 316.350000 558.500000 317.650000 ;
      RECT 516.500000 316.350000 549.500000 317.650000 ;
      RECT 507.500000 316.350000 508.500000 317.650000 ;
      RECT 416.500000 316.350000 499.500000 317.650000 ;
      RECT 407.500000 316.350000 408.500000 317.650000 ;
      RECT 366.500000 316.350000 399.500000 317.650000 ;
      RECT 357.500000 316.350000 358.500000 317.650000 ;
      RECT 316.500000 316.350000 349.500000 317.650000 ;
      RECT 307.500000 316.350000 308.500000 317.650000 ;
      RECT 266.500000 316.350000 299.500000 317.650000 ;
      RECT 257.500000 316.350000 258.500000 317.650000 ;
      RECT 216.500000 316.350000 249.500000 317.650000 ;
      RECT 207.500000 316.350000 208.500000 317.650000 ;
      RECT 166.500000 316.350000 199.500000 317.650000 ;
      RECT 157.500000 316.350000 158.500000 317.650000 ;
      RECT 116.500000 316.350000 149.500000 317.650000 ;
      RECT 107.500000 316.350000 108.500000 317.650000 ;
      RECT 66.500000 316.350000 99.500000 317.650000 ;
      RECT 57.500000 316.350000 58.500000 317.650000 ;
      RECT 29.500000 316.350000 49.500000 317.650000 ;
      RECT 15.500000 316.350000 16.500000 317.650000 ;
      RECT 0.000000 316.350000 2.500000 319.650000 ;
      RECT 1169.500000 315.650000 1186.000000 316.350000 ;
      RECT 1116.500000 315.650000 1156.500000 316.350000 ;
      RECT 1066.500000 315.650000 1108.500000 316.350000 ;
      RECT 1016.500000 315.650000 1058.500000 316.350000 ;
      RECT 966.500000 315.650000 1008.500000 316.350000 ;
      RECT 916.500000 315.650000 958.500000 316.350000 ;
      RECT 866.500000 315.650000 908.500000 316.350000 ;
      RECT 816.500000 315.650000 858.500000 316.350000 ;
      RECT 766.500000 315.650000 808.500000 316.350000 ;
      RECT 716.500000 315.650000 758.500000 316.350000 ;
      RECT 666.500000 315.650000 708.500000 316.350000 ;
      RECT 616.500000 315.650000 658.500000 316.350000 ;
      RECT 566.500000 315.650000 608.500000 316.350000 ;
      RECT 516.500000 315.650000 558.500000 316.350000 ;
      RECT 416.500000 315.650000 508.500000 316.350000 ;
      RECT 366.500000 315.650000 408.500000 316.350000 ;
      RECT 316.500000 315.650000 358.500000 316.350000 ;
      RECT 266.500000 315.650000 308.500000 316.350000 ;
      RECT 216.500000 315.650000 258.500000 316.350000 ;
      RECT 166.500000 315.650000 208.500000 316.350000 ;
      RECT 116.500000 315.650000 158.500000 316.350000 ;
      RECT 66.500000 315.650000 108.500000 316.350000 ;
      RECT 29.500000 315.650000 58.500000 316.350000 ;
      RECT 0.000000 315.650000 16.500000 316.350000 ;
      RECT 1169.500000 314.350000 1170.500000 315.650000 ;
      RECT 1116.500000 314.350000 1149.500000 315.650000 ;
      RECT 1107.500000 314.350000 1108.500000 315.650000 ;
      RECT 1066.500000 314.350000 1099.500000 315.650000 ;
      RECT 1057.500000 314.350000 1058.500000 315.650000 ;
      RECT 1016.500000 314.350000 1049.500000 315.650000 ;
      RECT 1007.500000 314.350000 1008.500000 315.650000 ;
      RECT 966.500000 314.350000 999.500000 315.650000 ;
      RECT 957.500000 314.350000 958.500000 315.650000 ;
      RECT 916.500000 314.350000 949.500000 315.650000 ;
      RECT 907.500000 314.350000 908.500000 315.650000 ;
      RECT 866.500000 314.350000 899.500000 315.650000 ;
      RECT 857.500000 314.350000 858.500000 315.650000 ;
      RECT 816.500000 314.350000 849.500000 315.650000 ;
      RECT 807.500000 314.350000 808.500000 315.650000 ;
      RECT 766.500000 314.350000 799.500000 315.650000 ;
      RECT 757.500000 314.350000 758.500000 315.650000 ;
      RECT 716.500000 314.350000 749.500000 315.650000 ;
      RECT 707.500000 314.350000 708.500000 315.650000 ;
      RECT 666.500000 314.350000 699.500000 315.650000 ;
      RECT 657.500000 314.350000 658.500000 315.650000 ;
      RECT 616.500000 314.350000 649.500000 315.650000 ;
      RECT 607.500000 314.350000 608.500000 315.650000 ;
      RECT 566.500000 314.350000 599.500000 315.650000 ;
      RECT 557.500000 314.350000 558.500000 315.650000 ;
      RECT 516.500000 314.350000 549.500000 315.650000 ;
      RECT 507.500000 314.350000 508.500000 315.650000 ;
      RECT 416.500000 314.350000 499.500000 315.650000 ;
      RECT 407.500000 314.350000 408.500000 315.650000 ;
      RECT 366.500000 314.350000 399.500000 315.650000 ;
      RECT 357.500000 314.350000 358.500000 315.650000 ;
      RECT 316.500000 314.350000 349.500000 315.650000 ;
      RECT 307.500000 314.350000 308.500000 315.650000 ;
      RECT 266.500000 314.350000 299.500000 315.650000 ;
      RECT 257.500000 314.350000 258.500000 315.650000 ;
      RECT 216.500000 314.350000 249.500000 315.650000 ;
      RECT 207.500000 314.350000 208.500000 315.650000 ;
      RECT 166.500000 314.350000 199.500000 315.650000 ;
      RECT 157.500000 314.350000 158.500000 315.650000 ;
      RECT 116.500000 314.350000 149.500000 315.650000 ;
      RECT 107.500000 314.350000 108.500000 315.650000 ;
      RECT 66.500000 314.350000 99.500000 315.650000 ;
      RECT 57.500000 314.350000 58.500000 315.650000 ;
      RECT 29.500000 314.350000 49.500000 315.650000 ;
      RECT 15.500000 314.350000 16.500000 315.650000 ;
      RECT 1157.500000 313.650000 1170.500000 314.350000 ;
      RECT 1107.500000 313.650000 1149.500000 314.350000 ;
      RECT 1057.500000 313.650000 1099.500000 314.350000 ;
      RECT 1007.500000 313.650000 1049.500000 314.350000 ;
      RECT 957.500000 313.650000 999.500000 314.350000 ;
      RECT 907.500000 313.650000 949.500000 314.350000 ;
      RECT 857.500000 313.650000 899.500000 314.350000 ;
      RECT 807.500000 313.650000 849.500000 314.350000 ;
      RECT 757.500000 313.650000 799.500000 314.350000 ;
      RECT 707.500000 313.650000 749.500000 314.350000 ;
      RECT 657.500000 313.650000 699.500000 314.350000 ;
      RECT 607.500000 313.650000 649.500000 314.350000 ;
      RECT 557.500000 313.650000 599.500000 314.350000 ;
      RECT 507.500000 313.650000 549.500000 314.350000 ;
      RECT 407.500000 313.650000 499.500000 314.350000 ;
      RECT 357.500000 313.650000 399.500000 314.350000 ;
      RECT 307.500000 313.650000 349.500000 314.350000 ;
      RECT 257.500000 313.650000 299.500000 314.350000 ;
      RECT 207.500000 313.650000 249.500000 314.350000 ;
      RECT 157.500000 313.650000 199.500000 314.350000 ;
      RECT 107.500000 313.650000 149.500000 314.350000 ;
      RECT 57.500000 313.650000 99.500000 314.350000 ;
      RECT 15.500000 313.650000 49.500000 314.350000 ;
      RECT 1183.500000 312.350000 1186.000000 315.650000 ;
      RECT 1169.500000 312.350000 1170.500000 313.650000 ;
      RECT 1116.500000 312.350000 1149.500000 313.650000 ;
      RECT 1107.500000 312.350000 1108.500000 313.650000 ;
      RECT 1066.500000 312.350000 1099.500000 313.650000 ;
      RECT 1057.500000 312.350000 1058.500000 313.650000 ;
      RECT 1016.500000 312.350000 1049.500000 313.650000 ;
      RECT 1007.500000 312.350000 1008.500000 313.650000 ;
      RECT 966.500000 312.350000 999.500000 313.650000 ;
      RECT 957.500000 312.350000 958.500000 313.650000 ;
      RECT 916.500000 312.350000 949.500000 313.650000 ;
      RECT 907.500000 312.350000 908.500000 313.650000 ;
      RECT 866.500000 312.350000 899.500000 313.650000 ;
      RECT 857.500000 312.350000 858.500000 313.650000 ;
      RECT 816.500000 312.350000 849.500000 313.650000 ;
      RECT 807.500000 312.350000 808.500000 313.650000 ;
      RECT 766.500000 312.350000 799.500000 313.650000 ;
      RECT 757.500000 312.350000 758.500000 313.650000 ;
      RECT 716.500000 312.350000 749.500000 313.650000 ;
      RECT 707.500000 312.350000 708.500000 313.650000 ;
      RECT 666.500000 312.350000 699.500000 313.650000 ;
      RECT 657.500000 312.350000 658.500000 313.650000 ;
      RECT 616.500000 312.350000 649.500000 313.650000 ;
      RECT 607.500000 312.350000 608.500000 313.650000 ;
      RECT 566.500000 312.350000 599.500000 313.650000 ;
      RECT 557.500000 312.350000 558.500000 313.650000 ;
      RECT 516.500000 312.350000 549.500000 313.650000 ;
      RECT 507.500000 312.350000 508.500000 313.650000 ;
      RECT 416.500000 312.350000 499.500000 313.650000 ;
      RECT 407.500000 312.350000 408.500000 313.650000 ;
      RECT 366.500000 312.350000 399.500000 313.650000 ;
      RECT 357.500000 312.350000 358.500000 313.650000 ;
      RECT 316.500000 312.350000 349.500000 313.650000 ;
      RECT 307.500000 312.350000 308.500000 313.650000 ;
      RECT 266.500000 312.350000 299.500000 313.650000 ;
      RECT 257.500000 312.350000 258.500000 313.650000 ;
      RECT 216.500000 312.350000 249.500000 313.650000 ;
      RECT 207.500000 312.350000 208.500000 313.650000 ;
      RECT 166.500000 312.350000 199.500000 313.650000 ;
      RECT 157.500000 312.350000 158.500000 313.650000 ;
      RECT 116.500000 312.350000 149.500000 313.650000 ;
      RECT 107.500000 312.350000 108.500000 313.650000 ;
      RECT 66.500000 312.350000 99.500000 313.650000 ;
      RECT 57.500000 312.350000 58.500000 313.650000 ;
      RECT 29.500000 312.350000 49.500000 313.650000 ;
      RECT 15.500000 312.350000 16.500000 313.650000 ;
      RECT 0.000000 312.350000 2.500000 315.650000 ;
      RECT 1169.500000 311.650000 1186.000000 312.350000 ;
      RECT 1116.500000 311.650000 1156.500000 312.350000 ;
      RECT 1066.500000 311.650000 1108.500000 312.350000 ;
      RECT 1016.500000 311.650000 1058.500000 312.350000 ;
      RECT 966.500000 311.650000 1008.500000 312.350000 ;
      RECT 916.500000 311.650000 958.500000 312.350000 ;
      RECT 866.500000 311.650000 908.500000 312.350000 ;
      RECT 816.500000 311.650000 858.500000 312.350000 ;
      RECT 766.500000 311.650000 808.500000 312.350000 ;
      RECT 716.500000 311.650000 758.500000 312.350000 ;
      RECT 666.500000 311.650000 708.500000 312.350000 ;
      RECT 616.500000 311.650000 658.500000 312.350000 ;
      RECT 566.500000 311.650000 608.500000 312.350000 ;
      RECT 516.500000 311.650000 558.500000 312.350000 ;
      RECT 416.500000 311.650000 508.500000 312.350000 ;
      RECT 366.500000 311.650000 408.500000 312.350000 ;
      RECT 316.500000 311.650000 358.500000 312.350000 ;
      RECT 266.500000 311.650000 308.500000 312.350000 ;
      RECT 216.500000 311.650000 258.500000 312.350000 ;
      RECT 166.500000 311.650000 208.500000 312.350000 ;
      RECT 116.500000 311.650000 158.500000 312.350000 ;
      RECT 66.500000 311.650000 108.500000 312.350000 ;
      RECT 29.500000 311.650000 58.500000 312.350000 ;
      RECT 0.000000 311.650000 16.500000 312.350000 ;
      RECT 0.000000 311.170000 2.500000 311.650000 ;
      RECT 1183.500000 311.165000 1186.000000 311.650000 ;
      RECT 1169.500000 310.350000 1170.500000 311.650000 ;
      RECT 1116.500000 310.350000 1149.500000 311.650000 ;
      RECT 1107.500000 310.350000 1108.500000 311.650000 ;
      RECT 1066.500000 310.350000 1099.500000 311.650000 ;
      RECT 1057.500000 310.350000 1058.500000 311.650000 ;
      RECT 1016.500000 310.350000 1049.500000 311.650000 ;
      RECT 1007.500000 310.350000 1008.500000 311.650000 ;
      RECT 966.500000 310.350000 999.500000 311.650000 ;
      RECT 957.500000 310.350000 958.500000 311.650000 ;
      RECT 916.500000 310.350000 949.500000 311.650000 ;
      RECT 907.500000 310.350000 908.500000 311.650000 ;
      RECT 866.500000 310.350000 899.500000 311.650000 ;
      RECT 857.500000 310.350000 858.500000 311.650000 ;
      RECT 816.500000 310.350000 849.500000 311.650000 ;
      RECT 807.500000 310.350000 808.500000 311.650000 ;
      RECT 766.500000 310.350000 799.500000 311.650000 ;
      RECT 757.500000 310.350000 758.500000 311.650000 ;
      RECT 716.500000 310.350000 749.500000 311.650000 ;
      RECT 707.500000 310.350000 708.500000 311.650000 ;
      RECT 666.500000 310.350000 699.500000 311.650000 ;
      RECT 657.500000 310.350000 658.500000 311.650000 ;
      RECT 616.500000 310.350000 649.500000 311.650000 ;
      RECT 607.500000 310.350000 608.500000 311.650000 ;
      RECT 566.500000 310.350000 599.500000 311.650000 ;
      RECT 557.500000 310.350000 558.500000 311.650000 ;
      RECT 516.500000 310.350000 549.500000 311.650000 ;
      RECT 507.500000 310.350000 508.500000 311.650000 ;
      RECT 416.500000 310.350000 499.500000 311.650000 ;
      RECT 407.500000 310.350000 408.500000 311.650000 ;
      RECT 366.500000 310.350000 399.500000 311.650000 ;
      RECT 357.500000 310.350000 358.500000 311.650000 ;
      RECT 316.500000 310.350000 349.500000 311.650000 ;
      RECT 307.500000 310.350000 308.500000 311.650000 ;
      RECT 266.500000 310.350000 299.500000 311.650000 ;
      RECT 257.500000 310.350000 258.500000 311.650000 ;
      RECT 216.500000 310.350000 249.500000 311.650000 ;
      RECT 207.500000 310.350000 208.500000 311.650000 ;
      RECT 166.500000 310.350000 199.500000 311.650000 ;
      RECT 157.500000 310.350000 158.500000 311.650000 ;
      RECT 116.500000 310.350000 149.500000 311.650000 ;
      RECT 107.500000 310.350000 108.500000 311.650000 ;
      RECT 66.500000 310.350000 99.500000 311.650000 ;
      RECT 57.500000 310.350000 58.500000 311.650000 ;
      RECT 29.500000 310.350000 49.500000 311.650000 ;
      RECT 15.500000 310.350000 16.500000 311.650000 ;
      RECT 1157.500000 309.650000 1170.500000 310.350000 ;
      RECT 1107.500000 309.650000 1149.500000 310.350000 ;
      RECT 1057.500000 309.650000 1099.500000 310.350000 ;
      RECT 1007.500000 309.650000 1049.500000 310.350000 ;
      RECT 957.500000 309.650000 999.500000 310.350000 ;
      RECT 907.500000 309.650000 949.500000 310.350000 ;
      RECT 857.500000 309.650000 899.500000 310.350000 ;
      RECT 807.500000 309.650000 849.500000 310.350000 ;
      RECT 757.500000 309.650000 799.500000 310.350000 ;
      RECT 707.500000 309.650000 749.500000 310.350000 ;
      RECT 657.500000 309.650000 699.500000 310.350000 ;
      RECT 607.500000 309.650000 649.500000 310.350000 ;
      RECT 557.500000 309.650000 599.500000 310.350000 ;
      RECT 507.500000 309.650000 549.500000 310.350000 ;
      RECT 407.500000 309.650000 499.500000 310.350000 ;
      RECT 357.500000 309.650000 399.500000 310.350000 ;
      RECT 307.500000 309.650000 349.500000 310.350000 ;
      RECT 257.500000 309.650000 299.500000 310.350000 ;
      RECT 207.500000 309.650000 249.500000 310.350000 ;
      RECT 157.500000 309.650000 199.500000 310.350000 ;
      RECT 107.500000 309.650000 149.500000 310.350000 ;
      RECT 57.500000 309.650000 99.500000 310.350000 ;
      RECT 15.500000 309.650000 49.500000 310.350000 ;
      RECT 1183.500000 308.350000 1183.980000 311.165000 ;
      RECT 1169.500000 308.350000 1170.500000 309.650000 ;
      RECT 1116.500000 308.350000 1149.500000 309.650000 ;
      RECT 1107.500000 308.350000 1108.500000 309.650000 ;
      RECT 1066.500000 308.350000 1099.500000 309.650000 ;
      RECT 1057.500000 308.350000 1058.500000 309.650000 ;
      RECT 1016.500000 308.350000 1049.500000 309.650000 ;
      RECT 1007.500000 308.350000 1008.500000 309.650000 ;
      RECT 966.500000 308.350000 999.500000 309.650000 ;
      RECT 957.500000 308.350000 958.500000 309.650000 ;
      RECT 916.500000 308.350000 949.500000 309.650000 ;
      RECT 907.500000 308.350000 908.500000 309.650000 ;
      RECT 866.500000 308.350000 899.500000 309.650000 ;
      RECT 857.500000 308.350000 858.500000 309.650000 ;
      RECT 816.500000 308.350000 849.500000 309.650000 ;
      RECT 807.500000 308.350000 808.500000 309.650000 ;
      RECT 766.500000 308.350000 799.500000 309.650000 ;
      RECT 757.500000 308.350000 758.500000 309.650000 ;
      RECT 716.500000 308.350000 749.500000 309.650000 ;
      RECT 707.500000 308.350000 708.500000 309.650000 ;
      RECT 666.500000 308.350000 699.500000 309.650000 ;
      RECT 657.500000 308.350000 658.500000 309.650000 ;
      RECT 616.500000 308.350000 649.500000 309.650000 ;
      RECT 607.500000 308.350000 608.500000 309.650000 ;
      RECT 566.500000 308.350000 599.500000 309.650000 ;
      RECT 557.500000 308.350000 558.500000 309.650000 ;
      RECT 516.500000 308.350000 549.500000 309.650000 ;
      RECT 507.500000 308.350000 508.500000 309.650000 ;
      RECT 416.500000 308.350000 499.500000 309.650000 ;
      RECT 407.500000 308.350000 408.500000 309.650000 ;
      RECT 366.500000 308.350000 399.500000 309.650000 ;
      RECT 357.500000 308.350000 358.500000 309.650000 ;
      RECT 316.500000 308.350000 349.500000 309.650000 ;
      RECT 307.500000 308.350000 308.500000 309.650000 ;
      RECT 266.500000 308.350000 299.500000 309.650000 ;
      RECT 257.500000 308.350000 258.500000 309.650000 ;
      RECT 216.500000 308.350000 249.500000 309.650000 ;
      RECT 207.500000 308.350000 208.500000 309.650000 ;
      RECT 166.500000 308.350000 199.500000 309.650000 ;
      RECT 157.500000 308.350000 158.500000 309.650000 ;
      RECT 116.500000 308.350000 149.500000 309.650000 ;
      RECT 107.500000 308.350000 108.500000 309.650000 ;
      RECT 66.500000 308.350000 99.500000 309.650000 ;
      RECT 57.500000 308.350000 58.500000 309.650000 ;
      RECT 29.500000 308.350000 49.500000 309.650000 ;
      RECT 15.500000 308.350000 16.500000 309.650000 ;
      RECT 2.020000 308.350000 2.500000 311.170000 ;
      RECT 2.020000 308.070000 16.500000 308.350000 ;
      RECT 1169.500000 308.065000 1183.980000 308.350000 ;
      RECT 1169.500000 307.650000 1186.000000 308.065000 ;
      RECT 1116.500000 307.650000 1156.500000 308.350000 ;
      RECT 1066.500000 307.650000 1108.500000 308.350000 ;
      RECT 1016.500000 307.650000 1058.500000 308.350000 ;
      RECT 966.500000 307.650000 1008.500000 308.350000 ;
      RECT 916.500000 307.650000 958.500000 308.350000 ;
      RECT 866.500000 307.650000 908.500000 308.350000 ;
      RECT 816.500000 307.650000 858.500000 308.350000 ;
      RECT 766.500000 307.650000 808.500000 308.350000 ;
      RECT 716.500000 307.650000 758.500000 308.350000 ;
      RECT 666.500000 307.650000 708.500000 308.350000 ;
      RECT 616.500000 307.650000 658.500000 308.350000 ;
      RECT 566.500000 307.650000 608.500000 308.350000 ;
      RECT 516.500000 307.650000 558.500000 308.350000 ;
      RECT 416.500000 307.650000 508.500000 308.350000 ;
      RECT 366.500000 307.650000 408.500000 308.350000 ;
      RECT 316.500000 307.650000 358.500000 308.350000 ;
      RECT 266.500000 307.650000 308.500000 308.350000 ;
      RECT 216.500000 307.650000 258.500000 308.350000 ;
      RECT 166.500000 307.650000 208.500000 308.350000 ;
      RECT 116.500000 307.650000 158.500000 308.350000 ;
      RECT 66.500000 307.650000 108.500000 308.350000 ;
      RECT 29.500000 307.650000 58.500000 308.350000 ;
      RECT 0.000000 307.650000 16.500000 308.070000 ;
      RECT 1169.500000 306.350000 1170.500000 307.650000 ;
      RECT 1116.500000 306.350000 1149.500000 307.650000 ;
      RECT 1107.500000 306.350000 1108.500000 307.650000 ;
      RECT 1066.500000 306.350000 1099.500000 307.650000 ;
      RECT 1057.500000 306.350000 1058.500000 307.650000 ;
      RECT 1016.500000 306.350000 1049.500000 307.650000 ;
      RECT 1007.500000 306.350000 1008.500000 307.650000 ;
      RECT 966.500000 306.350000 999.500000 307.650000 ;
      RECT 957.500000 306.350000 958.500000 307.650000 ;
      RECT 916.500000 306.350000 949.500000 307.650000 ;
      RECT 907.500000 306.350000 908.500000 307.650000 ;
      RECT 866.500000 306.350000 899.500000 307.650000 ;
      RECT 857.500000 306.350000 858.500000 307.650000 ;
      RECT 816.500000 306.350000 849.500000 307.650000 ;
      RECT 807.500000 306.350000 808.500000 307.650000 ;
      RECT 766.500000 306.350000 799.500000 307.650000 ;
      RECT 757.500000 306.350000 758.500000 307.650000 ;
      RECT 716.500000 306.350000 749.500000 307.650000 ;
      RECT 707.500000 306.350000 708.500000 307.650000 ;
      RECT 666.500000 306.350000 699.500000 307.650000 ;
      RECT 657.500000 306.350000 658.500000 307.650000 ;
      RECT 616.500000 306.350000 649.500000 307.650000 ;
      RECT 607.500000 306.350000 608.500000 307.650000 ;
      RECT 566.500000 306.350000 599.500000 307.650000 ;
      RECT 557.500000 306.350000 558.500000 307.650000 ;
      RECT 516.500000 306.350000 549.500000 307.650000 ;
      RECT 507.500000 306.350000 508.500000 307.650000 ;
      RECT 416.500000 306.350000 499.500000 307.650000 ;
      RECT 407.500000 306.350000 408.500000 307.650000 ;
      RECT 366.500000 306.350000 399.500000 307.650000 ;
      RECT 357.500000 306.350000 358.500000 307.650000 ;
      RECT 316.500000 306.350000 349.500000 307.650000 ;
      RECT 307.500000 306.350000 308.500000 307.650000 ;
      RECT 266.500000 306.350000 299.500000 307.650000 ;
      RECT 257.500000 306.350000 258.500000 307.650000 ;
      RECT 216.500000 306.350000 249.500000 307.650000 ;
      RECT 207.500000 306.350000 208.500000 307.650000 ;
      RECT 166.500000 306.350000 199.500000 307.650000 ;
      RECT 157.500000 306.350000 158.500000 307.650000 ;
      RECT 116.500000 306.350000 149.500000 307.650000 ;
      RECT 107.500000 306.350000 108.500000 307.650000 ;
      RECT 66.500000 306.350000 99.500000 307.650000 ;
      RECT 57.500000 306.350000 58.500000 307.650000 ;
      RECT 29.500000 306.350000 49.500000 307.650000 ;
      RECT 15.500000 306.350000 16.500000 307.650000 ;
      RECT 1157.500000 305.650000 1170.500000 306.350000 ;
      RECT 1107.500000 305.650000 1149.500000 306.350000 ;
      RECT 1057.500000 305.650000 1099.500000 306.350000 ;
      RECT 1007.500000 305.650000 1049.500000 306.350000 ;
      RECT 957.500000 305.650000 999.500000 306.350000 ;
      RECT 907.500000 305.650000 949.500000 306.350000 ;
      RECT 857.500000 305.650000 899.500000 306.350000 ;
      RECT 807.500000 305.650000 849.500000 306.350000 ;
      RECT 757.500000 305.650000 799.500000 306.350000 ;
      RECT 707.500000 305.650000 749.500000 306.350000 ;
      RECT 657.500000 305.650000 699.500000 306.350000 ;
      RECT 607.500000 305.650000 649.500000 306.350000 ;
      RECT 557.500000 305.650000 599.500000 306.350000 ;
      RECT 507.500000 305.650000 549.500000 306.350000 ;
      RECT 407.500000 305.650000 499.500000 306.350000 ;
      RECT 357.500000 305.650000 399.500000 306.350000 ;
      RECT 307.500000 305.650000 349.500000 306.350000 ;
      RECT 257.500000 305.650000 299.500000 306.350000 ;
      RECT 207.500000 305.650000 249.500000 306.350000 ;
      RECT 157.500000 305.650000 199.500000 306.350000 ;
      RECT 107.500000 305.650000 149.500000 306.350000 ;
      RECT 57.500000 305.650000 99.500000 306.350000 ;
      RECT 15.500000 305.650000 49.500000 306.350000 ;
      RECT 1183.500000 305.485000 1186.000000 307.650000 ;
      RECT 1183.500000 304.350000 1183.980000 305.485000 ;
      RECT 1169.500000 304.350000 1170.500000 305.650000 ;
      RECT 1116.500000 304.350000 1149.500000 305.650000 ;
      RECT 1107.500000 304.350000 1108.500000 305.650000 ;
      RECT 1066.500000 304.350000 1099.500000 305.650000 ;
      RECT 1057.500000 304.350000 1058.500000 305.650000 ;
      RECT 1016.500000 304.350000 1049.500000 305.650000 ;
      RECT 1007.500000 304.350000 1008.500000 305.650000 ;
      RECT 966.500000 304.350000 999.500000 305.650000 ;
      RECT 957.500000 304.350000 958.500000 305.650000 ;
      RECT 916.500000 304.350000 949.500000 305.650000 ;
      RECT 907.500000 304.350000 908.500000 305.650000 ;
      RECT 866.500000 304.350000 899.500000 305.650000 ;
      RECT 857.500000 304.350000 858.500000 305.650000 ;
      RECT 816.500000 304.350000 849.500000 305.650000 ;
      RECT 807.500000 304.350000 808.500000 305.650000 ;
      RECT 766.500000 304.350000 799.500000 305.650000 ;
      RECT 757.500000 304.350000 758.500000 305.650000 ;
      RECT 716.500000 304.350000 749.500000 305.650000 ;
      RECT 707.500000 304.350000 708.500000 305.650000 ;
      RECT 666.500000 304.350000 699.500000 305.650000 ;
      RECT 657.500000 304.350000 658.500000 305.650000 ;
      RECT 616.500000 304.350000 649.500000 305.650000 ;
      RECT 607.500000 304.350000 608.500000 305.650000 ;
      RECT 566.500000 304.350000 599.500000 305.650000 ;
      RECT 557.500000 304.350000 558.500000 305.650000 ;
      RECT 516.500000 304.350000 549.500000 305.650000 ;
      RECT 507.500000 304.350000 508.500000 305.650000 ;
      RECT 416.500000 304.350000 499.500000 305.650000 ;
      RECT 407.500000 304.350000 408.500000 305.650000 ;
      RECT 366.500000 304.350000 399.500000 305.650000 ;
      RECT 357.500000 304.350000 358.500000 305.650000 ;
      RECT 316.500000 304.350000 349.500000 305.650000 ;
      RECT 307.500000 304.350000 308.500000 305.650000 ;
      RECT 266.500000 304.350000 299.500000 305.650000 ;
      RECT 257.500000 304.350000 258.500000 305.650000 ;
      RECT 216.500000 304.350000 249.500000 305.650000 ;
      RECT 207.500000 304.350000 208.500000 305.650000 ;
      RECT 166.500000 304.350000 199.500000 305.650000 ;
      RECT 157.500000 304.350000 158.500000 305.650000 ;
      RECT 116.500000 304.350000 149.500000 305.650000 ;
      RECT 107.500000 304.350000 108.500000 305.650000 ;
      RECT 66.500000 304.350000 99.500000 305.650000 ;
      RECT 57.500000 304.350000 58.500000 305.650000 ;
      RECT 29.500000 304.350000 49.500000 305.650000 ;
      RECT 15.500000 304.350000 16.500000 305.650000 ;
      RECT 0.000000 304.350000 2.500000 307.650000 ;
      RECT 1169.500000 303.650000 1183.980000 304.350000 ;
      RECT 1116.500000 303.650000 1156.500000 304.350000 ;
      RECT 1066.500000 303.650000 1108.500000 304.350000 ;
      RECT 1016.500000 303.650000 1058.500000 304.350000 ;
      RECT 966.500000 303.650000 1008.500000 304.350000 ;
      RECT 916.500000 303.650000 958.500000 304.350000 ;
      RECT 866.500000 303.650000 908.500000 304.350000 ;
      RECT 816.500000 303.650000 858.500000 304.350000 ;
      RECT 766.500000 303.650000 808.500000 304.350000 ;
      RECT 716.500000 303.650000 758.500000 304.350000 ;
      RECT 666.500000 303.650000 708.500000 304.350000 ;
      RECT 616.500000 303.650000 658.500000 304.350000 ;
      RECT 566.500000 303.650000 608.500000 304.350000 ;
      RECT 516.500000 303.650000 558.500000 304.350000 ;
      RECT 416.500000 303.650000 508.500000 304.350000 ;
      RECT 366.500000 303.650000 408.500000 304.350000 ;
      RECT 316.500000 303.650000 358.500000 304.350000 ;
      RECT 266.500000 303.650000 308.500000 304.350000 ;
      RECT 216.500000 303.650000 258.500000 304.350000 ;
      RECT 166.500000 303.650000 208.500000 304.350000 ;
      RECT 116.500000 303.650000 158.500000 304.350000 ;
      RECT 66.500000 303.650000 108.500000 304.350000 ;
      RECT 29.500000 303.650000 58.500000 304.350000 ;
      RECT 0.000000 303.650000 16.500000 304.350000 ;
      RECT 1183.500000 302.385000 1183.980000 303.650000 ;
      RECT 1169.500000 302.350000 1170.500000 303.650000 ;
      RECT 1116.500000 302.350000 1149.500000 303.650000 ;
      RECT 1107.500000 302.350000 1108.500000 303.650000 ;
      RECT 1066.500000 302.350000 1099.500000 303.650000 ;
      RECT 1057.500000 302.350000 1058.500000 303.650000 ;
      RECT 1016.500000 302.350000 1049.500000 303.650000 ;
      RECT 1007.500000 302.350000 1008.500000 303.650000 ;
      RECT 966.500000 302.350000 999.500000 303.650000 ;
      RECT 957.500000 302.350000 958.500000 303.650000 ;
      RECT 916.500000 302.350000 949.500000 303.650000 ;
      RECT 907.500000 302.350000 908.500000 303.650000 ;
      RECT 866.500000 302.350000 899.500000 303.650000 ;
      RECT 857.500000 302.350000 858.500000 303.650000 ;
      RECT 816.500000 302.350000 849.500000 303.650000 ;
      RECT 807.500000 302.350000 808.500000 303.650000 ;
      RECT 766.500000 302.350000 799.500000 303.650000 ;
      RECT 757.500000 302.350000 758.500000 303.650000 ;
      RECT 716.500000 302.350000 749.500000 303.650000 ;
      RECT 707.500000 302.350000 708.500000 303.650000 ;
      RECT 666.500000 302.350000 699.500000 303.650000 ;
      RECT 657.500000 302.350000 658.500000 303.650000 ;
      RECT 616.500000 302.350000 649.500000 303.650000 ;
      RECT 607.500000 302.350000 608.500000 303.650000 ;
      RECT 566.500000 302.350000 599.500000 303.650000 ;
      RECT 557.500000 302.350000 558.500000 303.650000 ;
      RECT 516.500000 302.350000 549.500000 303.650000 ;
      RECT 507.500000 302.350000 508.500000 303.650000 ;
      RECT 416.500000 302.350000 499.500000 303.650000 ;
      RECT 407.500000 302.350000 408.500000 303.650000 ;
      RECT 366.500000 302.350000 399.500000 303.650000 ;
      RECT 357.500000 302.350000 358.500000 303.650000 ;
      RECT 316.500000 302.350000 349.500000 303.650000 ;
      RECT 307.500000 302.350000 308.500000 303.650000 ;
      RECT 266.500000 302.350000 299.500000 303.650000 ;
      RECT 257.500000 302.350000 258.500000 303.650000 ;
      RECT 216.500000 302.350000 249.500000 303.650000 ;
      RECT 207.500000 302.350000 208.500000 303.650000 ;
      RECT 166.500000 302.350000 199.500000 303.650000 ;
      RECT 157.500000 302.350000 158.500000 303.650000 ;
      RECT 116.500000 302.350000 149.500000 303.650000 ;
      RECT 107.500000 302.350000 108.500000 303.650000 ;
      RECT 66.500000 302.350000 99.500000 303.650000 ;
      RECT 57.500000 302.350000 58.500000 303.650000 ;
      RECT 29.500000 302.350000 49.500000 303.650000 ;
      RECT 15.500000 302.350000 16.500000 303.650000 ;
      RECT 1157.500000 301.650000 1170.500000 302.350000 ;
      RECT 1107.500000 301.650000 1149.500000 302.350000 ;
      RECT 1057.500000 301.650000 1099.500000 302.350000 ;
      RECT 1007.500000 301.650000 1049.500000 302.350000 ;
      RECT 957.500000 301.650000 999.500000 302.350000 ;
      RECT 907.500000 301.650000 949.500000 302.350000 ;
      RECT 857.500000 301.650000 899.500000 302.350000 ;
      RECT 807.500000 301.650000 849.500000 302.350000 ;
      RECT 757.500000 301.650000 799.500000 302.350000 ;
      RECT 707.500000 301.650000 749.500000 302.350000 ;
      RECT 657.500000 301.650000 699.500000 302.350000 ;
      RECT 607.500000 301.650000 649.500000 302.350000 ;
      RECT 557.500000 301.650000 599.500000 302.350000 ;
      RECT 507.500000 301.650000 549.500000 302.350000 ;
      RECT 407.500000 301.650000 499.500000 302.350000 ;
      RECT 357.500000 301.650000 399.500000 302.350000 ;
      RECT 307.500000 301.650000 349.500000 302.350000 ;
      RECT 257.500000 301.650000 299.500000 302.350000 ;
      RECT 207.500000 301.650000 249.500000 302.350000 ;
      RECT 157.500000 301.650000 199.500000 302.350000 ;
      RECT 107.500000 301.650000 149.500000 302.350000 ;
      RECT 57.500000 301.650000 99.500000 302.350000 ;
      RECT 15.500000 301.650000 49.500000 302.350000 ;
      RECT 1183.500000 301.525000 1186.000000 302.385000 ;
      RECT 0.000000 300.575000 2.500000 303.650000 ;
      RECT 1183.500000 300.350000 1183.980000 301.525000 ;
      RECT 1169.500000 300.350000 1170.500000 301.650000 ;
      RECT 1116.500000 300.350000 1149.500000 301.650000 ;
      RECT 1107.500000 300.350000 1108.500000 301.650000 ;
      RECT 1066.500000 300.350000 1099.500000 301.650000 ;
      RECT 1057.500000 300.350000 1058.500000 301.650000 ;
      RECT 1016.500000 300.350000 1049.500000 301.650000 ;
      RECT 1007.500000 300.350000 1008.500000 301.650000 ;
      RECT 966.500000 300.350000 999.500000 301.650000 ;
      RECT 957.500000 300.350000 958.500000 301.650000 ;
      RECT 916.500000 300.350000 949.500000 301.650000 ;
      RECT 907.500000 300.350000 908.500000 301.650000 ;
      RECT 866.500000 300.350000 899.500000 301.650000 ;
      RECT 857.500000 300.350000 858.500000 301.650000 ;
      RECT 816.500000 300.350000 849.500000 301.650000 ;
      RECT 807.500000 300.350000 808.500000 301.650000 ;
      RECT 766.500000 300.350000 799.500000 301.650000 ;
      RECT 757.500000 300.350000 758.500000 301.650000 ;
      RECT 716.500000 300.350000 749.500000 301.650000 ;
      RECT 707.500000 300.350000 708.500000 301.650000 ;
      RECT 666.500000 300.350000 699.500000 301.650000 ;
      RECT 657.500000 300.350000 658.500000 301.650000 ;
      RECT 616.500000 300.350000 649.500000 301.650000 ;
      RECT 607.500000 300.350000 608.500000 301.650000 ;
      RECT 566.500000 300.350000 599.500000 301.650000 ;
      RECT 557.500000 300.350000 558.500000 301.650000 ;
      RECT 516.500000 300.350000 549.500000 301.650000 ;
      RECT 507.500000 300.350000 508.500000 301.650000 ;
      RECT 416.500000 300.350000 499.500000 301.650000 ;
      RECT 407.500000 300.350000 408.500000 301.650000 ;
      RECT 366.500000 300.350000 399.500000 301.650000 ;
      RECT 357.500000 300.350000 358.500000 301.650000 ;
      RECT 316.500000 300.350000 349.500000 301.650000 ;
      RECT 307.500000 300.350000 308.500000 301.650000 ;
      RECT 266.500000 300.350000 299.500000 301.650000 ;
      RECT 257.500000 300.350000 258.500000 301.650000 ;
      RECT 216.500000 300.350000 249.500000 301.650000 ;
      RECT 207.500000 300.350000 208.500000 301.650000 ;
      RECT 166.500000 300.350000 199.500000 301.650000 ;
      RECT 157.500000 300.350000 158.500000 301.650000 ;
      RECT 116.500000 300.350000 149.500000 301.650000 ;
      RECT 107.500000 300.350000 108.500000 301.650000 ;
      RECT 66.500000 300.350000 99.500000 301.650000 ;
      RECT 57.500000 300.350000 58.500000 301.650000 ;
      RECT 29.500000 300.350000 49.500000 301.650000 ;
      RECT 15.500000 300.350000 16.500000 301.650000 ;
      RECT 2.020000 300.350000 2.500000 300.575000 ;
      RECT 1169.500000 299.650000 1183.980000 300.350000 ;
      RECT 1116.500000 299.650000 1156.500000 300.350000 ;
      RECT 1066.500000 299.650000 1108.500000 300.350000 ;
      RECT 1016.500000 299.650000 1058.500000 300.350000 ;
      RECT 966.500000 299.650000 1008.500000 300.350000 ;
      RECT 916.500000 299.650000 958.500000 300.350000 ;
      RECT 866.500000 299.650000 908.500000 300.350000 ;
      RECT 816.500000 299.650000 858.500000 300.350000 ;
      RECT 766.500000 299.650000 808.500000 300.350000 ;
      RECT 716.500000 299.650000 758.500000 300.350000 ;
      RECT 666.500000 299.650000 708.500000 300.350000 ;
      RECT 616.500000 299.650000 658.500000 300.350000 ;
      RECT 566.500000 299.650000 608.500000 300.350000 ;
      RECT 516.500000 299.650000 558.500000 300.350000 ;
      RECT 416.500000 299.650000 508.500000 300.350000 ;
      RECT 366.500000 299.650000 408.500000 300.350000 ;
      RECT 316.500000 299.650000 358.500000 300.350000 ;
      RECT 266.500000 299.650000 308.500000 300.350000 ;
      RECT 216.500000 299.650000 258.500000 300.350000 ;
      RECT 166.500000 299.650000 208.500000 300.350000 ;
      RECT 116.500000 299.650000 158.500000 300.350000 ;
      RECT 66.500000 299.650000 108.500000 300.350000 ;
      RECT 29.500000 299.650000 58.500000 300.350000 ;
      RECT 2.020000 299.650000 16.500000 300.350000 ;
      RECT 1183.500000 298.425000 1183.980000 299.650000 ;
      RECT 1169.500000 298.350000 1170.500000 299.650000 ;
      RECT 1116.500000 298.350000 1149.500000 299.650000 ;
      RECT 1107.500000 298.350000 1108.500000 299.650000 ;
      RECT 1066.500000 298.350000 1099.500000 299.650000 ;
      RECT 1057.500000 298.350000 1058.500000 299.650000 ;
      RECT 1016.500000 298.350000 1049.500000 299.650000 ;
      RECT 1007.500000 298.350000 1008.500000 299.650000 ;
      RECT 966.500000 298.350000 999.500000 299.650000 ;
      RECT 957.500000 298.350000 958.500000 299.650000 ;
      RECT 916.500000 298.350000 949.500000 299.650000 ;
      RECT 907.500000 298.350000 908.500000 299.650000 ;
      RECT 866.500000 298.350000 899.500000 299.650000 ;
      RECT 857.500000 298.350000 858.500000 299.650000 ;
      RECT 816.500000 298.350000 849.500000 299.650000 ;
      RECT 807.500000 298.350000 808.500000 299.650000 ;
      RECT 766.500000 298.350000 799.500000 299.650000 ;
      RECT 757.500000 298.350000 758.500000 299.650000 ;
      RECT 716.500000 298.350000 749.500000 299.650000 ;
      RECT 707.500000 298.350000 708.500000 299.650000 ;
      RECT 666.500000 298.350000 699.500000 299.650000 ;
      RECT 657.500000 298.350000 658.500000 299.650000 ;
      RECT 616.500000 298.350000 649.500000 299.650000 ;
      RECT 607.500000 298.350000 608.500000 299.650000 ;
      RECT 566.500000 298.350000 599.500000 299.650000 ;
      RECT 557.500000 298.350000 558.500000 299.650000 ;
      RECT 516.500000 298.350000 549.500000 299.650000 ;
      RECT 507.500000 298.350000 508.500000 299.650000 ;
      RECT 416.500000 298.350000 449.500000 299.650000 ;
      RECT 407.500000 298.350000 408.500000 299.650000 ;
      RECT 366.500000 298.350000 399.500000 299.650000 ;
      RECT 357.500000 298.350000 358.500000 299.650000 ;
      RECT 316.500000 298.350000 349.500000 299.650000 ;
      RECT 307.500000 298.350000 308.500000 299.650000 ;
      RECT 266.500000 298.350000 299.500000 299.650000 ;
      RECT 257.500000 298.350000 258.500000 299.650000 ;
      RECT 216.500000 298.350000 249.500000 299.650000 ;
      RECT 207.500000 298.350000 208.500000 299.650000 ;
      RECT 166.500000 298.350000 199.500000 299.650000 ;
      RECT 157.500000 298.350000 158.500000 299.650000 ;
      RECT 116.500000 298.350000 149.500000 299.650000 ;
      RECT 107.500000 298.350000 108.500000 299.650000 ;
      RECT 66.500000 298.350000 99.500000 299.650000 ;
      RECT 57.500000 298.350000 58.500000 299.650000 ;
      RECT 29.500000 298.350000 49.500000 299.650000 ;
      RECT 15.500000 298.350000 16.500000 299.650000 ;
      RECT 1157.500000 297.650000 1170.500000 298.350000 ;
      RECT 1107.500000 297.650000 1149.500000 298.350000 ;
      RECT 1057.500000 297.650000 1099.500000 298.350000 ;
      RECT 1007.500000 297.650000 1049.500000 298.350000 ;
      RECT 957.500000 297.650000 999.500000 298.350000 ;
      RECT 907.500000 297.650000 949.500000 298.350000 ;
      RECT 857.500000 297.650000 899.500000 298.350000 ;
      RECT 807.500000 297.650000 849.500000 298.350000 ;
      RECT 757.500000 297.650000 799.500000 298.350000 ;
      RECT 707.500000 297.650000 749.500000 298.350000 ;
      RECT 657.500000 297.650000 699.500000 298.350000 ;
      RECT 607.500000 297.650000 649.500000 298.350000 ;
      RECT 557.500000 297.650000 599.500000 298.350000 ;
      RECT 507.500000 297.650000 549.500000 298.350000 ;
      RECT 457.500000 297.650000 499.500000 299.650000 ;
      RECT 407.500000 297.650000 449.500000 298.350000 ;
      RECT 357.500000 297.650000 399.500000 298.350000 ;
      RECT 307.500000 297.650000 349.500000 298.350000 ;
      RECT 257.500000 297.650000 299.500000 298.350000 ;
      RECT 207.500000 297.650000 249.500000 298.350000 ;
      RECT 157.500000 297.650000 199.500000 298.350000 ;
      RECT 107.500000 297.650000 149.500000 298.350000 ;
      RECT 57.500000 297.650000 99.500000 298.350000 ;
      RECT 15.500000 297.650000 49.500000 298.350000 ;
      RECT 2.020000 297.475000 2.500000 299.650000 ;
      RECT 0.000000 296.615000 2.500000 297.475000 ;
      RECT 1183.500000 296.350000 1186.000000 298.425000 ;
      RECT 1169.500000 296.350000 1170.500000 297.650000 ;
      RECT 1116.500000 296.350000 1149.500000 297.650000 ;
      RECT 1107.500000 296.350000 1108.500000 297.650000 ;
      RECT 1066.500000 296.350000 1099.500000 297.650000 ;
      RECT 1057.500000 296.350000 1058.500000 297.650000 ;
      RECT 1016.500000 296.350000 1049.500000 297.650000 ;
      RECT 1007.500000 296.350000 1008.500000 297.650000 ;
      RECT 966.500000 296.350000 999.500000 297.650000 ;
      RECT 957.500000 296.350000 958.500000 297.650000 ;
      RECT 916.500000 296.350000 949.500000 297.650000 ;
      RECT 907.500000 296.350000 908.500000 297.650000 ;
      RECT 866.500000 296.350000 899.500000 297.650000 ;
      RECT 857.500000 296.350000 858.500000 297.650000 ;
      RECT 816.500000 296.350000 849.500000 297.650000 ;
      RECT 807.500000 296.350000 808.500000 297.650000 ;
      RECT 766.500000 296.350000 799.500000 297.650000 ;
      RECT 757.500000 296.350000 758.500000 297.650000 ;
      RECT 716.500000 296.350000 749.500000 297.650000 ;
      RECT 707.500000 296.350000 708.500000 297.650000 ;
      RECT 666.500000 296.350000 699.500000 297.650000 ;
      RECT 657.500000 296.350000 658.500000 297.650000 ;
      RECT 616.500000 296.350000 649.500000 297.650000 ;
      RECT 607.500000 296.350000 608.500000 297.650000 ;
      RECT 566.500000 296.350000 599.500000 297.650000 ;
      RECT 557.500000 296.350000 558.500000 297.650000 ;
      RECT 516.500000 296.350000 549.500000 297.650000 ;
      RECT 507.500000 296.350000 508.500000 297.650000 ;
      RECT 466.500000 296.350000 499.500000 297.650000 ;
      RECT 457.500000 296.350000 458.500000 297.650000 ;
      RECT 416.500000 296.350000 449.500000 297.650000 ;
      RECT 407.500000 296.350000 408.500000 297.650000 ;
      RECT 366.500000 296.350000 399.500000 297.650000 ;
      RECT 357.500000 296.350000 358.500000 297.650000 ;
      RECT 316.500000 296.350000 349.500000 297.650000 ;
      RECT 307.500000 296.350000 308.500000 297.650000 ;
      RECT 266.500000 296.350000 299.500000 297.650000 ;
      RECT 257.500000 296.350000 258.500000 297.650000 ;
      RECT 216.500000 296.350000 249.500000 297.650000 ;
      RECT 207.500000 296.350000 208.500000 297.650000 ;
      RECT 166.500000 296.350000 199.500000 297.650000 ;
      RECT 157.500000 296.350000 158.500000 297.650000 ;
      RECT 116.500000 296.350000 149.500000 297.650000 ;
      RECT 107.500000 296.350000 108.500000 297.650000 ;
      RECT 66.500000 296.350000 99.500000 297.650000 ;
      RECT 57.500000 296.350000 58.500000 297.650000 ;
      RECT 29.500000 296.350000 49.500000 297.650000 ;
      RECT 15.500000 296.350000 16.500000 297.650000 ;
      RECT 2.020000 296.350000 2.500000 296.615000 ;
      RECT 1169.500000 295.650000 1186.000000 296.350000 ;
      RECT 1116.500000 295.650000 1156.500000 296.350000 ;
      RECT 1066.500000 295.650000 1108.500000 296.350000 ;
      RECT 1016.500000 295.650000 1058.500000 296.350000 ;
      RECT 966.500000 295.650000 1008.500000 296.350000 ;
      RECT 916.500000 295.650000 958.500000 296.350000 ;
      RECT 866.500000 295.650000 908.500000 296.350000 ;
      RECT 816.500000 295.650000 858.500000 296.350000 ;
      RECT 766.500000 295.650000 808.500000 296.350000 ;
      RECT 716.500000 295.650000 758.500000 296.350000 ;
      RECT 666.500000 295.650000 708.500000 296.350000 ;
      RECT 616.500000 295.650000 658.500000 296.350000 ;
      RECT 566.500000 295.650000 608.500000 296.350000 ;
      RECT 516.500000 295.650000 558.500000 296.350000 ;
      RECT 466.500000 295.650000 508.500000 296.350000 ;
      RECT 416.500000 295.650000 458.500000 296.350000 ;
      RECT 366.500000 295.650000 408.500000 296.350000 ;
      RECT 316.500000 295.650000 358.500000 296.350000 ;
      RECT 266.500000 295.650000 308.500000 296.350000 ;
      RECT 216.500000 295.650000 258.500000 296.350000 ;
      RECT 166.500000 295.650000 208.500000 296.350000 ;
      RECT 116.500000 295.650000 158.500000 296.350000 ;
      RECT 66.500000 295.650000 108.500000 296.350000 ;
      RECT 29.500000 295.650000 58.500000 296.350000 ;
      RECT 2.020000 295.650000 16.500000 296.350000 ;
      RECT 1169.500000 294.350000 1170.500000 295.650000 ;
      RECT 1116.500000 294.350000 1149.500000 295.650000 ;
      RECT 1107.500000 294.350000 1108.500000 295.650000 ;
      RECT 1066.500000 294.350000 1099.500000 295.650000 ;
      RECT 1057.500000 294.350000 1058.500000 295.650000 ;
      RECT 1016.500000 294.350000 1049.500000 295.650000 ;
      RECT 1007.500000 294.350000 1008.500000 295.650000 ;
      RECT 966.500000 294.350000 999.500000 295.650000 ;
      RECT 957.500000 294.350000 958.500000 295.650000 ;
      RECT 916.500000 294.350000 949.500000 295.650000 ;
      RECT 907.500000 294.350000 908.500000 295.650000 ;
      RECT 866.500000 294.350000 899.500000 295.650000 ;
      RECT 857.500000 294.350000 858.500000 295.650000 ;
      RECT 816.500000 294.350000 849.500000 295.650000 ;
      RECT 807.500000 294.350000 808.500000 295.650000 ;
      RECT 766.500000 294.350000 799.500000 295.650000 ;
      RECT 757.500000 294.350000 758.500000 295.650000 ;
      RECT 716.500000 294.350000 749.500000 295.650000 ;
      RECT 707.500000 294.350000 708.500000 295.650000 ;
      RECT 666.500000 294.350000 699.500000 295.650000 ;
      RECT 657.500000 294.350000 658.500000 295.650000 ;
      RECT 616.500000 294.350000 649.500000 295.650000 ;
      RECT 607.500000 294.350000 608.500000 295.650000 ;
      RECT 566.500000 294.350000 599.500000 295.650000 ;
      RECT 557.500000 294.350000 558.500000 295.650000 ;
      RECT 516.500000 294.350000 549.500000 295.650000 ;
      RECT 507.500000 294.350000 508.500000 295.650000 ;
      RECT 466.500000 294.350000 499.500000 295.650000 ;
      RECT 457.500000 294.350000 458.500000 295.650000 ;
      RECT 416.500000 294.350000 449.500000 295.650000 ;
      RECT 407.500000 294.350000 408.500000 295.650000 ;
      RECT 366.500000 294.350000 399.500000 295.650000 ;
      RECT 357.500000 294.350000 358.500000 295.650000 ;
      RECT 316.500000 294.350000 349.500000 295.650000 ;
      RECT 307.500000 294.350000 308.500000 295.650000 ;
      RECT 266.500000 294.350000 299.500000 295.650000 ;
      RECT 257.500000 294.350000 258.500000 295.650000 ;
      RECT 216.500000 294.350000 249.500000 295.650000 ;
      RECT 207.500000 294.350000 208.500000 295.650000 ;
      RECT 166.500000 294.350000 199.500000 295.650000 ;
      RECT 157.500000 294.350000 158.500000 295.650000 ;
      RECT 116.500000 294.350000 149.500000 295.650000 ;
      RECT 107.500000 294.350000 108.500000 295.650000 ;
      RECT 66.500000 294.350000 99.500000 295.650000 ;
      RECT 57.500000 294.350000 58.500000 295.650000 ;
      RECT 29.500000 294.350000 49.500000 295.650000 ;
      RECT 15.500000 294.350000 16.500000 295.650000 ;
      RECT 1157.500000 293.650000 1170.500000 294.350000 ;
      RECT 1107.500000 293.650000 1149.500000 294.350000 ;
      RECT 1057.500000 293.650000 1099.500000 294.350000 ;
      RECT 1007.500000 293.650000 1049.500000 294.350000 ;
      RECT 957.500000 293.650000 999.500000 294.350000 ;
      RECT 907.500000 293.650000 949.500000 294.350000 ;
      RECT 857.500000 293.650000 899.500000 294.350000 ;
      RECT 807.500000 293.650000 849.500000 294.350000 ;
      RECT 757.500000 293.650000 799.500000 294.350000 ;
      RECT 707.500000 293.650000 749.500000 294.350000 ;
      RECT 657.500000 293.650000 699.500000 294.350000 ;
      RECT 607.500000 293.650000 649.500000 294.350000 ;
      RECT 557.500000 293.650000 599.500000 294.350000 ;
      RECT 507.500000 293.650000 549.500000 294.350000 ;
      RECT 457.500000 293.650000 499.500000 294.350000 ;
      RECT 407.500000 293.650000 449.500000 294.350000 ;
      RECT 357.500000 293.650000 399.500000 294.350000 ;
      RECT 307.500000 293.650000 349.500000 294.350000 ;
      RECT 257.500000 293.650000 299.500000 294.350000 ;
      RECT 207.500000 293.650000 249.500000 294.350000 ;
      RECT 157.500000 293.650000 199.500000 294.350000 ;
      RECT 107.500000 293.650000 149.500000 294.350000 ;
      RECT 57.500000 293.650000 99.500000 294.350000 ;
      RECT 15.500000 293.650000 49.500000 294.350000 ;
      RECT 2.020000 293.515000 2.500000 295.650000 ;
      RECT 1183.500000 292.350000 1186.000000 295.650000 ;
      RECT 1169.500000 292.350000 1170.500000 293.650000 ;
      RECT 1116.500000 292.350000 1149.500000 293.650000 ;
      RECT 1107.500000 292.350000 1108.500000 293.650000 ;
      RECT 1066.500000 292.350000 1099.500000 293.650000 ;
      RECT 1057.500000 292.350000 1058.500000 293.650000 ;
      RECT 1016.500000 292.350000 1049.500000 293.650000 ;
      RECT 1007.500000 292.350000 1008.500000 293.650000 ;
      RECT 966.500000 292.350000 999.500000 293.650000 ;
      RECT 957.500000 292.350000 958.500000 293.650000 ;
      RECT 916.500000 292.350000 949.500000 293.650000 ;
      RECT 907.500000 292.350000 908.500000 293.650000 ;
      RECT 866.500000 292.350000 899.500000 293.650000 ;
      RECT 857.500000 292.350000 858.500000 293.650000 ;
      RECT 816.500000 292.350000 849.500000 293.650000 ;
      RECT 807.500000 292.350000 808.500000 293.650000 ;
      RECT 766.500000 292.350000 799.500000 293.650000 ;
      RECT 757.500000 292.350000 758.500000 293.650000 ;
      RECT 716.500000 292.350000 749.500000 293.650000 ;
      RECT 707.500000 292.350000 708.500000 293.650000 ;
      RECT 666.500000 292.350000 699.500000 293.650000 ;
      RECT 657.500000 292.350000 658.500000 293.650000 ;
      RECT 616.500000 292.350000 649.500000 293.650000 ;
      RECT 607.500000 292.350000 608.500000 293.650000 ;
      RECT 566.500000 292.350000 599.500000 293.650000 ;
      RECT 557.500000 292.350000 558.500000 293.650000 ;
      RECT 516.500000 292.350000 549.500000 293.650000 ;
      RECT 507.500000 292.350000 508.500000 293.650000 ;
      RECT 466.500000 292.350000 499.500000 293.650000 ;
      RECT 457.500000 292.350000 458.500000 293.650000 ;
      RECT 416.500000 292.350000 449.500000 293.650000 ;
      RECT 407.500000 292.350000 408.500000 293.650000 ;
      RECT 366.500000 292.350000 399.500000 293.650000 ;
      RECT 357.500000 292.350000 358.500000 293.650000 ;
      RECT 316.500000 292.350000 349.500000 293.650000 ;
      RECT 307.500000 292.350000 308.500000 293.650000 ;
      RECT 266.500000 292.350000 299.500000 293.650000 ;
      RECT 257.500000 292.350000 258.500000 293.650000 ;
      RECT 216.500000 292.350000 249.500000 293.650000 ;
      RECT 207.500000 292.350000 208.500000 293.650000 ;
      RECT 166.500000 292.350000 199.500000 293.650000 ;
      RECT 157.500000 292.350000 158.500000 293.650000 ;
      RECT 116.500000 292.350000 149.500000 293.650000 ;
      RECT 107.500000 292.350000 108.500000 293.650000 ;
      RECT 66.500000 292.350000 99.500000 293.650000 ;
      RECT 57.500000 292.350000 58.500000 293.650000 ;
      RECT 29.500000 292.350000 49.500000 293.650000 ;
      RECT 15.500000 292.350000 16.500000 293.650000 ;
      RECT 0.000000 292.350000 2.500000 293.515000 ;
      RECT 1169.500000 291.650000 1186.000000 292.350000 ;
      RECT 1116.500000 291.650000 1156.500000 292.350000 ;
      RECT 1066.500000 291.650000 1108.500000 292.350000 ;
      RECT 1016.500000 291.650000 1058.500000 292.350000 ;
      RECT 966.500000 291.650000 1008.500000 292.350000 ;
      RECT 916.500000 291.650000 958.500000 292.350000 ;
      RECT 866.500000 291.650000 908.500000 292.350000 ;
      RECT 816.500000 291.650000 858.500000 292.350000 ;
      RECT 766.500000 291.650000 808.500000 292.350000 ;
      RECT 716.500000 291.650000 758.500000 292.350000 ;
      RECT 666.500000 291.650000 708.500000 292.350000 ;
      RECT 616.500000 291.650000 658.500000 292.350000 ;
      RECT 566.500000 291.650000 608.500000 292.350000 ;
      RECT 516.500000 291.650000 558.500000 292.350000 ;
      RECT 466.500000 291.650000 508.500000 292.350000 ;
      RECT 416.500000 291.650000 458.500000 292.350000 ;
      RECT 366.500000 291.650000 408.500000 292.350000 ;
      RECT 316.500000 291.650000 358.500000 292.350000 ;
      RECT 266.500000 291.650000 308.500000 292.350000 ;
      RECT 216.500000 291.650000 258.500000 292.350000 ;
      RECT 166.500000 291.650000 208.500000 292.350000 ;
      RECT 116.500000 291.650000 158.500000 292.350000 ;
      RECT 66.500000 291.650000 108.500000 292.350000 ;
      RECT 29.500000 291.650000 58.500000 292.350000 ;
      RECT 0.000000 291.650000 16.500000 292.350000 ;
      RECT 0.000000 290.935000 2.500000 291.650000 ;
      RECT 1183.500000 290.930000 1186.000000 291.650000 ;
      RECT 1169.500000 290.350000 1170.500000 291.650000 ;
      RECT 1116.500000 290.350000 1149.500000 291.650000 ;
      RECT 1107.500000 290.350000 1108.500000 291.650000 ;
      RECT 1066.500000 290.350000 1099.500000 291.650000 ;
      RECT 1057.500000 290.350000 1058.500000 291.650000 ;
      RECT 1016.500000 290.350000 1049.500000 291.650000 ;
      RECT 1007.500000 290.350000 1008.500000 291.650000 ;
      RECT 966.500000 290.350000 999.500000 291.650000 ;
      RECT 957.500000 290.350000 958.500000 291.650000 ;
      RECT 916.500000 290.350000 949.500000 291.650000 ;
      RECT 907.500000 290.350000 908.500000 291.650000 ;
      RECT 866.500000 290.350000 899.500000 291.650000 ;
      RECT 857.500000 290.350000 858.500000 291.650000 ;
      RECT 816.500000 290.350000 849.500000 291.650000 ;
      RECT 807.500000 290.350000 808.500000 291.650000 ;
      RECT 766.500000 290.350000 799.500000 291.650000 ;
      RECT 757.500000 290.350000 758.500000 291.650000 ;
      RECT 716.500000 290.350000 749.500000 291.650000 ;
      RECT 707.500000 290.350000 708.500000 291.650000 ;
      RECT 666.500000 290.350000 699.500000 291.650000 ;
      RECT 657.500000 290.350000 658.500000 291.650000 ;
      RECT 616.500000 290.350000 649.500000 291.650000 ;
      RECT 607.500000 290.350000 608.500000 291.650000 ;
      RECT 566.500000 290.350000 599.500000 291.650000 ;
      RECT 557.500000 290.350000 558.500000 291.650000 ;
      RECT 516.500000 290.350000 549.500000 291.650000 ;
      RECT 507.500000 290.350000 508.500000 291.650000 ;
      RECT 466.500000 290.350000 499.500000 291.650000 ;
      RECT 457.500000 290.350000 458.500000 291.650000 ;
      RECT 416.500000 290.350000 449.500000 291.650000 ;
      RECT 407.500000 290.350000 408.500000 291.650000 ;
      RECT 366.500000 290.350000 399.500000 291.650000 ;
      RECT 357.500000 290.350000 358.500000 291.650000 ;
      RECT 316.500000 290.350000 349.500000 291.650000 ;
      RECT 307.500000 290.350000 308.500000 291.650000 ;
      RECT 266.500000 290.350000 299.500000 291.650000 ;
      RECT 257.500000 290.350000 258.500000 291.650000 ;
      RECT 216.500000 290.350000 249.500000 291.650000 ;
      RECT 207.500000 290.350000 208.500000 291.650000 ;
      RECT 166.500000 290.350000 199.500000 291.650000 ;
      RECT 157.500000 290.350000 158.500000 291.650000 ;
      RECT 116.500000 290.350000 149.500000 291.650000 ;
      RECT 107.500000 290.350000 108.500000 291.650000 ;
      RECT 66.500000 290.350000 99.500000 291.650000 ;
      RECT 57.500000 290.350000 58.500000 291.650000 ;
      RECT 29.500000 290.350000 49.500000 291.650000 ;
      RECT 15.500000 290.350000 16.500000 291.650000 ;
      RECT 1157.500000 289.650000 1170.500000 290.350000 ;
      RECT 1107.500000 289.650000 1149.500000 290.350000 ;
      RECT 1057.500000 289.650000 1099.500000 290.350000 ;
      RECT 1007.500000 289.650000 1049.500000 290.350000 ;
      RECT 957.500000 289.650000 999.500000 290.350000 ;
      RECT 907.500000 289.650000 949.500000 290.350000 ;
      RECT 857.500000 289.650000 899.500000 290.350000 ;
      RECT 807.500000 289.650000 849.500000 290.350000 ;
      RECT 757.500000 289.650000 799.500000 290.350000 ;
      RECT 707.500000 289.650000 749.500000 290.350000 ;
      RECT 657.500000 289.650000 699.500000 290.350000 ;
      RECT 607.500000 289.650000 649.500000 290.350000 ;
      RECT 557.500000 289.650000 599.500000 290.350000 ;
      RECT 507.500000 289.650000 549.500000 290.350000 ;
      RECT 457.500000 289.650000 499.500000 290.350000 ;
      RECT 407.500000 289.650000 449.500000 290.350000 ;
      RECT 357.500000 289.650000 399.500000 290.350000 ;
      RECT 307.500000 289.650000 349.500000 290.350000 ;
      RECT 257.500000 289.650000 299.500000 290.350000 ;
      RECT 207.500000 289.650000 249.500000 290.350000 ;
      RECT 157.500000 289.650000 199.500000 290.350000 ;
      RECT 107.500000 289.650000 149.500000 290.350000 ;
      RECT 57.500000 289.650000 99.500000 290.350000 ;
      RECT 15.500000 289.650000 49.500000 290.350000 ;
      RECT 1183.500000 288.350000 1183.980000 290.930000 ;
      RECT 1169.500000 288.350000 1170.500000 289.650000 ;
      RECT 1116.500000 288.350000 1149.500000 289.650000 ;
      RECT 1107.500000 288.350000 1108.500000 289.650000 ;
      RECT 1066.500000 288.350000 1099.500000 289.650000 ;
      RECT 1057.500000 288.350000 1058.500000 289.650000 ;
      RECT 1016.500000 288.350000 1049.500000 289.650000 ;
      RECT 1007.500000 288.350000 1008.500000 289.650000 ;
      RECT 966.500000 288.350000 999.500000 289.650000 ;
      RECT 957.500000 288.350000 958.500000 289.650000 ;
      RECT 916.500000 288.350000 949.500000 289.650000 ;
      RECT 907.500000 288.350000 908.500000 289.650000 ;
      RECT 866.500000 288.350000 899.500000 289.650000 ;
      RECT 857.500000 288.350000 858.500000 289.650000 ;
      RECT 816.500000 288.350000 849.500000 289.650000 ;
      RECT 807.500000 288.350000 808.500000 289.650000 ;
      RECT 766.500000 288.350000 799.500000 289.650000 ;
      RECT 757.500000 288.350000 758.500000 289.650000 ;
      RECT 716.500000 288.350000 749.500000 289.650000 ;
      RECT 707.500000 288.350000 708.500000 289.650000 ;
      RECT 666.500000 288.350000 699.500000 289.650000 ;
      RECT 657.500000 288.350000 658.500000 289.650000 ;
      RECT 616.500000 288.350000 649.500000 289.650000 ;
      RECT 607.500000 288.350000 608.500000 289.650000 ;
      RECT 566.500000 288.350000 599.500000 289.650000 ;
      RECT 557.500000 288.350000 558.500000 289.650000 ;
      RECT 516.500000 288.350000 549.500000 289.650000 ;
      RECT 507.500000 288.350000 508.500000 289.650000 ;
      RECT 466.500000 288.350000 499.500000 289.650000 ;
      RECT 457.500000 288.350000 458.500000 289.650000 ;
      RECT 416.500000 288.350000 449.500000 289.650000 ;
      RECT 407.500000 288.350000 408.500000 289.650000 ;
      RECT 366.500000 288.350000 399.500000 289.650000 ;
      RECT 357.500000 288.350000 358.500000 289.650000 ;
      RECT 316.500000 288.350000 349.500000 289.650000 ;
      RECT 307.500000 288.350000 308.500000 289.650000 ;
      RECT 266.500000 288.350000 299.500000 289.650000 ;
      RECT 257.500000 288.350000 258.500000 289.650000 ;
      RECT 216.500000 288.350000 249.500000 289.650000 ;
      RECT 207.500000 288.350000 208.500000 289.650000 ;
      RECT 166.500000 288.350000 199.500000 289.650000 ;
      RECT 157.500000 288.350000 158.500000 289.650000 ;
      RECT 116.500000 288.350000 149.500000 289.650000 ;
      RECT 107.500000 288.350000 108.500000 289.650000 ;
      RECT 66.500000 288.350000 99.500000 289.650000 ;
      RECT 57.500000 288.350000 58.500000 289.650000 ;
      RECT 29.500000 288.350000 49.500000 289.650000 ;
      RECT 15.500000 288.350000 16.500000 289.650000 ;
      RECT 2.020000 288.350000 2.500000 290.935000 ;
      RECT 2.020000 287.835000 16.500000 288.350000 ;
      RECT 1169.500000 287.830000 1183.980000 288.350000 ;
      RECT 1169.500000 287.650000 1186.000000 287.830000 ;
      RECT 1116.500000 287.650000 1156.500000 288.350000 ;
      RECT 1066.500000 287.650000 1108.500000 288.350000 ;
      RECT 1016.500000 287.650000 1058.500000 288.350000 ;
      RECT 966.500000 287.650000 1008.500000 288.350000 ;
      RECT 916.500000 287.650000 958.500000 288.350000 ;
      RECT 866.500000 287.650000 908.500000 288.350000 ;
      RECT 816.500000 287.650000 858.500000 288.350000 ;
      RECT 766.500000 287.650000 808.500000 288.350000 ;
      RECT 716.500000 287.650000 758.500000 288.350000 ;
      RECT 666.500000 287.650000 708.500000 288.350000 ;
      RECT 616.500000 287.650000 658.500000 288.350000 ;
      RECT 566.500000 287.650000 608.500000 288.350000 ;
      RECT 516.500000 287.650000 558.500000 288.350000 ;
      RECT 466.500000 287.650000 508.500000 288.350000 ;
      RECT 416.500000 287.650000 458.500000 288.350000 ;
      RECT 366.500000 287.650000 408.500000 288.350000 ;
      RECT 316.500000 287.650000 358.500000 288.350000 ;
      RECT 266.500000 287.650000 308.500000 288.350000 ;
      RECT 216.500000 287.650000 258.500000 288.350000 ;
      RECT 166.500000 287.650000 208.500000 288.350000 ;
      RECT 116.500000 287.650000 158.500000 288.350000 ;
      RECT 66.500000 287.650000 108.500000 288.350000 ;
      RECT 29.500000 287.650000 58.500000 288.350000 ;
      RECT 0.000000 287.650000 16.500000 287.835000 ;
      RECT 1169.500000 286.350000 1170.500000 287.650000 ;
      RECT 1116.500000 286.350000 1149.500000 287.650000 ;
      RECT 1107.500000 286.350000 1108.500000 287.650000 ;
      RECT 1066.500000 286.350000 1099.500000 287.650000 ;
      RECT 1057.500000 286.350000 1058.500000 287.650000 ;
      RECT 1016.500000 286.350000 1049.500000 287.650000 ;
      RECT 1007.500000 286.350000 1008.500000 287.650000 ;
      RECT 966.500000 286.350000 999.500000 287.650000 ;
      RECT 957.500000 286.350000 958.500000 287.650000 ;
      RECT 916.500000 286.350000 949.500000 287.650000 ;
      RECT 907.500000 286.350000 908.500000 287.650000 ;
      RECT 866.500000 286.350000 899.500000 287.650000 ;
      RECT 857.500000 286.350000 858.500000 287.650000 ;
      RECT 816.500000 286.350000 849.500000 287.650000 ;
      RECT 807.500000 286.350000 808.500000 287.650000 ;
      RECT 766.500000 286.350000 799.500000 287.650000 ;
      RECT 757.500000 286.350000 758.500000 287.650000 ;
      RECT 716.500000 286.350000 749.500000 287.650000 ;
      RECT 707.500000 286.350000 708.500000 287.650000 ;
      RECT 666.500000 286.350000 699.500000 287.650000 ;
      RECT 657.500000 286.350000 658.500000 287.650000 ;
      RECT 616.500000 286.350000 649.500000 287.650000 ;
      RECT 607.500000 286.350000 608.500000 287.650000 ;
      RECT 566.500000 286.350000 599.500000 287.650000 ;
      RECT 557.500000 286.350000 558.500000 287.650000 ;
      RECT 516.500000 286.350000 549.500000 287.650000 ;
      RECT 507.500000 286.350000 508.500000 287.650000 ;
      RECT 466.500000 286.350000 499.500000 287.650000 ;
      RECT 457.500000 286.350000 458.500000 287.650000 ;
      RECT 416.500000 286.350000 449.500000 287.650000 ;
      RECT 407.500000 286.350000 408.500000 287.650000 ;
      RECT 366.500000 286.350000 399.500000 287.650000 ;
      RECT 357.500000 286.350000 358.500000 287.650000 ;
      RECT 316.500000 286.350000 349.500000 287.650000 ;
      RECT 307.500000 286.350000 308.500000 287.650000 ;
      RECT 266.500000 286.350000 299.500000 287.650000 ;
      RECT 257.500000 286.350000 258.500000 287.650000 ;
      RECT 216.500000 286.350000 249.500000 287.650000 ;
      RECT 207.500000 286.350000 208.500000 287.650000 ;
      RECT 166.500000 286.350000 199.500000 287.650000 ;
      RECT 157.500000 286.350000 158.500000 287.650000 ;
      RECT 116.500000 286.350000 149.500000 287.650000 ;
      RECT 107.500000 286.350000 108.500000 287.650000 ;
      RECT 66.500000 286.350000 99.500000 287.650000 ;
      RECT 57.500000 286.350000 58.500000 287.650000 ;
      RECT 29.500000 286.350000 49.500000 287.650000 ;
      RECT 15.500000 286.350000 16.500000 287.650000 ;
      RECT 1157.500000 285.650000 1170.500000 286.350000 ;
      RECT 1107.500000 285.650000 1149.500000 286.350000 ;
      RECT 1057.500000 285.650000 1099.500000 286.350000 ;
      RECT 1007.500000 285.650000 1049.500000 286.350000 ;
      RECT 957.500000 285.650000 999.500000 286.350000 ;
      RECT 907.500000 285.650000 949.500000 286.350000 ;
      RECT 857.500000 285.650000 899.500000 286.350000 ;
      RECT 807.500000 285.650000 849.500000 286.350000 ;
      RECT 757.500000 285.650000 799.500000 286.350000 ;
      RECT 707.500000 285.650000 749.500000 286.350000 ;
      RECT 657.500000 285.650000 699.500000 286.350000 ;
      RECT 607.500000 285.650000 649.500000 286.350000 ;
      RECT 557.500000 285.650000 599.500000 286.350000 ;
      RECT 507.500000 285.650000 549.500000 286.350000 ;
      RECT 457.500000 285.650000 499.500000 286.350000 ;
      RECT 407.500000 285.650000 449.500000 286.350000 ;
      RECT 357.500000 285.650000 399.500000 286.350000 ;
      RECT 307.500000 285.650000 349.500000 286.350000 ;
      RECT 257.500000 285.650000 299.500000 286.350000 ;
      RECT 207.500000 285.650000 249.500000 286.350000 ;
      RECT 157.500000 285.650000 199.500000 286.350000 ;
      RECT 107.500000 285.650000 149.500000 286.350000 ;
      RECT 57.500000 285.650000 99.500000 286.350000 ;
      RECT 15.500000 285.650000 49.500000 286.350000 ;
      RECT 1183.500000 284.350000 1186.000000 287.650000 ;
      RECT 1169.500000 284.350000 1170.500000 285.650000 ;
      RECT 1116.500000 284.350000 1149.500000 285.650000 ;
      RECT 1107.500000 284.350000 1108.500000 285.650000 ;
      RECT 1066.500000 284.350000 1099.500000 285.650000 ;
      RECT 1057.500000 284.350000 1058.500000 285.650000 ;
      RECT 1016.500000 284.350000 1049.500000 285.650000 ;
      RECT 1007.500000 284.350000 1008.500000 285.650000 ;
      RECT 966.500000 284.350000 999.500000 285.650000 ;
      RECT 957.500000 284.350000 958.500000 285.650000 ;
      RECT 916.500000 284.350000 949.500000 285.650000 ;
      RECT 907.500000 284.350000 908.500000 285.650000 ;
      RECT 866.500000 284.350000 899.500000 285.650000 ;
      RECT 857.500000 284.350000 858.500000 285.650000 ;
      RECT 816.500000 284.350000 849.500000 285.650000 ;
      RECT 807.500000 284.350000 808.500000 285.650000 ;
      RECT 766.500000 284.350000 799.500000 285.650000 ;
      RECT 757.500000 284.350000 758.500000 285.650000 ;
      RECT 716.500000 284.350000 749.500000 285.650000 ;
      RECT 707.500000 284.350000 708.500000 285.650000 ;
      RECT 666.500000 284.350000 699.500000 285.650000 ;
      RECT 657.500000 284.350000 658.500000 285.650000 ;
      RECT 616.500000 284.350000 649.500000 285.650000 ;
      RECT 607.500000 284.350000 608.500000 285.650000 ;
      RECT 566.500000 284.350000 599.500000 285.650000 ;
      RECT 557.500000 284.350000 558.500000 285.650000 ;
      RECT 516.500000 284.350000 549.500000 285.650000 ;
      RECT 507.500000 284.350000 508.500000 285.650000 ;
      RECT 466.500000 284.350000 499.500000 285.650000 ;
      RECT 457.500000 284.350000 458.500000 285.650000 ;
      RECT 416.500000 284.350000 449.500000 285.650000 ;
      RECT 407.500000 284.350000 408.500000 285.650000 ;
      RECT 366.500000 284.350000 399.500000 285.650000 ;
      RECT 357.500000 284.350000 358.500000 285.650000 ;
      RECT 316.500000 284.350000 349.500000 285.650000 ;
      RECT 307.500000 284.350000 308.500000 285.650000 ;
      RECT 266.500000 284.350000 299.500000 285.650000 ;
      RECT 257.500000 284.350000 258.500000 285.650000 ;
      RECT 216.500000 284.350000 249.500000 285.650000 ;
      RECT 207.500000 284.350000 208.500000 285.650000 ;
      RECT 166.500000 284.350000 199.500000 285.650000 ;
      RECT 157.500000 284.350000 158.500000 285.650000 ;
      RECT 116.500000 284.350000 149.500000 285.650000 ;
      RECT 107.500000 284.350000 108.500000 285.650000 ;
      RECT 66.500000 284.350000 99.500000 285.650000 ;
      RECT 57.500000 284.350000 58.500000 285.650000 ;
      RECT 29.500000 284.350000 49.500000 285.650000 ;
      RECT 15.500000 284.350000 16.500000 285.650000 ;
      RECT 0.000000 284.350000 2.500000 287.650000 ;
      RECT 1169.500000 283.650000 1186.000000 284.350000 ;
      RECT 1116.500000 283.650000 1156.500000 284.350000 ;
      RECT 1066.500000 283.650000 1108.500000 284.350000 ;
      RECT 1016.500000 283.650000 1058.500000 284.350000 ;
      RECT 966.500000 283.650000 1008.500000 284.350000 ;
      RECT 916.500000 283.650000 958.500000 284.350000 ;
      RECT 866.500000 283.650000 908.500000 284.350000 ;
      RECT 816.500000 283.650000 858.500000 284.350000 ;
      RECT 766.500000 283.650000 808.500000 284.350000 ;
      RECT 716.500000 283.650000 758.500000 284.350000 ;
      RECT 666.500000 283.650000 708.500000 284.350000 ;
      RECT 616.500000 283.650000 658.500000 284.350000 ;
      RECT 566.500000 283.650000 608.500000 284.350000 ;
      RECT 516.500000 283.650000 558.500000 284.350000 ;
      RECT 466.500000 283.650000 508.500000 284.350000 ;
      RECT 416.500000 283.650000 458.500000 284.350000 ;
      RECT 366.500000 283.650000 408.500000 284.350000 ;
      RECT 316.500000 283.650000 358.500000 284.350000 ;
      RECT 266.500000 283.650000 308.500000 284.350000 ;
      RECT 216.500000 283.650000 258.500000 284.350000 ;
      RECT 166.500000 283.650000 208.500000 284.350000 ;
      RECT 116.500000 283.650000 158.500000 284.350000 ;
      RECT 66.500000 283.650000 108.500000 284.350000 ;
      RECT 29.500000 283.650000 58.500000 284.350000 ;
      RECT 0.000000 283.650000 16.500000 284.350000 ;
      RECT 1169.500000 282.350000 1170.500000 283.650000 ;
      RECT 1116.500000 282.350000 1149.500000 283.650000 ;
      RECT 1107.500000 282.350000 1108.500000 283.650000 ;
      RECT 1066.500000 282.350000 1099.500000 283.650000 ;
      RECT 1057.500000 282.350000 1058.500000 283.650000 ;
      RECT 1016.500000 282.350000 1049.500000 283.650000 ;
      RECT 1007.500000 282.350000 1008.500000 283.650000 ;
      RECT 966.500000 282.350000 999.500000 283.650000 ;
      RECT 957.500000 282.350000 958.500000 283.650000 ;
      RECT 916.500000 282.350000 949.500000 283.650000 ;
      RECT 907.500000 282.350000 908.500000 283.650000 ;
      RECT 866.500000 282.350000 899.500000 283.650000 ;
      RECT 857.500000 282.350000 858.500000 283.650000 ;
      RECT 816.500000 282.350000 849.500000 283.650000 ;
      RECT 807.500000 282.350000 808.500000 283.650000 ;
      RECT 766.500000 282.350000 799.500000 283.650000 ;
      RECT 757.500000 282.350000 758.500000 283.650000 ;
      RECT 716.500000 282.350000 749.500000 283.650000 ;
      RECT 707.500000 282.350000 708.500000 283.650000 ;
      RECT 666.500000 282.350000 699.500000 283.650000 ;
      RECT 657.500000 282.350000 658.500000 283.650000 ;
      RECT 616.500000 282.350000 649.500000 283.650000 ;
      RECT 607.500000 282.350000 608.500000 283.650000 ;
      RECT 566.500000 282.350000 599.500000 283.650000 ;
      RECT 557.500000 282.350000 558.500000 283.650000 ;
      RECT 516.500000 282.350000 549.500000 283.650000 ;
      RECT 507.500000 282.350000 508.500000 283.650000 ;
      RECT 466.500000 282.350000 499.500000 283.650000 ;
      RECT 457.500000 282.350000 458.500000 283.650000 ;
      RECT 416.500000 282.350000 449.500000 283.650000 ;
      RECT 407.500000 282.350000 408.500000 283.650000 ;
      RECT 366.500000 282.350000 399.500000 283.650000 ;
      RECT 357.500000 282.350000 358.500000 283.650000 ;
      RECT 316.500000 282.350000 349.500000 283.650000 ;
      RECT 307.500000 282.350000 308.500000 283.650000 ;
      RECT 266.500000 282.350000 299.500000 283.650000 ;
      RECT 257.500000 282.350000 258.500000 283.650000 ;
      RECT 216.500000 282.350000 249.500000 283.650000 ;
      RECT 207.500000 282.350000 208.500000 283.650000 ;
      RECT 166.500000 282.350000 199.500000 283.650000 ;
      RECT 157.500000 282.350000 158.500000 283.650000 ;
      RECT 116.500000 282.350000 149.500000 283.650000 ;
      RECT 107.500000 282.350000 108.500000 283.650000 ;
      RECT 66.500000 282.350000 99.500000 283.650000 ;
      RECT 57.500000 282.350000 58.500000 283.650000 ;
      RECT 29.500000 282.350000 49.500000 283.650000 ;
      RECT 15.500000 282.350000 16.500000 283.650000 ;
      RECT 1157.500000 281.650000 1170.500000 282.350000 ;
      RECT 1107.500000 281.650000 1149.500000 282.350000 ;
      RECT 1057.500000 281.650000 1099.500000 282.350000 ;
      RECT 1007.500000 281.650000 1049.500000 282.350000 ;
      RECT 957.500000 281.650000 999.500000 282.350000 ;
      RECT 907.500000 281.650000 949.500000 282.350000 ;
      RECT 857.500000 281.650000 899.500000 282.350000 ;
      RECT 807.500000 281.650000 849.500000 282.350000 ;
      RECT 757.500000 281.650000 799.500000 282.350000 ;
      RECT 707.500000 281.650000 749.500000 282.350000 ;
      RECT 657.500000 281.650000 699.500000 282.350000 ;
      RECT 607.500000 281.650000 649.500000 282.350000 ;
      RECT 557.500000 281.650000 599.500000 282.350000 ;
      RECT 507.500000 281.650000 549.500000 282.350000 ;
      RECT 457.500000 281.650000 499.500000 282.350000 ;
      RECT 407.500000 281.650000 449.500000 282.350000 ;
      RECT 357.500000 281.650000 399.500000 282.350000 ;
      RECT 307.500000 281.650000 349.500000 282.350000 ;
      RECT 257.500000 281.650000 299.500000 282.350000 ;
      RECT 207.500000 281.650000 249.500000 282.350000 ;
      RECT 157.500000 281.650000 199.500000 282.350000 ;
      RECT 107.500000 281.650000 149.500000 282.350000 ;
      RECT 57.500000 281.650000 99.500000 282.350000 ;
      RECT 15.500000 281.650000 49.500000 282.350000 ;
      RECT 1183.500000 280.350000 1186.000000 283.650000 ;
      RECT 1169.500000 280.350000 1170.500000 281.650000 ;
      RECT 1116.500000 280.350000 1149.500000 281.650000 ;
      RECT 1107.500000 280.350000 1108.500000 281.650000 ;
      RECT 1066.500000 280.350000 1099.500000 281.650000 ;
      RECT 1057.500000 280.350000 1058.500000 281.650000 ;
      RECT 1016.500000 280.350000 1049.500000 281.650000 ;
      RECT 1007.500000 280.350000 1008.500000 281.650000 ;
      RECT 966.500000 280.350000 999.500000 281.650000 ;
      RECT 957.500000 280.350000 958.500000 281.650000 ;
      RECT 916.500000 280.350000 949.500000 281.650000 ;
      RECT 907.500000 280.350000 908.500000 281.650000 ;
      RECT 866.500000 280.350000 899.500000 281.650000 ;
      RECT 857.500000 280.350000 858.500000 281.650000 ;
      RECT 816.500000 280.350000 849.500000 281.650000 ;
      RECT 807.500000 280.350000 808.500000 281.650000 ;
      RECT 766.500000 280.350000 799.500000 281.650000 ;
      RECT 757.500000 280.350000 758.500000 281.650000 ;
      RECT 716.500000 280.350000 749.500000 281.650000 ;
      RECT 707.500000 280.350000 708.500000 281.650000 ;
      RECT 666.500000 280.350000 699.500000 281.650000 ;
      RECT 657.500000 280.350000 658.500000 281.650000 ;
      RECT 616.500000 280.350000 649.500000 281.650000 ;
      RECT 607.500000 280.350000 608.500000 281.650000 ;
      RECT 566.500000 280.350000 599.500000 281.650000 ;
      RECT 557.500000 280.350000 558.500000 281.650000 ;
      RECT 516.500000 280.350000 549.500000 281.650000 ;
      RECT 507.500000 280.350000 508.500000 281.650000 ;
      RECT 466.500000 280.350000 499.500000 281.650000 ;
      RECT 457.500000 280.350000 458.500000 281.650000 ;
      RECT 416.500000 280.350000 449.500000 281.650000 ;
      RECT 407.500000 280.350000 408.500000 281.650000 ;
      RECT 366.500000 280.350000 399.500000 281.650000 ;
      RECT 357.500000 280.350000 358.500000 281.650000 ;
      RECT 316.500000 280.350000 349.500000 281.650000 ;
      RECT 307.500000 280.350000 308.500000 281.650000 ;
      RECT 266.500000 280.350000 299.500000 281.650000 ;
      RECT 257.500000 280.350000 258.500000 281.650000 ;
      RECT 216.500000 280.350000 249.500000 281.650000 ;
      RECT 207.500000 280.350000 208.500000 281.650000 ;
      RECT 166.500000 280.350000 199.500000 281.650000 ;
      RECT 157.500000 280.350000 158.500000 281.650000 ;
      RECT 116.500000 280.350000 149.500000 281.650000 ;
      RECT 107.500000 280.350000 108.500000 281.650000 ;
      RECT 66.500000 280.350000 99.500000 281.650000 ;
      RECT 57.500000 280.350000 58.500000 281.650000 ;
      RECT 29.500000 280.350000 49.500000 281.650000 ;
      RECT 15.500000 280.350000 16.500000 281.650000 ;
      RECT 0.000000 280.350000 2.500000 283.650000 ;
      RECT 1169.500000 279.650000 1186.000000 280.350000 ;
      RECT 1116.500000 279.650000 1156.500000 280.350000 ;
      RECT 1066.500000 279.650000 1108.500000 280.350000 ;
      RECT 1016.500000 279.650000 1058.500000 280.350000 ;
      RECT 966.500000 279.650000 1008.500000 280.350000 ;
      RECT 916.500000 279.650000 958.500000 280.350000 ;
      RECT 866.500000 279.650000 908.500000 280.350000 ;
      RECT 816.500000 279.650000 858.500000 280.350000 ;
      RECT 766.500000 279.650000 808.500000 280.350000 ;
      RECT 716.500000 279.650000 758.500000 280.350000 ;
      RECT 666.500000 279.650000 708.500000 280.350000 ;
      RECT 616.500000 279.650000 658.500000 280.350000 ;
      RECT 566.500000 279.650000 608.500000 280.350000 ;
      RECT 516.500000 279.650000 558.500000 280.350000 ;
      RECT 466.500000 279.650000 508.500000 280.350000 ;
      RECT 416.500000 279.650000 458.500000 280.350000 ;
      RECT 366.500000 279.650000 408.500000 280.350000 ;
      RECT 316.500000 279.650000 358.500000 280.350000 ;
      RECT 266.500000 279.650000 308.500000 280.350000 ;
      RECT 216.500000 279.650000 258.500000 280.350000 ;
      RECT 166.500000 279.650000 208.500000 280.350000 ;
      RECT 116.500000 279.650000 158.500000 280.350000 ;
      RECT 66.500000 279.650000 108.500000 280.350000 ;
      RECT 29.500000 279.650000 58.500000 280.350000 ;
      RECT 0.000000 279.650000 16.500000 280.350000 ;
      RECT 1169.500000 278.350000 1170.500000 279.650000 ;
      RECT 1116.500000 278.350000 1149.500000 279.650000 ;
      RECT 1107.500000 278.350000 1108.500000 279.650000 ;
      RECT 1066.500000 278.350000 1099.500000 279.650000 ;
      RECT 1057.500000 278.350000 1058.500000 279.650000 ;
      RECT 1016.500000 278.350000 1049.500000 279.650000 ;
      RECT 1007.500000 278.350000 1008.500000 279.650000 ;
      RECT 966.500000 278.350000 999.500000 279.650000 ;
      RECT 957.500000 278.350000 958.500000 279.650000 ;
      RECT 916.500000 278.350000 949.500000 279.650000 ;
      RECT 907.500000 278.350000 908.500000 279.650000 ;
      RECT 866.500000 278.350000 899.500000 279.650000 ;
      RECT 857.500000 278.350000 858.500000 279.650000 ;
      RECT 816.500000 278.350000 849.500000 279.650000 ;
      RECT 807.500000 278.350000 808.500000 279.650000 ;
      RECT 766.500000 278.350000 799.500000 279.650000 ;
      RECT 757.500000 278.350000 758.500000 279.650000 ;
      RECT 716.500000 278.350000 749.500000 279.650000 ;
      RECT 707.500000 278.350000 708.500000 279.650000 ;
      RECT 666.500000 278.350000 699.500000 279.650000 ;
      RECT 657.500000 278.350000 658.500000 279.650000 ;
      RECT 616.500000 278.350000 649.500000 279.650000 ;
      RECT 607.500000 278.350000 608.500000 279.650000 ;
      RECT 566.500000 278.350000 599.500000 279.650000 ;
      RECT 557.500000 278.350000 558.500000 279.650000 ;
      RECT 516.500000 278.350000 549.500000 279.650000 ;
      RECT 507.500000 278.350000 508.500000 279.650000 ;
      RECT 466.500000 278.350000 499.500000 279.650000 ;
      RECT 457.500000 278.350000 458.500000 279.650000 ;
      RECT 416.500000 278.350000 449.500000 279.650000 ;
      RECT 407.500000 278.350000 408.500000 279.650000 ;
      RECT 366.500000 278.350000 399.500000 279.650000 ;
      RECT 357.500000 278.350000 358.500000 279.650000 ;
      RECT 316.500000 278.350000 349.500000 279.650000 ;
      RECT 307.500000 278.350000 308.500000 279.650000 ;
      RECT 266.500000 278.350000 299.500000 279.650000 ;
      RECT 257.500000 278.350000 258.500000 279.650000 ;
      RECT 216.500000 278.350000 249.500000 279.650000 ;
      RECT 207.500000 278.350000 208.500000 279.650000 ;
      RECT 166.500000 278.350000 199.500000 279.650000 ;
      RECT 157.500000 278.350000 158.500000 279.650000 ;
      RECT 116.500000 278.350000 149.500000 279.650000 ;
      RECT 107.500000 278.350000 108.500000 279.650000 ;
      RECT 66.500000 278.350000 99.500000 279.650000 ;
      RECT 57.500000 278.350000 58.500000 279.650000 ;
      RECT 29.500000 278.350000 49.500000 279.650000 ;
      RECT 15.500000 278.350000 16.500000 279.650000 ;
      RECT 1157.500000 277.650000 1170.500000 278.350000 ;
      RECT 1107.500000 277.650000 1149.500000 278.350000 ;
      RECT 1057.500000 277.650000 1099.500000 278.350000 ;
      RECT 1007.500000 277.650000 1049.500000 278.350000 ;
      RECT 957.500000 277.650000 999.500000 278.350000 ;
      RECT 907.500000 277.650000 949.500000 278.350000 ;
      RECT 857.500000 277.650000 899.500000 278.350000 ;
      RECT 807.500000 277.650000 849.500000 278.350000 ;
      RECT 757.500000 277.650000 799.500000 278.350000 ;
      RECT 707.500000 277.650000 749.500000 278.350000 ;
      RECT 657.500000 277.650000 699.500000 278.350000 ;
      RECT 607.500000 277.650000 649.500000 278.350000 ;
      RECT 557.500000 277.650000 599.500000 278.350000 ;
      RECT 507.500000 277.650000 549.500000 278.350000 ;
      RECT 457.500000 277.650000 499.500000 278.350000 ;
      RECT 407.500000 277.650000 449.500000 278.350000 ;
      RECT 357.500000 277.650000 399.500000 278.350000 ;
      RECT 307.500000 277.650000 349.500000 278.350000 ;
      RECT 257.500000 277.650000 299.500000 278.350000 ;
      RECT 207.500000 277.650000 249.500000 278.350000 ;
      RECT 157.500000 277.650000 199.500000 278.350000 ;
      RECT 107.500000 277.650000 149.500000 278.350000 ;
      RECT 57.500000 277.650000 99.500000 278.350000 ;
      RECT 15.500000 277.650000 49.500000 278.350000 ;
      RECT 1183.500000 276.350000 1186.000000 279.650000 ;
      RECT 1169.500000 276.350000 1170.500000 277.650000 ;
      RECT 1116.500000 276.350000 1149.500000 277.650000 ;
      RECT 1107.500000 276.350000 1108.500000 277.650000 ;
      RECT 1066.500000 276.350000 1099.500000 277.650000 ;
      RECT 1057.500000 276.350000 1058.500000 277.650000 ;
      RECT 1016.500000 276.350000 1049.500000 277.650000 ;
      RECT 1007.500000 276.350000 1008.500000 277.650000 ;
      RECT 966.500000 276.350000 999.500000 277.650000 ;
      RECT 957.500000 276.350000 958.500000 277.650000 ;
      RECT 916.500000 276.350000 949.500000 277.650000 ;
      RECT 907.500000 276.350000 908.500000 277.650000 ;
      RECT 866.500000 276.350000 899.500000 277.650000 ;
      RECT 857.500000 276.350000 858.500000 277.650000 ;
      RECT 816.500000 276.350000 849.500000 277.650000 ;
      RECT 807.500000 276.350000 808.500000 277.650000 ;
      RECT 766.500000 276.350000 799.500000 277.650000 ;
      RECT 757.500000 276.350000 758.500000 277.650000 ;
      RECT 716.500000 276.350000 749.500000 277.650000 ;
      RECT 707.500000 276.350000 708.500000 277.650000 ;
      RECT 666.500000 276.350000 699.500000 277.650000 ;
      RECT 657.500000 276.350000 658.500000 277.650000 ;
      RECT 616.500000 276.350000 649.500000 277.650000 ;
      RECT 607.500000 276.350000 608.500000 277.650000 ;
      RECT 566.500000 276.350000 599.500000 277.650000 ;
      RECT 557.500000 276.350000 558.500000 277.650000 ;
      RECT 516.500000 276.350000 549.500000 277.650000 ;
      RECT 507.500000 276.350000 508.500000 277.650000 ;
      RECT 466.500000 276.350000 499.500000 277.650000 ;
      RECT 457.500000 276.350000 458.500000 277.650000 ;
      RECT 416.500000 276.350000 449.500000 277.650000 ;
      RECT 407.500000 276.350000 408.500000 277.650000 ;
      RECT 366.500000 276.350000 399.500000 277.650000 ;
      RECT 357.500000 276.350000 358.500000 277.650000 ;
      RECT 316.500000 276.350000 349.500000 277.650000 ;
      RECT 307.500000 276.350000 308.500000 277.650000 ;
      RECT 266.500000 276.350000 299.500000 277.650000 ;
      RECT 257.500000 276.350000 258.500000 277.650000 ;
      RECT 216.500000 276.350000 249.500000 277.650000 ;
      RECT 207.500000 276.350000 208.500000 277.650000 ;
      RECT 166.500000 276.350000 199.500000 277.650000 ;
      RECT 157.500000 276.350000 158.500000 277.650000 ;
      RECT 116.500000 276.350000 149.500000 277.650000 ;
      RECT 107.500000 276.350000 108.500000 277.650000 ;
      RECT 66.500000 276.350000 99.500000 277.650000 ;
      RECT 57.500000 276.350000 58.500000 277.650000 ;
      RECT 29.500000 276.350000 49.500000 277.650000 ;
      RECT 15.500000 276.350000 16.500000 277.650000 ;
      RECT 0.000000 276.350000 2.500000 279.650000 ;
      RECT 1169.500000 275.650000 1186.000000 276.350000 ;
      RECT 1116.500000 275.650000 1156.500000 276.350000 ;
      RECT 1066.500000 275.650000 1108.500000 276.350000 ;
      RECT 1016.500000 275.650000 1058.500000 276.350000 ;
      RECT 966.500000 275.650000 1008.500000 276.350000 ;
      RECT 916.500000 275.650000 958.500000 276.350000 ;
      RECT 866.500000 275.650000 908.500000 276.350000 ;
      RECT 816.500000 275.650000 858.500000 276.350000 ;
      RECT 766.500000 275.650000 808.500000 276.350000 ;
      RECT 716.500000 275.650000 758.500000 276.350000 ;
      RECT 666.500000 275.650000 708.500000 276.350000 ;
      RECT 616.500000 275.650000 658.500000 276.350000 ;
      RECT 566.500000 275.650000 608.500000 276.350000 ;
      RECT 516.500000 275.650000 558.500000 276.350000 ;
      RECT 466.500000 275.650000 508.500000 276.350000 ;
      RECT 416.500000 275.650000 458.500000 276.350000 ;
      RECT 366.500000 275.650000 408.500000 276.350000 ;
      RECT 316.500000 275.650000 358.500000 276.350000 ;
      RECT 266.500000 275.650000 308.500000 276.350000 ;
      RECT 216.500000 275.650000 258.500000 276.350000 ;
      RECT 166.500000 275.650000 208.500000 276.350000 ;
      RECT 116.500000 275.650000 158.500000 276.350000 ;
      RECT 66.500000 275.650000 108.500000 276.350000 ;
      RECT 29.500000 275.650000 58.500000 276.350000 ;
      RECT 0.000000 275.650000 16.500000 276.350000 ;
      RECT 1169.500000 274.350000 1170.500000 275.650000 ;
      RECT 1116.500000 274.350000 1149.500000 275.650000 ;
      RECT 1107.500000 274.350000 1108.500000 275.650000 ;
      RECT 1066.500000 274.350000 1099.500000 275.650000 ;
      RECT 1057.500000 274.350000 1058.500000 275.650000 ;
      RECT 1016.500000 274.350000 1049.500000 275.650000 ;
      RECT 1007.500000 274.350000 1008.500000 275.650000 ;
      RECT 966.500000 274.350000 999.500000 275.650000 ;
      RECT 957.500000 274.350000 958.500000 275.650000 ;
      RECT 916.500000 274.350000 949.500000 275.650000 ;
      RECT 907.500000 274.350000 908.500000 275.650000 ;
      RECT 866.500000 274.350000 899.500000 275.650000 ;
      RECT 857.500000 274.350000 858.500000 275.650000 ;
      RECT 816.500000 274.350000 849.500000 275.650000 ;
      RECT 807.500000 274.350000 808.500000 275.650000 ;
      RECT 766.500000 274.350000 799.500000 275.650000 ;
      RECT 757.500000 274.350000 758.500000 275.650000 ;
      RECT 716.500000 274.350000 749.500000 275.650000 ;
      RECT 707.500000 274.350000 708.500000 275.650000 ;
      RECT 666.500000 274.350000 699.500000 275.650000 ;
      RECT 657.500000 274.350000 658.500000 275.650000 ;
      RECT 616.500000 274.350000 649.500000 275.650000 ;
      RECT 607.500000 274.350000 608.500000 275.650000 ;
      RECT 566.500000 274.350000 599.500000 275.650000 ;
      RECT 557.500000 274.350000 558.500000 275.650000 ;
      RECT 516.500000 274.350000 549.500000 275.650000 ;
      RECT 507.500000 274.350000 508.500000 275.650000 ;
      RECT 466.500000 274.350000 499.500000 275.650000 ;
      RECT 457.500000 274.350000 458.500000 275.650000 ;
      RECT 416.500000 274.350000 449.500000 275.650000 ;
      RECT 407.500000 274.350000 408.500000 275.650000 ;
      RECT 366.500000 274.350000 399.500000 275.650000 ;
      RECT 357.500000 274.350000 358.500000 275.650000 ;
      RECT 316.500000 274.350000 349.500000 275.650000 ;
      RECT 307.500000 274.350000 308.500000 275.650000 ;
      RECT 266.500000 274.350000 299.500000 275.650000 ;
      RECT 257.500000 274.350000 258.500000 275.650000 ;
      RECT 216.500000 274.350000 249.500000 275.650000 ;
      RECT 207.500000 274.350000 208.500000 275.650000 ;
      RECT 166.500000 274.350000 199.500000 275.650000 ;
      RECT 157.500000 274.350000 158.500000 275.650000 ;
      RECT 116.500000 274.350000 149.500000 275.650000 ;
      RECT 107.500000 274.350000 108.500000 275.650000 ;
      RECT 66.500000 274.350000 99.500000 275.650000 ;
      RECT 57.500000 274.350000 58.500000 275.650000 ;
      RECT 29.500000 274.350000 49.500000 275.650000 ;
      RECT 15.500000 274.350000 16.500000 275.650000 ;
      RECT 1157.500000 273.650000 1170.500000 274.350000 ;
      RECT 1107.500000 273.650000 1149.500000 274.350000 ;
      RECT 1057.500000 273.650000 1099.500000 274.350000 ;
      RECT 1007.500000 273.650000 1049.500000 274.350000 ;
      RECT 957.500000 273.650000 999.500000 274.350000 ;
      RECT 907.500000 273.650000 949.500000 274.350000 ;
      RECT 857.500000 273.650000 899.500000 274.350000 ;
      RECT 807.500000 273.650000 849.500000 274.350000 ;
      RECT 757.500000 273.650000 799.500000 274.350000 ;
      RECT 707.500000 273.650000 749.500000 274.350000 ;
      RECT 657.500000 273.650000 699.500000 274.350000 ;
      RECT 607.500000 273.650000 649.500000 274.350000 ;
      RECT 557.500000 273.650000 599.500000 274.350000 ;
      RECT 507.500000 273.650000 549.500000 274.350000 ;
      RECT 457.500000 273.650000 499.500000 274.350000 ;
      RECT 407.500000 273.650000 449.500000 274.350000 ;
      RECT 357.500000 273.650000 399.500000 274.350000 ;
      RECT 307.500000 273.650000 349.500000 274.350000 ;
      RECT 257.500000 273.650000 299.500000 274.350000 ;
      RECT 207.500000 273.650000 249.500000 274.350000 ;
      RECT 157.500000 273.650000 199.500000 274.350000 ;
      RECT 107.500000 273.650000 149.500000 274.350000 ;
      RECT 57.500000 273.650000 99.500000 274.350000 ;
      RECT 15.500000 273.650000 49.500000 274.350000 ;
      RECT 1183.500000 272.350000 1186.000000 275.650000 ;
      RECT 1169.500000 272.350000 1170.500000 273.650000 ;
      RECT 1116.500000 272.350000 1149.500000 273.650000 ;
      RECT 1107.500000 272.350000 1108.500000 273.650000 ;
      RECT 1066.500000 272.350000 1099.500000 273.650000 ;
      RECT 1057.500000 272.350000 1058.500000 273.650000 ;
      RECT 1016.500000 272.350000 1049.500000 273.650000 ;
      RECT 1007.500000 272.350000 1008.500000 273.650000 ;
      RECT 966.500000 272.350000 999.500000 273.650000 ;
      RECT 957.500000 272.350000 958.500000 273.650000 ;
      RECT 916.500000 272.350000 949.500000 273.650000 ;
      RECT 907.500000 272.350000 908.500000 273.650000 ;
      RECT 866.500000 272.350000 899.500000 273.650000 ;
      RECT 857.500000 272.350000 858.500000 273.650000 ;
      RECT 816.500000 272.350000 849.500000 273.650000 ;
      RECT 807.500000 272.350000 808.500000 273.650000 ;
      RECT 766.500000 272.350000 799.500000 273.650000 ;
      RECT 757.500000 272.350000 758.500000 273.650000 ;
      RECT 716.500000 272.350000 749.500000 273.650000 ;
      RECT 707.500000 272.350000 708.500000 273.650000 ;
      RECT 666.500000 272.350000 699.500000 273.650000 ;
      RECT 657.500000 272.350000 658.500000 273.650000 ;
      RECT 616.500000 272.350000 649.500000 273.650000 ;
      RECT 607.500000 272.350000 608.500000 273.650000 ;
      RECT 566.500000 272.350000 599.500000 273.650000 ;
      RECT 557.500000 272.350000 558.500000 273.650000 ;
      RECT 516.500000 272.350000 549.500000 273.650000 ;
      RECT 507.500000 272.350000 508.500000 273.650000 ;
      RECT 466.500000 272.350000 499.500000 273.650000 ;
      RECT 457.500000 272.350000 458.500000 273.650000 ;
      RECT 416.500000 272.350000 449.500000 273.650000 ;
      RECT 407.500000 272.350000 408.500000 273.650000 ;
      RECT 366.500000 272.350000 399.500000 273.650000 ;
      RECT 357.500000 272.350000 358.500000 273.650000 ;
      RECT 316.500000 272.350000 349.500000 273.650000 ;
      RECT 307.500000 272.350000 308.500000 273.650000 ;
      RECT 266.500000 272.350000 299.500000 273.650000 ;
      RECT 257.500000 272.350000 258.500000 273.650000 ;
      RECT 216.500000 272.350000 249.500000 273.650000 ;
      RECT 207.500000 272.350000 208.500000 273.650000 ;
      RECT 166.500000 272.350000 199.500000 273.650000 ;
      RECT 157.500000 272.350000 158.500000 273.650000 ;
      RECT 116.500000 272.350000 149.500000 273.650000 ;
      RECT 107.500000 272.350000 108.500000 273.650000 ;
      RECT 66.500000 272.350000 99.500000 273.650000 ;
      RECT 57.500000 272.350000 58.500000 273.650000 ;
      RECT 29.500000 272.350000 49.500000 273.650000 ;
      RECT 15.500000 272.350000 16.500000 273.650000 ;
      RECT 0.000000 272.350000 2.500000 275.650000 ;
      RECT 1169.500000 271.650000 1186.000000 272.350000 ;
      RECT 1116.500000 271.650000 1156.500000 272.350000 ;
      RECT 1066.500000 271.650000 1108.500000 272.350000 ;
      RECT 1016.500000 271.650000 1058.500000 272.350000 ;
      RECT 966.500000 271.650000 1008.500000 272.350000 ;
      RECT 916.500000 271.650000 958.500000 272.350000 ;
      RECT 866.500000 271.650000 908.500000 272.350000 ;
      RECT 816.500000 271.650000 858.500000 272.350000 ;
      RECT 766.500000 271.650000 808.500000 272.350000 ;
      RECT 716.500000 271.650000 758.500000 272.350000 ;
      RECT 666.500000 271.650000 708.500000 272.350000 ;
      RECT 616.500000 271.650000 658.500000 272.350000 ;
      RECT 566.500000 271.650000 608.500000 272.350000 ;
      RECT 516.500000 271.650000 558.500000 272.350000 ;
      RECT 466.500000 271.650000 508.500000 272.350000 ;
      RECT 416.500000 271.650000 458.500000 272.350000 ;
      RECT 366.500000 271.650000 408.500000 272.350000 ;
      RECT 316.500000 271.650000 358.500000 272.350000 ;
      RECT 266.500000 271.650000 308.500000 272.350000 ;
      RECT 216.500000 271.650000 258.500000 272.350000 ;
      RECT 166.500000 271.650000 208.500000 272.350000 ;
      RECT 116.500000 271.650000 158.500000 272.350000 ;
      RECT 66.500000 271.650000 108.500000 272.350000 ;
      RECT 29.500000 271.650000 58.500000 272.350000 ;
      RECT 0.000000 271.650000 16.500000 272.350000 ;
      RECT 1169.500000 270.350000 1170.500000 271.650000 ;
      RECT 1116.500000 270.350000 1149.500000 271.650000 ;
      RECT 1107.500000 270.350000 1108.500000 271.650000 ;
      RECT 1066.500000 270.350000 1099.500000 271.650000 ;
      RECT 1057.500000 270.350000 1058.500000 271.650000 ;
      RECT 1016.500000 270.350000 1049.500000 271.650000 ;
      RECT 1007.500000 270.350000 1008.500000 271.650000 ;
      RECT 966.500000 270.350000 999.500000 271.650000 ;
      RECT 957.500000 270.350000 958.500000 271.650000 ;
      RECT 916.500000 270.350000 949.500000 271.650000 ;
      RECT 907.500000 270.350000 908.500000 271.650000 ;
      RECT 866.500000 270.350000 899.500000 271.650000 ;
      RECT 857.500000 270.350000 858.500000 271.650000 ;
      RECT 816.500000 270.350000 849.500000 271.650000 ;
      RECT 807.500000 270.350000 808.500000 271.650000 ;
      RECT 766.500000 270.350000 799.500000 271.650000 ;
      RECT 757.500000 270.350000 758.500000 271.650000 ;
      RECT 716.500000 270.350000 749.500000 271.650000 ;
      RECT 707.500000 270.350000 708.500000 271.650000 ;
      RECT 666.500000 270.350000 699.500000 271.650000 ;
      RECT 657.500000 270.350000 658.500000 271.650000 ;
      RECT 616.500000 270.350000 649.500000 271.650000 ;
      RECT 607.500000 270.350000 608.500000 271.650000 ;
      RECT 566.500000 270.350000 599.500000 271.650000 ;
      RECT 557.500000 270.350000 558.500000 271.650000 ;
      RECT 516.500000 270.350000 549.500000 271.650000 ;
      RECT 507.500000 270.350000 508.500000 271.650000 ;
      RECT 466.500000 270.350000 499.500000 271.650000 ;
      RECT 457.500000 270.350000 458.500000 271.650000 ;
      RECT 416.500000 270.350000 449.500000 271.650000 ;
      RECT 407.500000 270.350000 408.500000 271.650000 ;
      RECT 366.500000 270.350000 399.500000 271.650000 ;
      RECT 357.500000 270.350000 358.500000 271.650000 ;
      RECT 316.500000 270.350000 349.500000 271.650000 ;
      RECT 307.500000 270.350000 308.500000 271.650000 ;
      RECT 266.500000 270.350000 299.500000 271.650000 ;
      RECT 257.500000 270.350000 258.500000 271.650000 ;
      RECT 216.500000 270.350000 249.500000 271.650000 ;
      RECT 207.500000 270.350000 208.500000 271.650000 ;
      RECT 166.500000 270.350000 199.500000 271.650000 ;
      RECT 157.500000 270.350000 158.500000 271.650000 ;
      RECT 116.500000 270.350000 149.500000 271.650000 ;
      RECT 107.500000 270.350000 108.500000 271.650000 ;
      RECT 66.500000 270.350000 99.500000 271.650000 ;
      RECT 57.500000 270.350000 58.500000 271.650000 ;
      RECT 29.500000 270.350000 49.500000 271.650000 ;
      RECT 15.500000 270.350000 16.500000 271.650000 ;
      RECT 1157.500000 269.650000 1170.500000 270.350000 ;
      RECT 1107.500000 269.650000 1149.500000 270.350000 ;
      RECT 1057.500000 269.650000 1099.500000 270.350000 ;
      RECT 1007.500000 269.650000 1049.500000 270.350000 ;
      RECT 957.500000 269.650000 999.500000 270.350000 ;
      RECT 907.500000 269.650000 949.500000 270.350000 ;
      RECT 857.500000 269.650000 899.500000 270.350000 ;
      RECT 807.500000 269.650000 849.500000 270.350000 ;
      RECT 757.500000 269.650000 799.500000 270.350000 ;
      RECT 707.500000 269.650000 749.500000 270.350000 ;
      RECT 657.500000 269.650000 699.500000 270.350000 ;
      RECT 607.500000 269.650000 649.500000 270.350000 ;
      RECT 557.500000 269.650000 599.500000 270.350000 ;
      RECT 507.500000 269.650000 549.500000 270.350000 ;
      RECT 457.500000 269.650000 499.500000 270.350000 ;
      RECT 407.500000 269.650000 449.500000 270.350000 ;
      RECT 357.500000 269.650000 399.500000 270.350000 ;
      RECT 307.500000 269.650000 349.500000 270.350000 ;
      RECT 257.500000 269.650000 299.500000 270.350000 ;
      RECT 207.500000 269.650000 249.500000 270.350000 ;
      RECT 157.500000 269.650000 199.500000 270.350000 ;
      RECT 107.500000 269.650000 149.500000 270.350000 ;
      RECT 57.500000 269.650000 99.500000 270.350000 ;
      RECT 15.500000 269.650000 49.500000 270.350000 ;
      RECT 1183.500000 268.350000 1186.000000 271.650000 ;
      RECT 1169.500000 268.350000 1170.500000 269.650000 ;
      RECT 1116.500000 268.350000 1149.500000 269.650000 ;
      RECT 1107.500000 268.350000 1108.500000 269.650000 ;
      RECT 1066.500000 268.350000 1099.500000 269.650000 ;
      RECT 1057.500000 268.350000 1058.500000 269.650000 ;
      RECT 1016.500000 268.350000 1049.500000 269.650000 ;
      RECT 1007.500000 268.350000 1008.500000 269.650000 ;
      RECT 966.500000 268.350000 999.500000 269.650000 ;
      RECT 957.500000 268.350000 958.500000 269.650000 ;
      RECT 916.500000 268.350000 949.500000 269.650000 ;
      RECT 907.500000 268.350000 908.500000 269.650000 ;
      RECT 866.500000 268.350000 899.500000 269.650000 ;
      RECT 857.500000 268.350000 858.500000 269.650000 ;
      RECT 816.500000 268.350000 849.500000 269.650000 ;
      RECT 807.500000 268.350000 808.500000 269.650000 ;
      RECT 766.500000 268.350000 799.500000 269.650000 ;
      RECT 757.500000 268.350000 758.500000 269.650000 ;
      RECT 716.500000 268.350000 749.500000 269.650000 ;
      RECT 707.500000 268.350000 708.500000 269.650000 ;
      RECT 666.500000 268.350000 699.500000 269.650000 ;
      RECT 657.500000 268.350000 658.500000 269.650000 ;
      RECT 616.500000 268.350000 649.500000 269.650000 ;
      RECT 607.500000 268.350000 608.500000 269.650000 ;
      RECT 566.500000 268.350000 599.500000 269.650000 ;
      RECT 557.500000 268.350000 558.500000 269.650000 ;
      RECT 516.500000 268.350000 549.500000 269.650000 ;
      RECT 507.500000 268.350000 508.500000 269.650000 ;
      RECT 466.500000 268.350000 499.500000 269.650000 ;
      RECT 457.500000 268.350000 458.500000 269.650000 ;
      RECT 416.500000 268.350000 449.500000 269.650000 ;
      RECT 407.500000 268.350000 408.500000 269.650000 ;
      RECT 366.500000 268.350000 399.500000 269.650000 ;
      RECT 357.500000 268.350000 358.500000 269.650000 ;
      RECT 316.500000 268.350000 349.500000 269.650000 ;
      RECT 307.500000 268.350000 308.500000 269.650000 ;
      RECT 266.500000 268.350000 299.500000 269.650000 ;
      RECT 257.500000 268.350000 258.500000 269.650000 ;
      RECT 216.500000 268.350000 249.500000 269.650000 ;
      RECT 207.500000 268.350000 208.500000 269.650000 ;
      RECT 166.500000 268.350000 199.500000 269.650000 ;
      RECT 157.500000 268.350000 158.500000 269.650000 ;
      RECT 116.500000 268.350000 149.500000 269.650000 ;
      RECT 107.500000 268.350000 108.500000 269.650000 ;
      RECT 66.500000 268.350000 99.500000 269.650000 ;
      RECT 57.500000 268.350000 58.500000 269.650000 ;
      RECT 29.500000 268.350000 49.500000 269.650000 ;
      RECT 15.500000 268.350000 16.500000 269.650000 ;
      RECT 0.000000 268.350000 2.500000 271.650000 ;
      RECT 1169.500000 267.650000 1186.000000 268.350000 ;
      RECT 1116.500000 267.650000 1156.500000 268.350000 ;
      RECT 1066.500000 267.650000 1108.500000 268.350000 ;
      RECT 1016.500000 267.650000 1058.500000 268.350000 ;
      RECT 966.500000 267.650000 1008.500000 268.350000 ;
      RECT 916.500000 267.650000 958.500000 268.350000 ;
      RECT 866.500000 267.650000 908.500000 268.350000 ;
      RECT 816.500000 267.650000 858.500000 268.350000 ;
      RECT 766.500000 267.650000 808.500000 268.350000 ;
      RECT 716.500000 267.650000 758.500000 268.350000 ;
      RECT 666.500000 267.650000 708.500000 268.350000 ;
      RECT 616.500000 267.650000 658.500000 268.350000 ;
      RECT 566.500000 267.650000 608.500000 268.350000 ;
      RECT 516.500000 267.650000 558.500000 268.350000 ;
      RECT 466.500000 267.650000 508.500000 268.350000 ;
      RECT 416.500000 267.650000 458.500000 268.350000 ;
      RECT 366.500000 267.650000 408.500000 268.350000 ;
      RECT 316.500000 267.650000 358.500000 268.350000 ;
      RECT 266.500000 267.650000 308.500000 268.350000 ;
      RECT 216.500000 267.650000 258.500000 268.350000 ;
      RECT 166.500000 267.650000 208.500000 268.350000 ;
      RECT 116.500000 267.650000 158.500000 268.350000 ;
      RECT 66.500000 267.650000 108.500000 268.350000 ;
      RECT 29.500000 267.650000 58.500000 268.350000 ;
      RECT 0.000000 267.650000 16.500000 268.350000 ;
      RECT 1169.500000 266.350000 1170.500000 267.650000 ;
      RECT 1116.500000 266.350000 1149.500000 267.650000 ;
      RECT 1107.500000 266.350000 1108.500000 267.650000 ;
      RECT 1066.500000 266.350000 1099.500000 267.650000 ;
      RECT 1057.500000 266.350000 1058.500000 267.650000 ;
      RECT 1016.500000 266.350000 1049.500000 267.650000 ;
      RECT 1007.500000 266.350000 1008.500000 267.650000 ;
      RECT 966.500000 266.350000 999.500000 267.650000 ;
      RECT 957.500000 266.350000 958.500000 267.650000 ;
      RECT 916.500000 266.350000 949.500000 267.650000 ;
      RECT 907.500000 266.350000 908.500000 267.650000 ;
      RECT 866.500000 266.350000 899.500000 267.650000 ;
      RECT 857.500000 266.350000 858.500000 267.650000 ;
      RECT 816.500000 266.350000 849.500000 267.650000 ;
      RECT 807.500000 266.350000 808.500000 267.650000 ;
      RECT 766.500000 266.350000 799.500000 267.650000 ;
      RECT 757.500000 266.350000 758.500000 267.650000 ;
      RECT 716.500000 266.350000 749.500000 267.650000 ;
      RECT 707.500000 266.350000 708.500000 267.650000 ;
      RECT 666.500000 266.350000 699.500000 267.650000 ;
      RECT 657.500000 266.350000 658.500000 267.650000 ;
      RECT 616.500000 266.350000 649.500000 267.650000 ;
      RECT 607.500000 266.350000 608.500000 267.650000 ;
      RECT 566.500000 266.350000 599.500000 267.650000 ;
      RECT 557.500000 266.350000 558.500000 267.650000 ;
      RECT 516.500000 266.350000 549.500000 267.650000 ;
      RECT 507.500000 266.350000 508.500000 267.650000 ;
      RECT 466.500000 266.350000 499.500000 267.650000 ;
      RECT 457.500000 266.350000 458.500000 267.650000 ;
      RECT 416.500000 266.350000 449.500000 267.650000 ;
      RECT 407.500000 266.350000 408.500000 267.650000 ;
      RECT 366.500000 266.350000 399.500000 267.650000 ;
      RECT 357.500000 266.350000 358.500000 267.650000 ;
      RECT 316.500000 266.350000 349.500000 267.650000 ;
      RECT 307.500000 266.350000 308.500000 267.650000 ;
      RECT 266.500000 266.350000 299.500000 267.650000 ;
      RECT 257.500000 266.350000 258.500000 267.650000 ;
      RECT 216.500000 266.350000 249.500000 267.650000 ;
      RECT 207.500000 266.350000 208.500000 267.650000 ;
      RECT 166.500000 266.350000 199.500000 267.650000 ;
      RECT 157.500000 266.350000 158.500000 267.650000 ;
      RECT 116.500000 266.350000 149.500000 267.650000 ;
      RECT 107.500000 266.350000 108.500000 267.650000 ;
      RECT 66.500000 266.350000 99.500000 267.650000 ;
      RECT 57.500000 266.350000 58.500000 267.650000 ;
      RECT 29.500000 266.350000 49.500000 267.650000 ;
      RECT 15.500000 266.350000 16.500000 267.650000 ;
      RECT 1157.500000 265.650000 1170.500000 266.350000 ;
      RECT 1107.500000 265.650000 1149.500000 266.350000 ;
      RECT 1057.500000 265.650000 1099.500000 266.350000 ;
      RECT 1007.500000 265.650000 1049.500000 266.350000 ;
      RECT 957.500000 265.650000 999.500000 266.350000 ;
      RECT 907.500000 265.650000 949.500000 266.350000 ;
      RECT 857.500000 265.650000 899.500000 266.350000 ;
      RECT 807.500000 265.650000 849.500000 266.350000 ;
      RECT 757.500000 265.650000 799.500000 266.350000 ;
      RECT 707.500000 265.650000 749.500000 266.350000 ;
      RECT 657.500000 265.650000 699.500000 266.350000 ;
      RECT 607.500000 265.650000 649.500000 266.350000 ;
      RECT 557.500000 265.650000 599.500000 266.350000 ;
      RECT 507.500000 265.650000 549.500000 266.350000 ;
      RECT 457.500000 265.650000 499.500000 266.350000 ;
      RECT 407.500000 265.650000 449.500000 266.350000 ;
      RECT 357.500000 265.650000 399.500000 266.350000 ;
      RECT 307.500000 265.650000 349.500000 266.350000 ;
      RECT 257.500000 265.650000 299.500000 266.350000 ;
      RECT 207.500000 265.650000 249.500000 266.350000 ;
      RECT 157.500000 265.650000 199.500000 266.350000 ;
      RECT 107.500000 265.650000 149.500000 266.350000 ;
      RECT 57.500000 265.650000 99.500000 266.350000 ;
      RECT 15.500000 265.650000 49.500000 266.350000 ;
      RECT 1183.500000 264.350000 1186.000000 267.650000 ;
      RECT 1169.500000 264.350000 1170.500000 265.650000 ;
      RECT 1116.500000 264.350000 1149.500000 265.650000 ;
      RECT 1107.500000 264.350000 1108.500000 265.650000 ;
      RECT 1066.500000 264.350000 1099.500000 265.650000 ;
      RECT 1057.500000 264.350000 1058.500000 265.650000 ;
      RECT 1016.500000 264.350000 1049.500000 265.650000 ;
      RECT 1007.500000 264.350000 1008.500000 265.650000 ;
      RECT 966.500000 264.350000 999.500000 265.650000 ;
      RECT 957.500000 264.350000 958.500000 265.650000 ;
      RECT 916.500000 264.350000 949.500000 265.650000 ;
      RECT 907.500000 264.350000 908.500000 265.650000 ;
      RECT 866.500000 264.350000 899.500000 265.650000 ;
      RECT 857.500000 264.350000 858.500000 265.650000 ;
      RECT 816.500000 264.350000 849.500000 265.650000 ;
      RECT 807.500000 264.350000 808.500000 265.650000 ;
      RECT 766.500000 264.350000 799.500000 265.650000 ;
      RECT 757.500000 264.350000 758.500000 265.650000 ;
      RECT 716.500000 264.350000 749.500000 265.650000 ;
      RECT 707.500000 264.350000 708.500000 265.650000 ;
      RECT 666.500000 264.350000 699.500000 265.650000 ;
      RECT 657.500000 264.350000 658.500000 265.650000 ;
      RECT 616.500000 264.350000 649.500000 265.650000 ;
      RECT 607.500000 264.350000 608.500000 265.650000 ;
      RECT 566.500000 264.350000 599.500000 265.650000 ;
      RECT 557.500000 264.350000 558.500000 265.650000 ;
      RECT 516.500000 264.350000 549.500000 265.650000 ;
      RECT 507.500000 264.350000 508.500000 265.650000 ;
      RECT 466.500000 264.350000 499.500000 265.650000 ;
      RECT 457.500000 264.350000 458.500000 265.650000 ;
      RECT 416.500000 264.350000 449.500000 265.650000 ;
      RECT 407.500000 264.350000 408.500000 265.650000 ;
      RECT 366.500000 264.350000 399.500000 265.650000 ;
      RECT 357.500000 264.350000 358.500000 265.650000 ;
      RECT 316.500000 264.350000 349.500000 265.650000 ;
      RECT 307.500000 264.350000 308.500000 265.650000 ;
      RECT 266.500000 264.350000 299.500000 265.650000 ;
      RECT 257.500000 264.350000 258.500000 265.650000 ;
      RECT 216.500000 264.350000 249.500000 265.650000 ;
      RECT 207.500000 264.350000 208.500000 265.650000 ;
      RECT 166.500000 264.350000 199.500000 265.650000 ;
      RECT 157.500000 264.350000 158.500000 265.650000 ;
      RECT 116.500000 264.350000 149.500000 265.650000 ;
      RECT 107.500000 264.350000 108.500000 265.650000 ;
      RECT 66.500000 264.350000 99.500000 265.650000 ;
      RECT 57.500000 264.350000 58.500000 265.650000 ;
      RECT 29.500000 264.350000 49.500000 265.650000 ;
      RECT 15.500000 264.350000 16.500000 265.650000 ;
      RECT 0.000000 264.350000 2.500000 267.650000 ;
      RECT 1169.500000 263.650000 1186.000000 264.350000 ;
      RECT 1116.500000 263.650000 1156.500000 264.350000 ;
      RECT 1066.500000 263.650000 1108.500000 264.350000 ;
      RECT 1016.500000 263.650000 1058.500000 264.350000 ;
      RECT 966.500000 263.650000 1008.500000 264.350000 ;
      RECT 916.500000 263.650000 958.500000 264.350000 ;
      RECT 866.500000 263.650000 908.500000 264.350000 ;
      RECT 816.500000 263.650000 858.500000 264.350000 ;
      RECT 766.500000 263.650000 808.500000 264.350000 ;
      RECT 716.500000 263.650000 758.500000 264.350000 ;
      RECT 666.500000 263.650000 708.500000 264.350000 ;
      RECT 616.500000 263.650000 658.500000 264.350000 ;
      RECT 566.500000 263.650000 608.500000 264.350000 ;
      RECT 516.500000 263.650000 558.500000 264.350000 ;
      RECT 466.500000 263.650000 508.500000 264.350000 ;
      RECT 416.500000 263.650000 458.500000 264.350000 ;
      RECT 366.500000 263.650000 408.500000 264.350000 ;
      RECT 316.500000 263.650000 358.500000 264.350000 ;
      RECT 266.500000 263.650000 308.500000 264.350000 ;
      RECT 216.500000 263.650000 258.500000 264.350000 ;
      RECT 166.500000 263.650000 208.500000 264.350000 ;
      RECT 116.500000 263.650000 158.500000 264.350000 ;
      RECT 66.500000 263.650000 108.500000 264.350000 ;
      RECT 29.500000 263.650000 58.500000 264.350000 ;
      RECT 0.000000 263.650000 16.500000 264.350000 ;
      RECT 1169.500000 262.350000 1170.500000 263.650000 ;
      RECT 1116.500000 262.350000 1149.500000 263.650000 ;
      RECT 1107.500000 262.350000 1108.500000 263.650000 ;
      RECT 1066.500000 262.350000 1099.500000 263.650000 ;
      RECT 1057.500000 262.350000 1058.500000 263.650000 ;
      RECT 1016.500000 262.350000 1049.500000 263.650000 ;
      RECT 1007.500000 262.350000 1008.500000 263.650000 ;
      RECT 966.500000 262.350000 999.500000 263.650000 ;
      RECT 957.500000 262.350000 958.500000 263.650000 ;
      RECT 916.500000 262.350000 949.500000 263.650000 ;
      RECT 907.500000 262.350000 908.500000 263.650000 ;
      RECT 866.500000 262.350000 899.500000 263.650000 ;
      RECT 857.500000 262.350000 858.500000 263.650000 ;
      RECT 816.500000 262.350000 849.500000 263.650000 ;
      RECT 807.500000 262.350000 808.500000 263.650000 ;
      RECT 766.500000 262.350000 799.500000 263.650000 ;
      RECT 757.500000 262.350000 758.500000 263.650000 ;
      RECT 716.500000 262.350000 749.500000 263.650000 ;
      RECT 707.500000 262.350000 708.500000 263.650000 ;
      RECT 666.500000 262.350000 699.500000 263.650000 ;
      RECT 657.500000 262.350000 658.500000 263.650000 ;
      RECT 616.500000 262.350000 649.500000 263.650000 ;
      RECT 607.500000 262.350000 608.500000 263.650000 ;
      RECT 566.500000 262.350000 599.500000 263.650000 ;
      RECT 557.500000 262.350000 558.500000 263.650000 ;
      RECT 516.500000 262.350000 549.500000 263.650000 ;
      RECT 507.500000 262.350000 508.500000 263.650000 ;
      RECT 466.500000 262.350000 499.500000 263.650000 ;
      RECT 457.500000 262.350000 458.500000 263.650000 ;
      RECT 416.500000 262.350000 449.500000 263.650000 ;
      RECT 407.500000 262.350000 408.500000 263.650000 ;
      RECT 366.500000 262.350000 399.500000 263.650000 ;
      RECT 357.500000 262.350000 358.500000 263.650000 ;
      RECT 316.500000 262.350000 349.500000 263.650000 ;
      RECT 307.500000 262.350000 308.500000 263.650000 ;
      RECT 266.500000 262.350000 299.500000 263.650000 ;
      RECT 257.500000 262.350000 258.500000 263.650000 ;
      RECT 216.500000 262.350000 249.500000 263.650000 ;
      RECT 207.500000 262.350000 208.500000 263.650000 ;
      RECT 166.500000 262.350000 199.500000 263.650000 ;
      RECT 157.500000 262.350000 158.500000 263.650000 ;
      RECT 116.500000 262.350000 149.500000 263.650000 ;
      RECT 107.500000 262.350000 108.500000 263.650000 ;
      RECT 66.500000 262.350000 99.500000 263.650000 ;
      RECT 57.500000 262.350000 58.500000 263.650000 ;
      RECT 29.500000 262.350000 49.500000 263.650000 ;
      RECT 15.500000 262.350000 16.500000 263.650000 ;
      RECT 1157.500000 261.650000 1170.500000 262.350000 ;
      RECT 1107.500000 261.650000 1149.500000 262.350000 ;
      RECT 1057.500000 261.650000 1099.500000 262.350000 ;
      RECT 1007.500000 261.650000 1049.500000 262.350000 ;
      RECT 957.500000 261.650000 999.500000 262.350000 ;
      RECT 907.500000 261.650000 949.500000 262.350000 ;
      RECT 857.500000 261.650000 899.500000 262.350000 ;
      RECT 807.500000 261.650000 849.500000 262.350000 ;
      RECT 757.500000 261.650000 799.500000 262.350000 ;
      RECT 707.500000 261.650000 749.500000 262.350000 ;
      RECT 657.500000 261.650000 699.500000 262.350000 ;
      RECT 607.500000 261.650000 649.500000 262.350000 ;
      RECT 557.500000 261.650000 599.500000 262.350000 ;
      RECT 507.500000 261.650000 549.500000 262.350000 ;
      RECT 457.500000 261.650000 499.500000 262.350000 ;
      RECT 407.500000 261.650000 449.500000 262.350000 ;
      RECT 357.500000 261.650000 399.500000 262.350000 ;
      RECT 307.500000 261.650000 349.500000 262.350000 ;
      RECT 257.500000 261.650000 299.500000 262.350000 ;
      RECT 207.500000 261.650000 249.500000 262.350000 ;
      RECT 157.500000 261.650000 199.500000 262.350000 ;
      RECT 107.500000 261.650000 149.500000 262.350000 ;
      RECT 57.500000 261.650000 99.500000 262.350000 ;
      RECT 15.500000 261.650000 49.500000 262.350000 ;
      RECT 1183.500000 260.350000 1186.000000 263.650000 ;
      RECT 1169.500000 260.350000 1170.500000 261.650000 ;
      RECT 1116.500000 260.350000 1149.500000 261.650000 ;
      RECT 1107.500000 260.350000 1108.500000 261.650000 ;
      RECT 1066.500000 260.350000 1099.500000 261.650000 ;
      RECT 1057.500000 260.350000 1058.500000 261.650000 ;
      RECT 1016.500000 260.350000 1049.500000 261.650000 ;
      RECT 1007.500000 260.350000 1008.500000 261.650000 ;
      RECT 966.500000 260.350000 999.500000 261.650000 ;
      RECT 957.500000 260.350000 958.500000 261.650000 ;
      RECT 916.500000 260.350000 949.500000 261.650000 ;
      RECT 907.500000 260.350000 908.500000 261.650000 ;
      RECT 866.500000 260.350000 899.500000 261.650000 ;
      RECT 857.500000 260.350000 858.500000 261.650000 ;
      RECT 816.500000 260.350000 849.500000 261.650000 ;
      RECT 807.500000 260.350000 808.500000 261.650000 ;
      RECT 766.500000 260.350000 799.500000 261.650000 ;
      RECT 757.500000 260.350000 758.500000 261.650000 ;
      RECT 716.500000 260.350000 749.500000 261.650000 ;
      RECT 707.500000 260.350000 708.500000 261.650000 ;
      RECT 666.500000 260.350000 699.500000 261.650000 ;
      RECT 657.500000 260.350000 658.500000 261.650000 ;
      RECT 616.500000 260.350000 649.500000 261.650000 ;
      RECT 607.500000 260.350000 608.500000 261.650000 ;
      RECT 566.500000 260.350000 599.500000 261.650000 ;
      RECT 557.500000 260.350000 558.500000 261.650000 ;
      RECT 516.500000 260.350000 549.500000 261.650000 ;
      RECT 507.500000 260.350000 508.500000 261.650000 ;
      RECT 466.500000 260.350000 499.500000 261.650000 ;
      RECT 457.500000 260.350000 458.500000 261.650000 ;
      RECT 416.500000 260.350000 449.500000 261.650000 ;
      RECT 407.500000 260.350000 408.500000 261.650000 ;
      RECT 366.500000 260.350000 399.500000 261.650000 ;
      RECT 357.500000 260.350000 358.500000 261.650000 ;
      RECT 316.500000 260.350000 349.500000 261.650000 ;
      RECT 307.500000 260.350000 308.500000 261.650000 ;
      RECT 266.500000 260.350000 299.500000 261.650000 ;
      RECT 257.500000 260.350000 258.500000 261.650000 ;
      RECT 216.500000 260.350000 249.500000 261.650000 ;
      RECT 207.500000 260.350000 208.500000 261.650000 ;
      RECT 166.500000 260.350000 199.500000 261.650000 ;
      RECT 157.500000 260.350000 158.500000 261.650000 ;
      RECT 116.500000 260.350000 149.500000 261.650000 ;
      RECT 107.500000 260.350000 108.500000 261.650000 ;
      RECT 66.500000 260.350000 99.500000 261.650000 ;
      RECT 57.500000 260.350000 58.500000 261.650000 ;
      RECT 29.500000 260.350000 49.500000 261.650000 ;
      RECT 15.500000 260.350000 16.500000 261.650000 ;
      RECT 0.000000 260.350000 2.500000 263.650000 ;
      RECT 1169.500000 259.650000 1186.000000 260.350000 ;
      RECT 1116.500000 259.650000 1156.500000 260.350000 ;
      RECT 1169.500000 258.350000 1170.500000 259.650000 ;
      RECT 1116.500000 258.350000 1149.500000 259.650000 ;
      RECT 1066.500000 258.350000 1108.500000 260.350000 ;
      RECT 1016.500000 258.350000 1058.500000 260.350000 ;
      RECT 966.500000 258.350000 1008.500000 260.350000 ;
      RECT 916.500000 258.350000 958.500000 260.350000 ;
      RECT 866.500000 258.350000 908.500000 260.350000 ;
      RECT 816.500000 258.350000 858.500000 260.350000 ;
      RECT 766.500000 258.350000 808.500000 260.350000 ;
      RECT 716.500000 258.350000 758.500000 260.350000 ;
      RECT 666.500000 258.350000 708.500000 260.350000 ;
      RECT 616.500000 258.350000 658.500000 260.350000 ;
      RECT 566.500000 258.350000 608.500000 260.350000 ;
      RECT 516.500000 258.350000 558.500000 260.350000 ;
      RECT 466.500000 258.350000 508.500000 260.350000 ;
      RECT 416.500000 258.350000 458.500000 260.350000 ;
      RECT 366.500000 258.350000 408.500000 260.350000 ;
      RECT 316.500000 258.350000 358.500000 260.350000 ;
      RECT 266.500000 258.350000 308.500000 260.350000 ;
      RECT 216.500000 258.350000 258.500000 260.350000 ;
      RECT 166.500000 258.350000 208.500000 260.350000 ;
      RECT 116.500000 258.350000 158.500000 260.350000 ;
      RECT 66.500000 258.350000 108.500000 260.350000 ;
      RECT 29.500000 258.350000 58.500000 260.350000 ;
      RECT 0.000000 258.350000 16.500000 260.350000 ;
      RECT 1157.500000 257.650000 1170.500000 258.350000 ;
      RECT 1183.500000 256.350000 1186.000000 259.650000 ;
      RECT 1169.500000 256.350000 1170.500000 257.650000 ;
      RECT 0.000000 256.350000 1149.500000 258.350000 ;
      RECT 1169.500000 255.650000 1186.000000 256.350000 ;
      RECT 1169.500000 254.350000 1170.500000 255.650000 ;
      RECT 0.000000 254.350000 1156.500000 256.350000 ;
      RECT 0.000000 253.650000 1170.500000 254.350000 ;
      RECT 1183.500000 252.350000 1186.000000 255.650000 ;
      RECT 1169.500000 252.350000 1170.500000 253.650000 ;
      RECT 1169.500000 251.650000 1186.000000 252.350000 ;
      RECT 1169.500000 250.350000 1170.500000 251.650000 ;
      RECT 0.000000 250.350000 1156.500000 253.650000 ;
      RECT 0.000000 249.650000 1170.500000 250.350000 ;
      RECT 1183.500000 248.350000 1186.000000 251.650000 ;
      RECT 1169.500000 248.350000 1170.500000 249.650000 ;
      RECT 1169.500000 247.650000 1186.000000 248.350000 ;
      RECT 1169.500000 246.350000 1170.500000 247.650000 ;
      RECT 0.000000 246.350000 1156.500000 249.650000 ;
      RECT 0.000000 245.650000 1170.500000 246.350000 ;
      RECT 1183.500000 244.350000 1186.000000 247.650000 ;
      RECT 1169.500000 244.350000 1170.500000 245.650000 ;
      RECT 1169.500000 243.650000 1186.000000 244.350000 ;
      RECT 1169.500000 242.350000 1170.500000 243.650000 ;
      RECT 0.000000 242.350000 1156.500000 245.650000 ;
      RECT 0.000000 241.650000 1170.500000 242.350000 ;
      RECT 1183.500000 240.350000 1186.000000 243.650000 ;
      RECT 1169.500000 240.350000 1170.500000 241.650000 ;
      RECT 1169.500000 239.650000 1186.000000 240.350000 ;
      RECT 1169.500000 238.350000 1170.500000 239.650000 ;
      RECT 0.000000 238.350000 1156.500000 241.650000 ;
      RECT 0.000000 237.650000 1170.500000 238.350000 ;
      RECT 1183.500000 236.350000 1186.000000 239.650000 ;
      RECT 1169.500000 236.350000 1170.500000 237.650000 ;
      RECT 1169.500000 235.650000 1186.000000 236.350000 ;
      RECT 1169.500000 234.350000 1170.500000 235.650000 ;
      RECT 0.000000 234.350000 1156.500000 237.650000 ;
      RECT 0.000000 233.650000 1170.500000 234.350000 ;
      RECT 1183.500000 232.350000 1186.000000 235.650000 ;
      RECT 1169.500000 232.350000 1170.500000 233.650000 ;
      RECT 1169.500000 231.650000 1186.000000 232.350000 ;
      RECT 1169.500000 230.350000 1170.500000 231.650000 ;
      RECT 0.000000 230.350000 1156.500000 233.650000 ;
      RECT 0.000000 229.650000 1170.500000 230.350000 ;
      RECT 1183.500000 228.350000 1186.000000 231.650000 ;
      RECT 1169.500000 228.350000 1170.500000 229.650000 ;
      RECT 1169.500000 227.650000 1186.000000 228.350000 ;
      RECT 1169.500000 226.350000 1170.500000 227.650000 ;
      RECT 0.000000 226.350000 1156.500000 229.650000 ;
      RECT 0.000000 225.650000 1170.500000 226.350000 ;
      RECT 1183.500000 224.350000 1186.000000 227.650000 ;
      RECT 1169.500000 224.350000 1170.500000 225.650000 ;
      RECT 1169.500000 223.650000 1186.000000 224.350000 ;
      RECT 0.000000 223.170000 1156.500000 225.650000 ;
      RECT 1183.500000 223.165000 1186.000000 223.650000 ;
      RECT 1169.500000 222.350000 1170.500000 223.650000 ;
      RECT 2.020000 222.350000 1156.500000 223.170000 ;
      RECT 2.020000 221.650000 1170.500000 222.350000 ;
      RECT 1183.500000 220.350000 1183.980000 223.165000 ;
      RECT 1169.500000 220.350000 1170.500000 221.650000 ;
      RECT 2.020000 220.070000 1156.500000 221.650000 ;
      RECT 1169.500000 220.065000 1183.980000 220.350000 ;
      RECT 1169.500000 219.650000 1186.000000 220.065000 ;
      RECT 1169.500000 218.350000 1170.500000 219.650000 ;
      RECT 0.000000 218.350000 1156.500000 220.070000 ;
      RECT 0.000000 217.650000 1170.500000 218.350000 ;
      RECT 1183.500000 217.485000 1186.000000 219.650000 ;
      RECT 1183.500000 216.350000 1183.980000 217.485000 ;
      RECT 1169.500000 216.350000 1170.500000 217.650000 ;
      RECT 1169.500000 215.650000 1183.980000 216.350000 ;
      RECT 1183.500000 214.385000 1183.980000 215.650000 ;
      RECT 1169.500000 214.350000 1170.500000 215.650000 ;
      RECT 0.000000 214.350000 1156.500000 217.650000 ;
      RECT 0.000000 213.650000 1170.500000 214.350000 ;
      RECT 1183.500000 213.525000 1186.000000 214.385000 ;
      RECT 0.000000 212.575000 1156.500000 213.650000 ;
      RECT 1183.500000 212.350000 1183.980000 213.525000 ;
      RECT 1169.500000 212.350000 1170.500000 213.650000 ;
      RECT 1169.500000 211.650000 1183.980000 212.350000 ;
      RECT 1183.500000 210.425000 1183.980000 211.650000 ;
      RECT 1169.500000 210.350000 1170.500000 211.650000 ;
      RECT 2.020000 210.350000 1156.500000 212.575000 ;
      RECT 2.020000 209.650000 1170.500000 210.350000 ;
      RECT 2.020000 209.475000 1156.500000 209.650000 ;
      RECT 0.000000 208.615000 1156.500000 209.475000 ;
      RECT 1183.500000 208.350000 1186.000000 210.425000 ;
      RECT 1169.500000 208.350000 1170.500000 209.650000 ;
      RECT 1169.500000 207.650000 1186.000000 208.350000 ;
      RECT 1169.500000 206.350000 1170.500000 207.650000 ;
      RECT 2.020000 206.350000 1156.500000 208.615000 ;
      RECT 2.020000 205.650000 1170.500000 206.350000 ;
      RECT 2.020000 205.515000 1156.500000 205.650000 ;
      RECT 1183.500000 204.350000 1186.000000 207.650000 ;
      RECT 1169.500000 204.350000 1170.500000 205.650000 ;
      RECT 1169.500000 203.650000 1186.000000 204.350000 ;
      RECT 0.000000 202.935000 1156.500000 205.515000 ;
      RECT 1183.500000 202.930000 1186.000000 203.650000 ;
      RECT 1169.500000 202.350000 1170.500000 203.650000 ;
      RECT 2.020000 202.350000 1156.500000 202.935000 ;
      RECT 2.020000 201.650000 1170.500000 202.350000 ;
      RECT 1183.500000 200.350000 1183.980000 202.930000 ;
      RECT 1169.500000 200.350000 1170.500000 201.650000 ;
      RECT 2.020000 199.835000 1156.500000 201.650000 ;
      RECT 1169.500000 199.830000 1183.980000 200.350000 ;
      RECT 1169.500000 199.650000 1186.000000 199.830000 ;
      RECT 1169.500000 198.350000 1170.500000 199.650000 ;
      RECT 0.000000 198.350000 1156.500000 199.835000 ;
      RECT 0.000000 197.650000 1170.500000 198.350000 ;
      RECT 1183.500000 196.350000 1186.000000 199.650000 ;
      RECT 1169.500000 196.350000 1170.500000 197.650000 ;
      RECT 1169.500000 195.650000 1186.000000 196.350000 ;
      RECT 1169.500000 194.350000 1170.500000 195.650000 ;
      RECT 0.000000 194.350000 1156.500000 197.650000 ;
      RECT 0.000000 193.650000 1170.500000 194.350000 ;
      RECT 1183.500000 192.350000 1186.000000 195.650000 ;
      RECT 1169.500000 192.350000 1170.500000 193.650000 ;
      RECT 1169.500000 191.650000 1186.000000 192.350000 ;
      RECT 1169.500000 190.350000 1170.500000 191.650000 ;
      RECT 0.000000 190.350000 1156.500000 193.650000 ;
      RECT 0.000000 189.650000 1170.500000 190.350000 ;
      RECT 1183.500000 188.350000 1186.000000 191.650000 ;
      RECT 1169.500000 188.350000 1170.500000 189.650000 ;
      RECT 1169.500000 187.650000 1186.000000 188.350000 ;
      RECT 1169.500000 186.350000 1170.500000 187.650000 ;
      RECT 0.000000 186.350000 1156.500000 189.650000 ;
      RECT 0.000000 185.650000 1170.500000 186.350000 ;
      RECT 1183.500000 184.350000 1186.000000 187.650000 ;
      RECT 1169.500000 184.350000 1170.500000 185.650000 ;
      RECT 1169.500000 183.650000 1186.000000 184.350000 ;
      RECT 1169.500000 182.350000 1170.500000 183.650000 ;
      RECT 0.000000 182.350000 1156.500000 185.650000 ;
      RECT 0.000000 181.650000 1170.500000 182.350000 ;
      RECT 1183.500000 180.350000 1186.000000 183.650000 ;
      RECT 1169.500000 180.350000 1170.500000 181.650000 ;
      RECT 1169.500000 179.650000 1186.000000 180.350000 ;
      RECT 1169.500000 178.350000 1170.500000 179.650000 ;
      RECT 0.000000 178.350000 1156.500000 181.650000 ;
      RECT 0.000000 177.650000 1170.500000 178.350000 ;
      RECT 1183.500000 176.350000 1186.000000 179.650000 ;
      RECT 1169.500000 176.350000 1170.500000 177.650000 ;
      RECT 1169.500000 175.650000 1186.000000 176.350000 ;
      RECT 1169.500000 174.350000 1170.500000 175.650000 ;
      RECT 0.000000 174.350000 1156.500000 177.650000 ;
      RECT 0.000000 173.650000 1170.500000 174.350000 ;
      RECT 1183.500000 172.350000 1186.000000 175.650000 ;
      RECT 1169.500000 172.350000 1170.500000 173.650000 ;
      RECT 1169.500000 171.650000 1186.000000 172.350000 ;
      RECT 1169.500000 170.350000 1170.500000 171.650000 ;
      RECT 0.000000 170.350000 1156.500000 173.650000 ;
      RECT 0.000000 169.650000 1170.500000 170.350000 ;
      RECT 1183.500000 168.350000 1186.000000 171.650000 ;
      RECT 1169.500000 168.350000 1170.500000 169.650000 ;
      RECT 1169.500000 167.650000 1186.000000 168.350000 ;
      RECT 1169.500000 166.350000 1170.500000 167.650000 ;
      RECT 0.000000 166.350000 1156.500000 169.650000 ;
      RECT 0.000000 165.650000 1170.500000 166.350000 ;
      RECT 1183.500000 164.350000 1186.000000 167.650000 ;
      RECT 1169.500000 164.350000 1170.500000 165.650000 ;
      RECT 1169.500000 163.650000 1186.000000 164.350000 ;
      RECT 1169.500000 162.350000 1170.500000 163.650000 ;
      RECT 0.000000 162.350000 1156.500000 165.650000 ;
      RECT 0.000000 161.650000 1170.500000 162.350000 ;
      RECT 1183.500000 160.350000 1186.000000 163.650000 ;
      RECT 1169.500000 160.350000 1170.500000 161.650000 ;
      RECT 1169.500000 159.650000 1186.000000 160.350000 ;
      RECT 1169.500000 158.350000 1170.500000 159.650000 ;
      RECT 0.000000 158.350000 1156.500000 161.650000 ;
      RECT 0.000000 157.650000 1170.500000 158.350000 ;
      RECT 1183.500000 156.350000 1186.000000 159.650000 ;
      RECT 1169.500000 156.350000 1170.500000 157.650000 ;
      RECT 1169.500000 155.650000 1186.000000 156.350000 ;
      RECT 1169.500000 154.350000 1170.500000 155.650000 ;
      RECT 0.000000 154.350000 1156.500000 157.650000 ;
      RECT 0.000000 153.650000 1170.500000 154.350000 ;
      RECT 1183.500000 152.350000 1186.000000 155.650000 ;
      RECT 1169.500000 152.350000 1170.500000 153.650000 ;
      RECT 1169.500000 151.650000 1186.000000 152.350000 ;
      RECT 1169.500000 150.350000 1170.500000 151.650000 ;
      RECT 0.000000 150.350000 1156.500000 153.650000 ;
      RECT 0.000000 149.650000 1170.500000 150.350000 ;
      RECT 1183.500000 148.350000 1186.000000 151.650000 ;
      RECT 1169.500000 148.350000 1170.500000 149.650000 ;
      RECT 1169.500000 147.650000 1186.000000 148.350000 ;
      RECT 1169.500000 146.350000 1170.500000 147.650000 ;
      RECT 0.000000 146.350000 1156.500000 149.650000 ;
      RECT 0.000000 145.650000 1170.500000 146.350000 ;
      RECT 1183.500000 144.350000 1186.000000 147.650000 ;
      RECT 1169.500000 144.350000 1170.500000 145.650000 ;
      RECT 1169.500000 143.650000 1186.000000 144.350000 ;
      RECT 1169.500000 142.350000 1170.500000 143.650000 ;
      RECT 0.000000 142.350000 1156.500000 145.650000 ;
      RECT 0.000000 141.650000 1170.500000 142.350000 ;
      RECT 1183.500000 140.350000 1186.000000 143.650000 ;
      RECT 1169.500000 140.350000 1170.500000 141.650000 ;
      RECT 1169.500000 139.650000 1186.000000 140.350000 ;
      RECT 1169.500000 138.350000 1170.500000 139.650000 ;
      RECT 0.000000 138.350000 1156.500000 141.650000 ;
      RECT 0.000000 137.650000 1170.500000 138.350000 ;
      RECT 1183.500000 136.350000 1186.000000 139.650000 ;
      RECT 1169.500000 136.350000 1170.500000 137.650000 ;
      RECT 1169.500000 135.650000 1186.000000 136.350000 ;
      RECT 0.000000 135.650000 1156.500000 137.650000 ;
      RECT 0.000000 135.170000 1149.500000 135.650000 ;
      RECT 1183.500000 135.165000 1186.000000 135.650000 ;
      RECT 1169.500000 134.350000 1170.500000 135.650000 ;
      RECT 1157.500000 133.650000 1170.500000 134.350000 ;
      RECT 1183.500000 132.350000 1183.980000 135.165000 ;
      RECT 1169.500000 132.350000 1170.500000 133.650000 ;
      RECT 2.020000 132.350000 1149.500000 135.170000 ;
      RECT 2.020000 132.070000 1156.500000 132.350000 ;
      RECT 1169.500000 132.065000 1183.980000 132.350000 ;
      RECT 1169.500000 131.650000 1186.000000 132.065000 ;
      RECT 1169.500000 130.350000 1170.500000 131.650000 ;
      RECT 0.000000 130.350000 1156.500000 132.070000 ;
      RECT 0.000000 129.650000 1170.500000 130.350000 ;
      RECT 1183.500000 129.485000 1186.000000 131.650000 ;
      RECT 1183.500000 128.350000 1183.980000 129.485000 ;
      RECT 1169.500000 128.350000 1170.500000 129.650000 ;
      RECT 1169.500000 127.650000 1183.980000 128.350000 ;
      RECT 1183.500000 126.385000 1183.980000 127.650000 ;
      RECT 1169.500000 126.350000 1170.500000 127.650000 ;
      RECT 0.000000 126.350000 1156.500000 129.650000 ;
      RECT 0.000000 125.650000 1170.500000 126.350000 ;
      RECT 1183.500000 125.525000 1186.000000 126.385000 ;
      RECT 0.000000 124.575000 1156.500000 125.650000 ;
      RECT 1183.500000 124.350000 1183.980000 125.525000 ;
      RECT 1169.500000 124.350000 1170.500000 125.650000 ;
      RECT 1169.500000 123.650000 1183.980000 124.350000 ;
      RECT 1183.500000 122.425000 1183.980000 123.650000 ;
      RECT 1169.500000 122.350000 1170.500000 123.650000 ;
      RECT 2.020000 122.350000 1156.500000 124.575000 ;
      RECT 2.020000 121.650000 1170.500000 122.350000 ;
      RECT 2.020000 121.475000 1156.500000 121.650000 ;
      RECT 0.000000 120.615000 1156.500000 121.475000 ;
      RECT 1183.500000 120.350000 1186.000000 122.425000 ;
      RECT 1169.500000 120.350000 1170.500000 121.650000 ;
      RECT 1169.500000 119.650000 1186.000000 120.350000 ;
      RECT 1169.500000 118.350000 1170.500000 119.650000 ;
      RECT 2.020000 118.350000 1156.500000 120.615000 ;
      RECT 2.020000 117.650000 1170.500000 118.350000 ;
      RECT 2.020000 117.515000 1156.500000 117.650000 ;
      RECT 1183.500000 116.350000 1186.000000 119.650000 ;
      RECT 1169.500000 116.350000 1170.500000 117.650000 ;
      RECT 1169.500000 115.650000 1186.000000 116.350000 ;
      RECT 0.000000 114.935000 1156.500000 117.515000 ;
      RECT 1183.500000 114.930000 1186.000000 115.650000 ;
      RECT 1169.500000 114.350000 1170.500000 115.650000 ;
      RECT 2.020000 114.350000 1156.500000 114.935000 ;
      RECT 2.020000 113.650000 1170.500000 114.350000 ;
      RECT 1183.500000 112.350000 1183.980000 114.930000 ;
      RECT 1169.500000 112.350000 1170.500000 113.650000 ;
      RECT 2.020000 111.835000 1156.500000 113.650000 ;
      RECT 1169.500000 111.830000 1183.980000 112.350000 ;
      RECT 1169.500000 111.650000 1186.000000 111.830000 ;
      RECT 1169.500000 110.350000 1170.500000 111.650000 ;
      RECT 0.000000 110.350000 1156.500000 111.835000 ;
      RECT 0.000000 109.650000 1170.500000 110.350000 ;
      RECT 1183.500000 108.350000 1186.000000 111.650000 ;
      RECT 1169.500000 108.350000 1170.500000 109.650000 ;
      RECT 1169.500000 107.650000 1186.000000 108.350000 ;
      RECT 1169.500000 106.350000 1170.500000 107.650000 ;
      RECT 0.000000 106.350000 1156.500000 109.650000 ;
      RECT 0.000000 105.650000 1170.500000 106.350000 ;
      RECT 1183.500000 104.350000 1186.000000 107.650000 ;
      RECT 1169.500000 104.350000 1170.500000 105.650000 ;
      RECT 1169.500000 103.650000 1186.000000 104.350000 ;
      RECT 1169.500000 102.350000 1170.500000 103.650000 ;
      RECT 0.000000 102.350000 1156.500000 105.650000 ;
      RECT 0.000000 101.650000 1170.500000 102.350000 ;
      RECT 1183.500000 100.350000 1186.000000 103.650000 ;
      RECT 1169.500000 100.350000 1170.500000 101.650000 ;
      RECT 1169.500000 99.650000 1186.000000 100.350000 ;
      RECT 1169.500000 98.350000 1170.500000 99.650000 ;
      RECT 0.000000 98.350000 1156.500000 101.650000 ;
      RECT 0.000000 97.650000 1170.500000 98.350000 ;
      RECT 1183.500000 96.350000 1186.000000 99.650000 ;
      RECT 1169.500000 96.350000 1170.500000 97.650000 ;
      RECT 1169.500000 95.650000 1186.000000 96.350000 ;
      RECT 1169.500000 94.350000 1170.500000 95.650000 ;
      RECT 0.000000 94.350000 1156.500000 97.650000 ;
      RECT 0.000000 93.650000 1170.500000 94.350000 ;
      RECT 1183.500000 92.350000 1186.000000 95.650000 ;
      RECT 1169.500000 92.350000 1170.500000 93.650000 ;
      RECT 1169.500000 91.650000 1186.000000 92.350000 ;
      RECT 1169.500000 90.350000 1170.500000 91.650000 ;
      RECT 0.000000 90.350000 1156.500000 93.650000 ;
      RECT 0.000000 89.650000 1170.500000 90.350000 ;
      RECT 1183.500000 88.350000 1186.000000 91.650000 ;
      RECT 1169.500000 88.350000 1170.500000 89.650000 ;
      RECT 1169.500000 87.650000 1186.000000 88.350000 ;
      RECT 1169.500000 86.350000 1170.500000 87.650000 ;
      RECT 0.000000 86.350000 1156.500000 89.650000 ;
      RECT 0.000000 85.650000 1170.500000 86.350000 ;
      RECT 1183.500000 84.350000 1186.000000 87.650000 ;
      RECT 1169.500000 84.350000 1170.500000 85.650000 ;
      RECT 1169.500000 83.650000 1186.000000 84.350000 ;
      RECT 1169.500000 82.350000 1170.500000 83.650000 ;
      RECT 0.000000 82.350000 1156.500000 85.650000 ;
      RECT 0.000000 81.650000 1170.500000 82.350000 ;
      RECT 1183.500000 80.350000 1186.000000 83.650000 ;
      RECT 1169.500000 80.350000 1170.500000 81.650000 ;
      RECT 1169.500000 79.650000 1186.000000 80.350000 ;
      RECT 1169.500000 78.350000 1170.500000 79.650000 ;
      RECT 0.000000 78.350000 1156.500000 81.650000 ;
      RECT 0.000000 77.650000 1170.500000 78.350000 ;
      RECT 1183.500000 76.350000 1186.000000 79.650000 ;
      RECT 1169.500000 76.350000 1170.500000 77.650000 ;
      RECT 1169.500000 75.650000 1186.000000 76.350000 ;
      RECT 1169.500000 74.350000 1170.500000 75.650000 ;
      RECT 0.000000 74.350000 1156.500000 77.650000 ;
      RECT 0.000000 73.650000 1170.500000 74.350000 ;
      RECT 1183.500000 72.350000 1186.000000 75.650000 ;
      RECT 1169.500000 72.350000 1170.500000 73.650000 ;
      RECT 1169.500000 71.650000 1186.000000 72.350000 ;
      RECT 1169.500000 70.350000 1170.500000 71.650000 ;
      RECT 0.000000 70.350000 1156.500000 73.650000 ;
      RECT 0.000000 69.650000 1170.500000 70.350000 ;
      RECT 1183.500000 68.350000 1186.000000 71.650000 ;
      RECT 1169.500000 68.350000 1170.500000 69.650000 ;
      RECT 1169.500000 67.650000 1186.000000 68.350000 ;
      RECT 1169.500000 66.350000 1170.500000 67.650000 ;
      RECT 0.000000 66.350000 1156.500000 69.650000 ;
      RECT 0.000000 65.650000 1170.500000 66.350000 ;
      RECT 1183.500000 64.350000 1186.000000 67.650000 ;
      RECT 1169.500000 64.350000 1170.500000 65.650000 ;
      RECT 1169.500000 63.650000 1186.000000 64.350000 ;
      RECT 1169.500000 62.350000 1170.500000 63.650000 ;
      RECT 0.000000 62.350000 1156.500000 65.650000 ;
      RECT 0.000000 61.650000 1170.500000 62.350000 ;
      RECT 1183.500000 60.350000 1186.000000 63.650000 ;
      RECT 1169.500000 60.350000 1170.500000 61.650000 ;
      RECT 1169.500000 59.650000 1186.000000 60.350000 ;
      RECT 1169.500000 58.350000 1170.500000 59.650000 ;
      RECT 0.000000 58.350000 1156.500000 61.650000 ;
      RECT 0.000000 57.650000 1170.500000 58.350000 ;
      RECT 1183.500000 56.350000 1186.000000 59.650000 ;
      RECT 1169.500000 56.350000 1170.500000 57.650000 ;
      RECT 1169.500000 55.650000 1186.000000 56.350000 ;
      RECT 1169.500000 54.350000 1170.500000 55.650000 ;
      RECT 0.000000 54.350000 1156.500000 57.650000 ;
      RECT 0.000000 53.650000 1170.500000 54.350000 ;
      RECT 1183.500000 52.350000 1186.000000 55.650000 ;
      RECT 1169.500000 52.350000 1170.500000 53.650000 ;
      RECT 1169.500000 51.650000 1186.000000 52.350000 ;
      RECT 1169.500000 50.350000 1170.500000 51.650000 ;
      RECT 0.000000 50.350000 1156.500000 53.650000 ;
      RECT 0.000000 49.650000 1170.500000 50.350000 ;
      RECT 1183.500000 48.350000 1186.000000 51.650000 ;
      RECT 1169.500000 48.350000 1170.500000 49.650000 ;
      RECT 1169.500000 47.650000 1186.000000 48.350000 ;
      RECT 0.000000 47.170000 1156.500000 49.650000 ;
      RECT 1183.500000 47.165000 1186.000000 47.650000 ;
      RECT 1169.500000 46.350000 1170.500000 47.650000 ;
      RECT 2.020000 46.350000 1156.500000 47.170000 ;
      RECT 2.020000 45.650000 1170.500000 46.350000 ;
      RECT 1183.500000 44.350000 1183.980000 47.165000 ;
      RECT 1169.500000 44.350000 1170.500000 45.650000 ;
      RECT 2.020000 44.070000 1156.500000 45.650000 ;
      RECT 1169.500000 44.065000 1183.980000 44.350000 ;
      RECT 1169.500000 43.650000 1186.000000 44.065000 ;
      RECT 1169.500000 42.350000 1170.500000 43.650000 ;
      RECT 0.000000 42.350000 1156.500000 44.070000 ;
      RECT 0.000000 41.650000 1170.500000 42.350000 ;
      RECT 1183.500000 41.485000 1186.000000 43.650000 ;
      RECT 1183.500000 40.350000 1183.980000 41.485000 ;
      RECT 1169.500000 40.350000 1170.500000 41.650000 ;
      RECT 1169.500000 39.650000 1183.980000 40.350000 ;
      RECT 1183.500000 38.385000 1183.980000 39.650000 ;
      RECT 1169.500000 38.350000 1170.500000 39.650000 ;
      RECT 0.000000 38.350000 1156.500000 41.650000 ;
      RECT 0.000000 37.650000 1170.500000 38.350000 ;
      RECT 1183.500000 37.525000 1186.000000 38.385000 ;
      RECT 0.000000 36.575000 1156.500000 37.650000 ;
      RECT 1183.500000 36.350000 1183.980000 37.525000 ;
      RECT 1169.500000 36.350000 1170.500000 37.650000 ;
      RECT 1169.500000 35.650000 1183.980000 36.350000 ;
      RECT 1183.500000 34.425000 1183.980000 35.650000 ;
      RECT 1169.500000 34.350000 1170.500000 35.650000 ;
      RECT 2.020000 34.350000 1156.500000 36.575000 ;
      RECT 2.020000 33.650000 1170.500000 34.350000 ;
      RECT 2.020000 33.475000 1156.500000 33.650000 ;
      RECT 0.000000 32.615000 1156.500000 33.475000 ;
      RECT 1183.500000 32.350000 1186.000000 34.425000 ;
      RECT 1169.500000 32.350000 1170.500000 33.650000 ;
      RECT 1169.500000 31.650000 1186.000000 32.350000 ;
      RECT 1169.500000 30.350000 1170.500000 31.650000 ;
      RECT 2.020000 30.350000 1156.500000 32.615000 ;
      RECT 2.020000 29.650000 1170.500000 30.350000 ;
      RECT 2.020000 29.515000 1156.500000 29.650000 ;
      RECT 1183.500000 28.350000 1186.000000 31.650000 ;
      RECT 1169.500000 28.350000 1170.500000 29.650000 ;
      RECT 1169.500000 27.650000 1186.000000 28.350000 ;
      RECT 0.000000 26.935000 1156.500000 29.515000 ;
      RECT 1183.500000 26.930000 1186.000000 27.650000 ;
      RECT 1169.500000 26.350000 1170.500000 27.650000 ;
      RECT 2.020000 26.350000 1156.500000 26.935000 ;
      RECT 2.020000 25.650000 1170.500000 26.350000 ;
      RECT 1183.500000 24.350000 1183.980000 26.930000 ;
      RECT 1169.500000 24.350000 1170.500000 25.650000 ;
      RECT 2.020000 23.835000 1156.500000 25.650000 ;
      RECT 1169.500000 23.830000 1183.980000 24.350000 ;
      RECT 1169.500000 23.650000 1186.000000 23.830000 ;
      RECT 1169.500000 22.350000 1170.500000 23.650000 ;
      RECT 0.000000 22.350000 1156.500000 23.835000 ;
      RECT 0.000000 21.650000 1170.500000 22.350000 ;
      RECT 1183.500000 20.350000 1186.000000 23.650000 ;
      RECT 1169.500000 20.350000 1170.500000 21.650000 ;
      RECT 1169.500000 19.650000 1186.000000 20.350000 ;
      RECT 1169.500000 18.350000 1170.500000 19.650000 ;
      RECT 0.000000 18.350000 1156.500000 21.650000 ;
      RECT 0.000000 17.650000 1170.500000 18.350000 ;
      RECT 1183.500000 16.350000 1186.000000 19.650000 ;
      RECT 1166.500000 16.350000 1170.500000 17.650000 ;
      RECT 1166.500000 15.650000 1186.000000 16.350000 ;
      RECT 1166.500000 14.350000 1170.500000 15.650000 ;
      RECT 0.000000 14.350000 1158.500000 17.650000 ;
      RECT 0.000000 13.650000 1170.500000 14.350000 ;
      RECT 1183.500000 12.350000 1186.000000 15.650000 ;
      RECT 1166.500000 12.350000 1170.500000 13.650000 ;
      RECT 1166.500000 11.650000 1186.000000 12.350000 ;
      RECT 1166.500000 10.350000 1170.500000 11.650000 ;
      RECT 0.000000 10.350000 1158.500000 13.650000 ;
      RECT 0.000000 9.650000 1170.500000 10.350000 ;
      RECT 1183.500000 8.350000 1186.000000 11.650000 ;
      RECT 1166.500000 8.350000 1170.500000 9.650000 ;
      RECT 1166.500000 7.650000 1186.000000 8.350000 ;
      RECT 1116.500000 7.650000 1158.500000 9.650000 ;
      RECT 1066.500000 7.650000 1108.500000 9.650000 ;
      RECT 1016.500000 7.650000 1058.500000 9.650000 ;
      RECT 966.500000 7.650000 1008.500000 9.650000 ;
      RECT 916.500000 7.650000 958.500000 9.650000 ;
      RECT 866.500000 7.650000 908.500000 9.650000 ;
      RECT 816.500000 7.650000 858.500000 9.650000 ;
      RECT 766.500000 7.650000 808.500000 9.650000 ;
      RECT 716.500000 7.650000 758.500000 9.650000 ;
      RECT 666.500000 7.650000 708.500000 9.650000 ;
      RECT 616.500000 7.650000 658.500000 9.650000 ;
      RECT 566.500000 7.650000 608.500000 9.650000 ;
      RECT 516.500000 7.650000 558.500000 9.650000 ;
      RECT 466.500000 7.650000 508.500000 9.650000 ;
      RECT 416.500000 7.650000 458.500000 9.650000 ;
      RECT 366.500000 7.650000 408.500000 9.650000 ;
      RECT 316.500000 7.650000 358.500000 9.650000 ;
      RECT 266.500000 7.650000 308.500000 9.650000 ;
      RECT 216.500000 7.650000 258.500000 9.650000 ;
      RECT 166.500000 7.650000 208.500000 9.650000 ;
      RECT 116.500000 7.650000 158.500000 9.650000 ;
      RECT 66.500000 7.650000 108.500000 9.650000 ;
      RECT 0.000000 7.650000 58.500000 9.650000 ;
      RECT 1166.500000 6.350000 1170.500000 7.650000 ;
      RECT 1157.500000 6.350000 1158.500000 7.650000 ;
      RECT 1116.500000 6.350000 1149.500000 7.650000 ;
      RECT 1107.500000 6.350000 1108.500000 7.650000 ;
      RECT 1066.500000 6.350000 1099.500000 7.650000 ;
      RECT 1057.500000 6.350000 1058.500000 7.650000 ;
      RECT 1016.500000 6.350000 1049.500000 7.650000 ;
      RECT 1007.500000 6.350000 1008.500000 7.650000 ;
      RECT 966.500000 6.350000 999.500000 7.650000 ;
      RECT 957.500000 6.350000 958.500000 7.650000 ;
      RECT 916.500000 6.350000 949.500000 7.650000 ;
      RECT 907.500000 6.350000 908.500000 7.650000 ;
      RECT 866.500000 6.350000 899.500000 7.650000 ;
      RECT 857.500000 6.350000 858.500000 7.650000 ;
      RECT 816.500000 6.350000 849.500000 7.650000 ;
      RECT 807.500000 6.350000 808.500000 7.650000 ;
      RECT 766.500000 6.350000 799.500000 7.650000 ;
      RECT 757.500000 6.350000 758.500000 7.650000 ;
      RECT 716.500000 6.350000 749.500000 7.650000 ;
      RECT 707.500000 6.350000 708.500000 7.650000 ;
      RECT 666.500000 6.350000 699.500000 7.650000 ;
      RECT 657.500000 6.350000 658.500000 7.650000 ;
      RECT 616.500000 6.350000 649.500000 7.650000 ;
      RECT 607.500000 6.350000 608.500000 7.650000 ;
      RECT 566.500000 6.350000 599.500000 7.650000 ;
      RECT 557.500000 6.350000 558.500000 7.650000 ;
      RECT 516.500000 6.350000 549.500000 7.650000 ;
      RECT 507.500000 6.350000 508.500000 7.650000 ;
      RECT 466.500000 6.350000 499.500000 7.650000 ;
      RECT 457.500000 6.350000 458.500000 7.650000 ;
      RECT 416.500000 6.350000 449.500000 7.650000 ;
      RECT 407.500000 6.350000 408.500000 7.650000 ;
      RECT 366.500000 6.350000 399.500000 7.650000 ;
      RECT 357.500000 6.350000 358.500000 7.650000 ;
      RECT 316.500000 6.350000 349.500000 7.650000 ;
      RECT 307.500000 6.350000 308.500000 7.650000 ;
      RECT 266.500000 6.350000 299.500000 7.650000 ;
      RECT 257.500000 6.350000 258.500000 7.650000 ;
      RECT 216.500000 6.350000 249.500000 7.650000 ;
      RECT 207.500000 6.350000 208.500000 7.650000 ;
      RECT 166.500000 6.350000 199.500000 7.650000 ;
      RECT 157.500000 6.350000 158.500000 7.650000 ;
      RECT 116.500000 6.350000 149.500000 7.650000 ;
      RECT 107.500000 6.350000 108.500000 7.650000 ;
      RECT 66.500000 6.350000 99.500000 7.650000 ;
      RECT 57.500000 6.350000 58.500000 7.650000 ;
      RECT 1157.500000 5.650000 1170.500000 6.350000 ;
      RECT 1107.500000 5.650000 1149.500000 6.350000 ;
      RECT 1057.500000 5.650000 1099.500000 6.350000 ;
      RECT 1007.500000 5.650000 1049.500000 6.350000 ;
      RECT 957.500000 5.650000 999.500000 6.350000 ;
      RECT 907.500000 5.650000 949.500000 6.350000 ;
      RECT 857.500000 5.650000 899.500000 6.350000 ;
      RECT 807.500000 5.650000 849.500000 6.350000 ;
      RECT 757.500000 5.650000 799.500000 6.350000 ;
      RECT 707.500000 5.650000 749.500000 6.350000 ;
      RECT 657.500000 5.650000 699.500000 6.350000 ;
      RECT 607.500000 5.650000 649.500000 6.350000 ;
      RECT 557.500000 5.650000 599.500000 6.350000 ;
      RECT 507.500000 5.650000 549.500000 6.350000 ;
      RECT 457.500000 5.650000 499.500000 6.350000 ;
      RECT 407.500000 5.650000 449.500000 6.350000 ;
      RECT 357.500000 5.650000 399.500000 6.350000 ;
      RECT 307.500000 5.650000 349.500000 6.350000 ;
      RECT 257.500000 5.650000 299.500000 6.350000 ;
      RECT 207.500000 5.650000 249.500000 6.350000 ;
      RECT 157.500000 5.650000 199.500000 6.350000 ;
      RECT 107.500000 5.650000 149.500000 6.350000 ;
      RECT 57.500000 5.650000 99.500000 6.350000 ;
      RECT 1183.500000 4.350000 1186.000000 7.650000 ;
      RECT 1166.500000 4.350000 1170.500000 5.650000 ;
      RECT 1157.500000 4.350000 1158.500000 5.650000 ;
      RECT 1116.500000 4.350000 1149.500000 5.650000 ;
      RECT 1107.500000 4.350000 1108.500000 5.650000 ;
      RECT 1066.500000 4.350000 1099.500000 5.650000 ;
      RECT 1057.500000 4.350000 1058.500000 5.650000 ;
      RECT 1016.500000 4.350000 1049.500000 5.650000 ;
      RECT 1007.500000 4.350000 1008.500000 5.650000 ;
      RECT 966.500000 4.350000 999.500000 5.650000 ;
      RECT 957.500000 4.350000 958.500000 5.650000 ;
      RECT 916.500000 4.350000 949.500000 5.650000 ;
      RECT 907.500000 4.350000 908.500000 5.650000 ;
      RECT 866.500000 4.350000 899.500000 5.650000 ;
      RECT 857.500000 4.350000 858.500000 5.650000 ;
      RECT 816.500000 4.350000 849.500000 5.650000 ;
      RECT 807.500000 4.350000 808.500000 5.650000 ;
      RECT 766.500000 4.350000 799.500000 5.650000 ;
      RECT 757.500000 4.350000 758.500000 5.650000 ;
      RECT 716.500000 4.350000 749.500000 5.650000 ;
      RECT 707.500000 4.350000 708.500000 5.650000 ;
      RECT 666.500000 4.350000 699.500000 5.650000 ;
      RECT 657.500000 4.350000 658.500000 5.650000 ;
      RECT 616.500000 4.350000 649.500000 5.650000 ;
      RECT 607.500000 4.350000 608.500000 5.650000 ;
      RECT 566.500000 4.350000 599.500000 5.650000 ;
      RECT 557.500000 4.350000 558.500000 5.650000 ;
      RECT 516.500000 4.350000 549.500000 5.650000 ;
      RECT 507.500000 4.350000 508.500000 5.650000 ;
      RECT 466.500000 4.350000 499.500000 5.650000 ;
      RECT 457.500000 4.350000 458.500000 5.650000 ;
      RECT 416.500000 4.350000 449.500000 5.650000 ;
      RECT 407.500000 4.350000 408.500000 5.650000 ;
      RECT 366.500000 4.350000 399.500000 5.650000 ;
      RECT 357.500000 4.350000 358.500000 5.650000 ;
      RECT 316.500000 4.350000 349.500000 5.650000 ;
      RECT 307.500000 4.350000 308.500000 5.650000 ;
      RECT 266.500000 4.350000 299.500000 5.650000 ;
      RECT 257.500000 4.350000 258.500000 5.650000 ;
      RECT 216.500000 4.350000 249.500000 5.650000 ;
      RECT 207.500000 4.350000 208.500000 5.650000 ;
      RECT 166.500000 4.350000 199.500000 5.650000 ;
      RECT 157.500000 4.350000 158.500000 5.650000 ;
      RECT 116.500000 4.350000 149.500000 5.650000 ;
      RECT 107.500000 4.350000 108.500000 5.650000 ;
      RECT 66.500000 4.350000 99.500000 5.650000 ;
      RECT 57.500000 4.350000 58.500000 5.650000 ;
      RECT 15.500000 4.350000 49.500000 7.650000 ;
      RECT 0.000000 4.350000 2.500000 7.650000 ;
      RECT 1116.500000 3.650000 1158.500000 4.350000 ;
      RECT 1066.500000 3.650000 1108.500000 4.350000 ;
      RECT 1016.500000 3.650000 1058.500000 4.350000 ;
      RECT 966.500000 3.650000 1008.500000 4.350000 ;
      RECT 916.500000 3.650000 958.500000 4.350000 ;
      RECT 866.500000 3.650000 908.500000 4.350000 ;
      RECT 816.500000 3.650000 858.500000 4.350000 ;
      RECT 766.500000 3.650000 808.500000 4.350000 ;
      RECT 716.500000 3.650000 758.500000 4.350000 ;
      RECT 666.500000 3.650000 708.500000 4.350000 ;
      RECT 616.500000 3.650000 658.500000 4.350000 ;
      RECT 566.500000 3.650000 608.500000 4.350000 ;
      RECT 516.500000 3.650000 558.500000 4.350000 ;
      RECT 466.500000 3.650000 508.500000 4.350000 ;
      RECT 416.500000 3.650000 458.500000 4.350000 ;
      RECT 366.500000 3.650000 408.500000 4.350000 ;
      RECT 316.500000 3.650000 358.500000 4.350000 ;
      RECT 266.500000 3.650000 308.500000 4.350000 ;
      RECT 216.500000 3.650000 258.500000 4.350000 ;
      RECT 166.500000 3.650000 208.500000 4.350000 ;
      RECT 116.500000 3.650000 158.500000 4.350000 ;
      RECT 66.500000 3.650000 108.500000 4.350000 ;
      RECT 0.000000 3.650000 58.500000 4.350000 ;
      RECT 1166.500000 2.350000 1186.000000 4.350000 ;
      RECT 1157.500000 2.350000 1158.500000 3.650000 ;
      RECT 1116.500000 2.350000 1149.500000 3.650000 ;
      RECT 1107.500000 2.350000 1108.500000 3.650000 ;
      RECT 1066.500000 2.350000 1099.500000 3.650000 ;
      RECT 1057.500000 2.350000 1058.500000 3.650000 ;
      RECT 1016.500000 2.350000 1049.500000 3.650000 ;
      RECT 1007.500000 2.350000 1008.500000 3.650000 ;
      RECT 966.500000 2.350000 999.500000 3.650000 ;
      RECT 957.500000 2.350000 958.500000 3.650000 ;
      RECT 916.500000 2.350000 949.500000 3.650000 ;
      RECT 907.500000 2.350000 908.500000 3.650000 ;
      RECT 866.500000 2.350000 899.500000 3.650000 ;
      RECT 857.500000 2.350000 858.500000 3.650000 ;
      RECT 816.500000 2.350000 849.500000 3.650000 ;
      RECT 807.500000 2.350000 808.500000 3.650000 ;
      RECT 766.500000 2.350000 799.500000 3.650000 ;
      RECT 757.500000 2.350000 758.500000 3.650000 ;
      RECT 716.500000 2.350000 749.500000 3.650000 ;
      RECT 707.500000 2.350000 708.500000 3.650000 ;
      RECT 666.500000 2.350000 699.500000 3.650000 ;
      RECT 657.500000 2.350000 658.500000 3.650000 ;
      RECT 616.500000 2.350000 649.500000 3.650000 ;
      RECT 607.500000 2.350000 608.500000 3.650000 ;
      RECT 566.500000 2.350000 599.500000 3.650000 ;
      RECT 557.500000 2.350000 558.500000 3.650000 ;
      RECT 516.500000 2.350000 549.500000 3.650000 ;
      RECT 507.500000 2.350000 508.500000 3.650000 ;
      RECT 466.500000 2.350000 499.500000 3.650000 ;
      RECT 457.500000 2.350000 458.500000 3.650000 ;
      RECT 416.500000 2.350000 449.500000 3.650000 ;
      RECT 407.500000 2.350000 408.500000 3.650000 ;
      RECT 366.500000 2.350000 399.500000 3.650000 ;
      RECT 357.500000 2.350000 358.500000 3.650000 ;
      RECT 316.500000 2.350000 349.500000 3.650000 ;
      RECT 307.500000 2.350000 308.500000 3.650000 ;
      RECT 266.500000 2.350000 299.500000 3.650000 ;
      RECT 257.500000 2.350000 258.500000 3.650000 ;
      RECT 216.500000 2.350000 249.500000 3.650000 ;
      RECT 207.500000 2.350000 208.500000 3.650000 ;
      RECT 166.500000 2.350000 199.500000 3.650000 ;
      RECT 157.500000 2.350000 158.500000 3.650000 ;
      RECT 116.500000 2.350000 149.500000 3.650000 ;
      RECT 107.500000 2.350000 108.500000 3.650000 ;
      RECT 66.500000 2.350000 99.500000 3.650000 ;
      RECT 57.500000 2.350000 58.500000 3.650000 ;
      RECT 857.500000 2.020000 899.500000 2.350000 ;
      RECT 807.500000 2.020000 849.500000 2.350000 ;
      RECT 757.500000 2.020000 799.500000 2.350000 ;
      RECT 707.500000 2.020000 749.500000 2.350000 ;
      RECT 607.500000 2.020000 649.500000 2.350000 ;
      RECT 557.500000 2.020000 599.500000 2.350000 ;
      RECT 507.500000 2.020000 549.500000 2.350000 ;
      RECT 457.500000 2.020000 499.500000 2.350000 ;
      RECT 357.500000 2.020000 399.500000 2.350000 ;
      RECT 257.500000 2.020000 299.500000 2.350000 ;
      RECT 107.500000 2.020000 149.500000 2.350000 ;
      RECT 1157.500000 0.350000 1186.000000 2.350000 ;
      RECT 1107.500000 0.350000 1149.500000 2.350000 ;
      RECT 1057.500000 0.350000 1099.500000 2.350000 ;
      RECT 1007.500000 0.350000 1049.500000 2.350000 ;
      RECT 957.500000 0.350000 999.500000 2.350000 ;
      RECT 907.500000 0.350000 949.500000 2.350000 ;
      RECT 899.485000 0.350000 899.500000 2.020000 ;
      RECT 857.500000 0.350000 881.830000 2.020000 ;
      RECT 819.365000 0.350000 849.500000 2.020000 ;
      RECT 799.130000 0.350000 799.500000 2.020000 ;
      RECT 757.500000 0.350000 796.030000 2.020000 ;
      RECT 733.565000 0.350000 749.500000 2.020000 ;
      RECT 707.500000 0.350000 710.230000 2.020000 ;
      RECT 657.500000 0.350000 699.500000 2.350000 ;
      RECT 647.765000 0.350000 649.500000 2.020000 ;
      RECT 607.500000 0.350000 624.430000 2.020000 ;
      RECT 561.965000 0.350000 599.500000 2.020000 ;
      RECT 557.500000 0.350000 558.865000 2.020000 ;
      RECT 507.500000 0.350000 538.630000 2.020000 ;
      RECT 476.165000 0.350000 499.500000 2.020000 ;
      RECT 457.500000 0.350000 463.425000 2.020000 ;
      RECT 407.500000 0.350000 449.500000 2.350000 ;
      RECT 390.365000 0.350000 399.500000 2.020000 ;
      RECT 357.500000 0.350000 367.030000 2.020000 ;
      RECT 307.500000 0.350000 349.500000 2.350000 ;
      RECT 298.885000 0.350000 299.500000 2.020000 ;
      RECT 257.500000 0.350000 281.230000 2.020000 ;
      RECT 207.500000 0.350000 249.500000 2.350000 ;
      RECT 157.500000 0.350000 199.500000 2.350000 ;
      RECT 132.965000 0.350000 149.500000 2.020000 ;
      RECT 107.500000 0.350000 109.630000 2.020000 ;
      RECT 57.500000 0.350000 99.500000 2.350000 ;
      RECT 0.000000 0.350000 49.500000 3.650000 ;
      RECT 905.165000 0.000000 1186.000000 0.350000 ;
      RECT 899.485000 0.000000 902.065000 0.350000 ;
      RECT 895.525000 0.000000 896.385000 2.020000 ;
      RECT 884.930000 0.000000 892.425000 2.020000 ;
      RECT 819.365000 0.000000 881.830000 0.350000 ;
      RECT 813.685000 0.000000 816.265000 2.020000 ;
      RECT 809.725000 0.000000 810.585000 2.020000 ;
      RECT 799.130000 0.000000 806.625000 0.350000 ;
      RECT 733.565000 0.000000 796.030000 0.350000 ;
      RECT 727.885000 0.000000 730.465000 2.020000 ;
      RECT 723.925000 0.000000 724.785000 2.020000 ;
      RECT 713.330000 0.000000 720.825000 2.020000 ;
      RECT 647.765000 0.000000 710.230000 0.350000 ;
      RECT 642.085000 0.000000 644.665000 2.020000 ;
      RECT 638.125000 0.000000 638.985000 2.020000 ;
      RECT 627.530000 0.000000 635.025000 2.020000 ;
      RECT 561.965000 0.000000 624.430000 0.350000 ;
      RECT 556.285000 0.000000 558.865000 0.350000 ;
      RECT 552.325000 0.000000 553.185000 0.350000 ;
      RECT 541.730000 0.000000 549.225000 2.020000 ;
      RECT 476.165000 0.000000 538.630000 0.350000 ;
      RECT 470.485000 0.000000 473.065000 2.020000 ;
      RECT 466.525000 0.000000 467.385000 2.020000 ;
      RECT 455.930000 0.000000 463.425000 0.350000 ;
      RECT 390.365000 0.000000 452.830000 0.350000 ;
      RECT 384.685000 0.000000 387.265000 2.020000 ;
      RECT 380.725000 0.000000 381.585000 2.020000 ;
      RECT 370.130000 0.000000 377.625000 2.020000 ;
      RECT 304.565000 0.000000 367.030000 0.350000 ;
      RECT 298.885000 0.000000 301.465000 0.350000 ;
      RECT 294.925000 0.000000 295.785000 2.020000 ;
      RECT 284.330000 0.000000 291.825000 2.020000 ;
      RECT 132.965000 0.000000 281.230000 0.350000 ;
      RECT 127.285000 0.000000 129.865000 2.020000 ;
      RECT 123.325000 0.000000 124.185000 2.020000 ;
      RECT 112.730000 0.000000 120.225000 2.020000 ;
      RECT 0.000000 0.000000 109.630000 0.350000 ;
    LAYER M3 ;
      RECT 1139.000000 685.650000 1186.000000 686.000000 ;
      RECT 0.000000 685.650000 670.000000 686.000000 ;
      RECT 1139.000000 683.650000 1158.500000 685.650000 ;
      RECT 616.500000 683.650000 658.500000 685.650000 ;
      RECT 566.500000 683.650000 608.500000 685.650000 ;
      RECT 516.500000 683.650000 558.500000 685.650000 ;
      RECT 466.500000 683.650000 508.500000 685.650000 ;
      RECT 416.500000 683.650000 458.500000 685.650000 ;
      RECT 366.500000 683.650000 408.500000 685.650000 ;
      RECT 316.500000 683.650000 358.500000 685.650000 ;
      RECT 0.000000 683.650000 308.500000 685.650000 ;
      RECT 1166.500000 682.350000 1186.000000 685.650000 ;
      RECT 1157.500000 682.350000 1158.500000 683.650000 ;
      RECT 666.500000 682.350000 670.000000 685.650000 ;
      RECT 657.500000 682.350000 658.500000 683.650000 ;
      RECT 616.500000 682.350000 649.500000 683.650000 ;
      RECT 607.500000 682.350000 608.500000 683.650000 ;
      RECT 566.500000 682.350000 599.500000 683.650000 ;
      RECT 557.500000 682.350000 558.500000 683.650000 ;
      RECT 516.500000 682.350000 549.500000 683.650000 ;
      RECT 507.500000 682.350000 508.500000 683.650000 ;
      RECT 466.500000 682.350000 499.500000 683.650000 ;
      RECT 457.500000 682.350000 458.500000 683.650000 ;
      RECT 416.500000 682.350000 449.500000 683.650000 ;
      RECT 407.500000 682.350000 408.500000 683.650000 ;
      RECT 366.500000 682.350000 373.500000 683.650000 ;
      RECT 357.500000 682.350000 358.500000 683.650000 ;
      RECT 316.500000 682.350000 349.500000 683.650000 ;
      RECT 307.500000 682.350000 308.500000 683.650000 ;
      RECT 1157.500000 681.650000 1186.000000 682.350000 ;
      RECT 657.500000 681.650000 670.000000 682.350000 ;
      RECT 607.500000 681.650000 649.500000 682.350000 ;
      RECT 557.500000 681.650000 599.500000 682.350000 ;
      RECT 507.500000 681.650000 549.500000 682.350000 ;
      RECT 457.500000 681.650000 499.500000 682.350000 ;
      RECT 407.500000 681.650000 449.500000 682.350000 ;
      RECT 357.500000 681.650000 373.500000 682.350000 ;
      RECT 307.500000 681.650000 349.500000 682.350000 ;
      RECT 1157.500000 680.350000 1158.500000 681.650000 ;
      RECT 1139.000000 680.350000 1149.500000 683.650000 ;
      RECT 657.500000 680.350000 658.500000 681.650000 ;
      RECT 616.500000 680.350000 649.500000 681.650000 ;
      RECT 607.500000 680.350000 608.500000 681.650000 ;
      RECT 566.500000 680.350000 599.500000 681.650000 ;
      RECT 557.500000 680.350000 558.500000 681.650000 ;
      RECT 516.500000 680.350000 549.500000 681.650000 ;
      RECT 507.500000 680.350000 508.500000 681.650000 ;
      RECT 466.500000 680.350000 499.500000 681.650000 ;
      RECT 457.500000 680.350000 458.500000 681.650000 ;
      RECT 416.500000 680.350000 449.500000 681.650000 ;
      RECT 407.500000 680.350000 408.500000 681.650000 ;
      RECT 386.500000 680.350000 399.500000 683.650000 ;
      RECT 366.500000 680.350000 373.500000 681.650000 ;
      RECT 357.500000 680.350000 358.500000 681.650000 ;
      RECT 316.500000 680.350000 349.500000 681.650000 ;
      RECT 307.500000 680.350000 308.500000 681.650000 ;
      RECT 0.000000 680.350000 299.500000 683.650000 ;
      RECT 1139.000000 679.650000 1158.500000 680.350000 ;
      RECT 616.500000 679.650000 658.500000 680.350000 ;
      RECT 566.500000 679.650000 608.500000 680.350000 ;
      RECT 516.500000 679.650000 558.500000 680.350000 ;
      RECT 466.500000 679.650000 508.500000 680.350000 ;
      RECT 416.500000 679.650000 458.500000 680.350000 ;
      RECT 366.500000 679.650000 408.500000 680.350000 ;
      RECT 316.500000 679.650000 358.500000 680.350000 ;
      RECT 0.000000 679.650000 308.500000 680.350000 ;
      RECT 1166.500000 678.350000 1186.000000 681.650000 ;
      RECT 1157.500000 678.350000 1158.500000 679.650000 ;
      RECT 666.500000 678.350000 670.000000 681.650000 ;
      RECT 657.500000 678.350000 658.500000 679.650000 ;
      RECT 616.500000 678.350000 649.500000 679.650000 ;
      RECT 607.500000 678.350000 608.500000 679.650000 ;
      RECT 566.500000 678.350000 599.500000 679.650000 ;
      RECT 557.500000 678.350000 558.500000 679.650000 ;
      RECT 516.500000 678.350000 549.500000 679.650000 ;
      RECT 507.500000 678.350000 508.500000 679.650000 ;
      RECT 466.500000 678.350000 499.500000 679.650000 ;
      RECT 457.500000 678.350000 458.500000 679.650000 ;
      RECT 416.500000 678.350000 449.500000 679.650000 ;
      RECT 407.500000 678.350000 408.500000 679.650000 ;
      RECT 366.500000 678.350000 373.500000 679.650000 ;
      RECT 357.500000 678.350000 358.500000 679.650000 ;
      RECT 316.500000 678.350000 349.500000 679.650000 ;
      RECT 307.500000 678.350000 308.500000 679.650000 ;
      RECT 1157.500000 677.650000 1186.000000 678.350000 ;
      RECT 657.500000 677.650000 670.000000 678.350000 ;
      RECT 607.500000 677.650000 649.500000 678.350000 ;
      RECT 557.500000 677.650000 599.500000 678.350000 ;
      RECT 507.500000 677.650000 549.500000 678.350000 ;
      RECT 457.500000 677.650000 499.500000 678.350000 ;
      RECT 407.500000 677.650000 449.500000 678.350000 ;
      RECT 357.500000 677.650000 373.500000 678.350000 ;
      RECT 1157.500000 676.350000 1158.500000 677.650000 ;
      RECT 1139.000000 676.350000 1149.500000 679.650000 ;
      RECT 657.500000 676.350000 658.500000 677.650000 ;
      RECT 616.500000 676.350000 649.500000 677.650000 ;
      RECT 607.500000 676.350000 608.500000 677.650000 ;
      RECT 566.500000 676.350000 599.500000 677.650000 ;
      RECT 557.500000 676.350000 558.500000 677.650000 ;
      RECT 516.500000 676.350000 549.500000 677.650000 ;
      RECT 507.500000 676.350000 508.500000 677.650000 ;
      RECT 466.500000 676.350000 499.500000 677.650000 ;
      RECT 457.500000 676.350000 458.500000 677.650000 ;
      RECT 416.500000 676.350000 449.500000 677.650000 ;
      RECT 407.500000 676.350000 408.500000 677.650000 ;
      RECT 386.500000 676.350000 399.500000 679.650000 ;
      RECT 366.500000 676.350000 373.500000 677.650000 ;
      RECT 357.500000 676.350000 358.500000 677.650000 ;
      RECT 307.500000 676.350000 349.500000 678.350000 ;
      RECT 0.000000 676.350000 299.500000 679.650000 ;
      RECT 1139.000000 675.650000 1158.500000 676.350000 ;
      RECT 616.500000 675.650000 658.500000 676.350000 ;
      RECT 566.500000 675.650000 608.500000 676.350000 ;
      RECT 516.500000 675.650000 558.500000 676.350000 ;
      RECT 466.500000 675.650000 508.500000 676.350000 ;
      RECT 416.500000 675.650000 458.500000 676.350000 ;
      RECT 366.500000 675.650000 408.500000 676.350000 ;
      RECT 0.000000 675.650000 358.500000 676.350000 ;
      RECT 1166.500000 674.350000 1186.000000 677.650000 ;
      RECT 1157.500000 674.350000 1158.500000 675.650000 ;
      RECT 666.500000 674.350000 670.000000 677.650000 ;
      RECT 657.500000 674.350000 658.500000 675.650000 ;
      RECT 616.500000 674.350000 649.500000 675.650000 ;
      RECT 607.500000 674.350000 608.500000 675.650000 ;
      RECT 566.500000 674.350000 599.500000 675.650000 ;
      RECT 557.500000 674.350000 558.500000 675.650000 ;
      RECT 516.500000 674.350000 549.500000 675.650000 ;
      RECT 507.500000 674.350000 508.500000 675.650000 ;
      RECT 466.500000 674.350000 499.500000 675.650000 ;
      RECT 457.500000 674.350000 458.500000 675.650000 ;
      RECT 416.500000 674.350000 449.500000 675.650000 ;
      RECT 407.500000 674.350000 408.500000 675.650000 ;
      RECT 366.500000 674.350000 373.500000 675.650000 ;
      RECT 357.500000 674.350000 358.500000 675.650000 ;
      RECT 1157.500000 673.650000 1186.000000 674.350000 ;
      RECT 657.500000 673.650000 670.000000 674.350000 ;
      RECT 607.500000 673.650000 649.500000 674.350000 ;
      RECT 557.500000 673.650000 599.500000 674.350000 ;
      RECT 507.500000 673.650000 549.500000 674.350000 ;
      RECT 457.500000 673.650000 499.500000 674.350000 ;
      RECT 407.500000 673.650000 449.500000 674.350000 ;
      RECT 357.500000 673.650000 373.500000 674.350000 ;
      RECT 1157.500000 672.350000 1158.500000 673.650000 ;
      RECT 1139.000000 672.350000 1149.500000 675.650000 ;
      RECT 657.500000 672.350000 658.500000 673.650000 ;
      RECT 616.500000 672.350000 649.500000 673.650000 ;
      RECT 607.500000 672.350000 608.500000 673.650000 ;
      RECT 566.500000 672.350000 599.500000 673.650000 ;
      RECT 557.500000 672.350000 558.500000 673.650000 ;
      RECT 516.500000 672.350000 549.500000 673.650000 ;
      RECT 507.500000 672.350000 508.500000 673.650000 ;
      RECT 466.500000 672.350000 499.500000 673.650000 ;
      RECT 457.500000 672.350000 458.500000 673.650000 ;
      RECT 416.500000 672.350000 449.500000 673.650000 ;
      RECT 407.500000 672.350000 408.500000 673.650000 ;
      RECT 386.500000 672.350000 399.500000 675.650000 ;
      RECT 366.500000 672.350000 373.500000 673.650000 ;
      RECT 357.500000 672.350000 358.500000 673.650000 ;
      RECT 0.000000 672.350000 349.500000 675.650000 ;
      RECT 1139.000000 671.650000 1158.500000 672.350000 ;
      RECT 616.500000 671.650000 658.500000 672.350000 ;
      RECT 566.500000 671.650000 608.500000 672.350000 ;
      RECT 516.500000 671.650000 558.500000 672.350000 ;
      RECT 466.500000 671.650000 508.500000 672.350000 ;
      RECT 416.500000 671.650000 458.500000 672.350000 ;
      RECT 366.500000 671.650000 408.500000 672.350000 ;
      RECT 0.000000 671.650000 358.500000 672.350000 ;
      RECT 1166.500000 670.350000 1186.000000 673.650000 ;
      RECT 1157.500000 670.350000 1158.500000 671.650000 ;
      RECT 666.500000 670.350000 670.000000 673.650000 ;
      RECT 657.500000 670.350000 658.500000 671.650000 ;
      RECT 616.500000 670.350000 649.500000 671.650000 ;
      RECT 607.500000 670.350000 608.500000 671.650000 ;
      RECT 566.500000 670.350000 599.500000 671.650000 ;
      RECT 557.500000 670.350000 558.500000 671.650000 ;
      RECT 516.500000 670.350000 549.500000 671.650000 ;
      RECT 507.500000 670.350000 508.500000 671.650000 ;
      RECT 466.500000 670.350000 499.500000 671.650000 ;
      RECT 457.500000 670.350000 458.500000 671.650000 ;
      RECT 416.500000 670.350000 449.500000 671.650000 ;
      RECT 407.500000 670.350000 408.500000 671.650000 ;
      RECT 366.500000 670.350000 373.500000 671.650000 ;
      RECT 357.500000 670.350000 358.500000 671.650000 ;
      RECT 1157.500000 669.650000 1186.000000 670.350000 ;
      RECT 657.500000 669.650000 670.000000 670.350000 ;
      RECT 607.500000 669.650000 649.500000 670.350000 ;
      RECT 557.500000 669.650000 599.500000 670.350000 ;
      RECT 507.500000 669.650000 549.500000 670.350000 ;
      RECT 457.500000 669.650000 499.500000 670.350000 ;
      RECT 407.500000 669.650000 449.500000 670.350000 ;
      RECT 357.500000 669.650000 373.500000 670.350000 ;
      RECT 1157.500000 668.350000 1158.500000 669.650000 ;
      RECT 1139.000000 668.350000 1149.500000 671.650000 ;
      RECT 657.500000 668.350000 658.500000 669.650000 ;
      RECT 616.500000 668.350000 649.500000 669.650000 ;
      RECT 607.500000 668.350000 608.500000 669.650000 ;
      RECT 566.500000 668.350000 599.500000 669.650000 ;
      RECT 557.500000 668.350000 558.500000 669.650000 ;
      RECT 516.500000 668.350000 549.500000 669.650000 ;
      RECT 507.500000 668.350000 508.500000 669.650000 ;
      RECT 466.500000 668.350000 499.500000 669.650000 ;
      RECT 457.500000 668.350000 458.500000 669.650000 ;
      RECT 416.500000 668.350000 449.500000 669.650000 ;
      RECT 407.500000 668.350000 408.500000 669.650000 ;
      RECT 386.500000 668.350000 399.500000 671.650000 ;
      RECT 372.500000 668.350000 373.500000 669.650000 ;
      RECT 357.500000 668.350000 358.500000 669.650000 ;
      RECT 0.000000 668.350000 349.500000 671.650000 ;
      RECT 1139.000000 667.650000 1158.500000 668.350000 ;
      RECT 616.500000 667.650000 658.500000 668.350000 ;
      RECT 566.500000 667.650000 608.500000 668.350000 ;
      RECT 516.500000 667.650000 558.500000 668.350000 ;
      RECT 466.500000 667.650000 508.500000 668.350000 ;
      RECT 416.500000 667.650000 458.500000 668.350000 ;
      RECT 372.500000 667.650000 408.500000 668.350000 ;
      RECT 0.000000 667.650000 358.500000 668.350000 ;
      RECT 1166.500000 666.350000 1186.000000 669.650000 ;
      RECT 1157.500000 666.350000 1158.500000 667.650000 ;
      RECT 666.500000 666.350000 670.000000 669.650000 ;
      RECT 657.500000 666.350000 658.500000 667.650000 ;
      RECT 616.500000 666.350000 649.500000 667.650000 ;
      RECT 607.500000 666.350000 608.500000 667.650000 ;
      RECT 566.500000 666.350000 599.500000 667.650000 ;
      RECT 557.500000 666.350000 558.500000 667.650000 ;
      RECT 516.500000 666.350000 549.500000 667.650000 ;
      RECT 507.500000 666.350000 508.500000 667.650000 ;
      RECT 466.500000 666.350000 499.500000 667.650000 ;
      RECT 457.500000 666.350000 458.500000 667.650000 ;
      RECT 416.500000 666.350000 449.500000 667.650000 ;
      RECT 407.500000 666.350000 408.500000 667.650000 ;
      RECT 372.500000 666.350000 373.500000 667.650000 ;
      RECT 357.500000 666.350000 358.500000 667.650000 ;
      RECT 1157.500000 665.650000 1186.000000 666.350000 ;
      RECT 657.500000 665.650000 670.000000 666.350000 ;
      RECT 607.500000 665.650000 649.500000 666.350000 ;
      RECT 557.500000 665.650000 599.500000 666.350000 ;
      RECT 507.500000 665.650000 549.500000 666.350000 ;
      RECT 457.500000 665.650000 499.500000 666.350000 ;
      RECT 407.500000 665.650000 449.500000 666.350000 ;
      RECT 357.500000 665.650000 373.500000 666.350000 ;
      RECT 1157.500000 664.350000 1158.500000 665.650000 ;
      RECT 1139.000000 664.350000 1149.500000 667.650000 ;
      RECT 657.500000 664.350000 658.500000 665.650000 ;
      RECT 616.500000 664.350000 649.500000 665.650000 ;
      RECT 607.500000 664.350000 608.500000 665.650000 ;
      RECT 566.500000 664.350000 599.500000 665.650000 ;
      RECT 557.500000 664.350000 558.500000 665.650000 ;
      RECT 516.500000 664.350000 549.500000 665.650000 ;
      RECT 507.500000 664.350000 508.500000 665.650000 ;
      RECT 466.500000 664.350000 499.500000 665.650000 ;
      RECT 457.500000 664.350000 458.500000 665.650000 ;
      RECT 416.500000 664.350000 449.500000 665.650000 ;
      RECT 407.500000 664.350000 408.500000 665.650000 ;
      RECT 386.500000 664.350000 399.500000 667.650000 ;
      RECT 372.500000 664.350000 373.500000 665.650000 ;
      RECT 357.500000 664.350000 358.500000 665.650000 ;
      RECT 0.000000 664.350000 349.500000 667.650000 ;
      RECT 1139.000000 663.650000 1158.500000 664.350000 ;
      RECT 616.500000 663.650000 658.500000 664.350000 ;
      RECT 566.500000 663.650000 608.500000 664.350000 ;
      RECT 516.500000 663.650000 558.500000 664.350000 ;
      RECT 466.500000 663.650000 508.500000 664.350000 ;
      RECT 416.500000 663.650000 458.500000 664.350000 ;
      RECT 372.500000 663.650000 408.500000 664.350000 ;
      RECT 0.000000 663.650000 358.500000 664.350000 ;
      RECT 1166.500000 662.350000 1186.000000 665.650000 ;
      RECT 1157.500000 662.350000 1158.500000 663.650000 ;
      RECT 666.500000 662.350000 670.000000 665.650000 ;
      RECT 657.500000 662.350000 658.500000 663.650000 ;
      RECT 616.500000 662.350000 649.500000 663.650000 ;
      RECT 607.500000 662.350000 608.500000 663.650000 ;
      RECT 566.500000 662.350000 599.500000 663.650000 ;
      RECT 557.500000 662.350000 558.500000 663.650000 ;
      RECT 516.500000 662.350000 549.500000 663.650000 ;
      RECT 507.500000 662.350000 508.500000 663.650000 ;
      RECT 466.500000 662.350000 499.500000 663.650000 ;
      RECT 457.500000 662.350000 458.500000 663.650000 ;
      RECT 416.500000 662.350000 449.500000 663.650000 ;
      RECT 407.500000 662.350000 408.500000 663.650000 ;
      RECT 372.500000 662.350000 373.500000 663.650000 ;
      RECT 357.500000 662.350000 358.500000 663.650000 ;
      RECT 1157.500000 661.650000 1186.000000 662.350000 ;
      RECT 657.500000 661.650000 670.000000 662.350000 ;
      RECT 607.500000 661.650000 649.500000 662.350000 ;
      RECT 557.500000 661.650000 599.500000 662.350000 ;
      RECT 507.500000 661.650000 549.500000 662.350000 ;
      RECT 457.500000 661.650000 499.500000 662.350000 ;
      RECT 407.500000 661.650000 449.500000 662.350000 ;
      RECT 357.500000 661.650000 373.500000 662.350000 ;
      RECT 1157.500000 660.350000 1158.500000 661.650000 ;
      RECT 1139.000000 660.350000 1149.500000 663.650000 ;
      RECT 657.500000 660.350000 658.500000 661.650000 ;
      RECT 616.500000 660.350000 649.500000 661.650000 ;
      RECT 607.500000 660.350000 608.500000 661.650000 ;
      RECT 566.500000 660.350000 599.500000 661.650000 ;
      RECT 557.500000 660.350000 558.500000 661.650000 ;
      RECT 516.500000 660.350000 549.500000 661.650000 ;
      RECT 507.500000 660.350000 508.500000 661.650000 ;
      RECT 466.500000 660.350000 499.500000 661.650000 ;
      RECT 457.500000 660.350000 458.500000 661.650000 ;
      RECT 416.500000 660.350000 449.500000 661.650000 ;
      RECT 407.500000 660.350000 408.500000 661.650000 ;
      RECT 386.500000 660.350000 399.500000 663.650000 ;
      RECT 372.500000 660.350000 373.500000 661.650000 ;
      RECT 357.500000 660.350000 358.500000 661.650000 ;
      RECT 0.000000 660.350000 349.500000 663.650000 ;
      RECT 1139.000000 659.650000 1158.500000 660.350000 ;
      RECT 616.500000 659.650000 658.500000 660.350000 ;
      RECT 566.500000 659.650000 608.500000 660.350000 ;
      RECT 516.500000 659.650000 558.500000 660.350000 ;
      RECT 466.500000 659.650000 508.500000 660.350000 ;
      RECT 416.500000 659.650000 458.500000 660.350000 ;
      RECT 372.500000 659.650000 408.500000 660.350000 ;
      RECT 0.000000 659.650000 358.500000 660.350000 ;
      RECT 1166.500000 658.350000 1186.000000 661.650000 ;
      RECT 1157.500000 658.350000 1158.500000 659.650000 ;
      RECT 666.500000 658.350000 670.000000 661.650000 ;
      RECT 657.500000 658.350000 658.500000 659.650000 ;
      RECT 616.500000 658.350000 649.500000 659.650000 ;
      RECT 607.500000 658.350000 608.500000 659.650000 ;
      RECT 566.500000 658.350000 599.500000 659.650000 ;
      RECT 557.500000 658.350000 558.500000 659.650000 ;
      RECT 516.500000 658.350000 549.500000 659.650000 ;
      RECT 507.500000 658.350000 508.500000 659.650000 ;
      RECT 466.500000 658.350000 499.500000 659.650000 ;
      RECT 457.500000 658.350000 458.500000 659.650000 ;
      RECT 416.500000 658.350000 449.500000 659.650000 ;
      RECT 407.500000 658.350000 408.500000 659.650000 ;
      RECT 372.500000 658.350000 373.500000 659.650000 ;
      RECT 357.500000 658.350000 358.500000 659.650000 ;
      RECT 1157.500000 657.650000 1186.000000 658.350000 ;
      RECT 357.500000 657.650000 373.500000 658.350000 ;
      RECT 1157.500000 656.350000 1158.500000 657.650000 ;
      RECT 1139.000000 656.350000 1149.500000 659.650000 ;
      RECT 657.500000 656.350000 670.000000 658.350000 ;
      RECT 607.500000 656.350000 649.500000 658.350000 ;
      RECT 557.500000 656.350000 599.500000 658.350000 ;
      RECT 507.500000 656.350000 549.500000 658.350000 ;
      RECT 457.500000 656.350000 499.500000 658.350000 ;
      RECT 407.500000 656.350000 449.500000 658.350000 ;
      RECT 386.500000 656.350000 399.500000 659.650000 ;
      RECT 372.500000 656.350000 373.500000 657.650000 ;
      RECT 357.500000 656.350000 358.500000 657.650000 ;
      RECT 0.000000 656.350000 349.500000 659.650000 ;
      RECT 372.500000 656.000000 670.000000 656.350000 ;
      RECT 1139.000000 655.650000 1158.500000 656.350000 ;
      RECT 372.500000 655.650000 389.000000 656.000000 ;
      RECT 0.000000 655.650000 358.500000 656.350000 ;
      RECT 1166.500000 654.350000 1186.000000 657.650000 ;
      RECT 1157.500000 654.350000 1158.500000 655.650000 ;
      RECT 372.500000 654.350000 373.500000 655.650000 ;
      RECT 357.500000 654.350000 358.500000 655.650000 ;
      RECT 1157.500000 653.650000 1186.000000 654.350000 ;
      RECT 357.500000 653.650000 373.500000 654.350000 ;
      RECT 1157.500000 652.350000 1158.500000 653.650000 ;
      RECT 1139.000000 652.350000 1149.500000 655.650000 ;
      RECT 386.500000 652.350000 389.000000 655.650000 ;
      RECT 372.500000 652.350000 373.500000 653.650000 ;
      RECT 357.500000 652.350000 358.500000 653.650000 ;
      RECT 0.000000 652.350000 349.500000 655.650000 ;
      RECT 1139.000000 651.650000 1158.500000 652.350000 ;
      RECT 372.500000 651.650000 389.000000 652.350000 ;
      RECT 0.000000 651.650000 358.500000 652.350000 ;
      RECT 1166.500000 650.350000 1186.000000 653.650000 ;
      RECT 1157.500000 650.350000 1158.500000 651.650000 ;
      RECT 372.500000 650.350000 373.500000 651.650000 ;
      RECT 357.500000 650.350000 358.500000 651.650000 ;
      RECT 1157.500000 649.650000 1186.000000 650.350000 ;
      RECT 357.500000 649.650000 373.500000 650.350000 ;
      RECT 1157.500000 648.350000 1158.500000 649.650000 ;
      RECT 1139.000000 648.350000 1149.500000 651.650000 ;
      RECT 386.500000 648.350000 389.000000 651.650000 ;
      RECT 372.500000 648.350000 373.500000 649.650000 ;
      RECT 357.500000 648.350000 358.500000 649.650000 ;
      RECT 0.000000 648.350000 349.500000 651.650000 ;
      RECT 1139.000000 647.650000 1158.500000 648.350000 ;
      RECT 372.500000 647.650000 389.000000 648.350000 ;
      RECT 0.000000 647.650000 358.500000 648.350000 ;
      RECT 1166.500000 646.350000 1186.000000 649.650000 ;
      RECT 1157.500000 646.350000 1158.500000 647.650000 ;
      RECT 372.500000 646.350000 373.500000 647.650000 ;
      RECT 357.500000 646.350000 358.500000 647.650000 ;
      RECT 1157.500000 645.650000 1186.000000 646.350000 ;
      RECT 357.500000 645.650000 373.500000 646.350000 ;
      RECT 1157.500000 644.350000 1158.500000 645.650000 ;
      RECT 1139.000000 644.350000 1149.500000 647.650000 ;
      RECT 386.500000 644.350000 389.000000 647.650000 ;
      RECT 372.500000 644.350000 373.500000 645.650000 ;
      RECT 357.500000 644.350000 358.500000 645.650000 ;
      RECT 0.000000 644.350000 349.500000 647.650000 ;
      RECT 1139.000000 643.650000 1158.500000 644.350000 ;
      RECT 372.500000 643.650000 389.000000 644.350000 ;
      RECT 0.000000 643.650000 358.500000 644.350000 ;
      RECT 1166.500000 642.350000 1186.000000 645.650000 ;
      RECT 1157.500000 642.350000 1158.500000 643.650000 ;
      RECT 372.500000 642.350000 373.500000 643.650000 ;
      RECT 357.500000 642.350000 358.500000 643.650000 ;
      RECT 1157.500000 641.650000 1186.000000 642.350000 ;
      RECT 357.500000 641.650000 373.500000 642.350000 ;
      RECT 1157.500000 640.350000 1158.500000 641.650000 ;
      RECT 1139.000000 640.350000 1149.500000 643.650000 ;
      RECT 386.500000 640.350000 389.000000 643.650000 ;
      RECT 372.500000 640.350000 373.500000 641.650000 ;
      RECT 357.500000 640.350000 358.500000 641.650000 ;
      RECT 0.000000 640.350000 349.500000 643.650000 ;
      RECT 1139.000000 639.650000 1158.500000 640.350000 ;
      RECT 372.500000 639.650000 389.000000 640.350000 ;
      RECT 0.000000 639.650000 358.500000 640.350000 ;
      RECT 1166.500000 638.350000 1186.000000 641.650000 ;
      RECT 1157.500000 638.350000 1158.500000 639.650000 ;
      RECT 372.500000 638.350000 373.500000 639.650000 ;
      RECT 357.500000 638.350000 358.500000 639.650000 ;
      RECT 1157.500000 637.650000 1186.000000 638.350000 ;
      RECT 357.500000 637.650000 373.500000 638.350000 ;
      RECT 1157.500000 636.350000 1158.500000 637.650000 ;
      RECT 1139.000000 636.350000 1149.500000 639.650000 ;
      RECT 386.500000 636.350000 389.000000 639.650000 ;
      RECT 372.500000 636.350000 373.500000 637.650000 ;
      RECT 357.500000 636.350000 358.500000 637.650000 ;
      RECT 0.000000 636.350000 349.500000 639.650000 ;
      RECT 1139.000000 635.650000 1158.500000 636.350000 ;
      RECT 372.500000 635.650000 389.000000 636.350000 ;
      RECT 0.000000 635.650000 358.500000 636.350000 ;
      RECT 1166.500000 634.350000 1186.000000 637.650000 ;
      RECT 1157.500000 634.350000 1158.500000 635.650000 ;
      RECT 372.500000 634.350000 373.500000 635.650000 ;
      RECT 357.500000 634.350000 358.500000 635.650000 ;
      RECT 1157.500000 633.650000 1186.000000 634.350000 ;
      RECT 357.500000 633.650000 373.500000 634.350000 ;
      RECT 1157.500000 632.350000 1158.500000 633.650000 ;
      RECT 1139.000000 632.350000 1149.500000 635.650000 ;
      RECT 386.500000 632.350000 389.000000 635.650000 ;
      RECT 372.500000 632.350000 373.500000 633.650000 ;
      RECT 357.500000 632.350000 358.500000 633.650000 ;
      RECT 0.000000 632.350000 349.500000 635.650000 ;
      RECT 1139.000000 631.650000 1158.500000 632.350000 ;
      RECT 372.500000 631.650000 389.000000 632.350000 ;
      RECT 0.000000 631.650000 358.500000 632.350000 ;
      RECT 1166.500000 630.350000 1186.000000 633.650000 ;
      RECT 1157.500000 630.350000 1158.500000 631.650000 ;
      RECT 372.500000 630.350000 373.500000 631.650000 ;
      RECT 357.500000 630.350000 358.500000 631.650000 ;
      RECT 1157.500000 629.650000 1186.000000 630.350000 ;
      RECT 357.500000 629.650000 373.500000 630.350000 ;
      RECT 1157.500000 628.350000 1158.500000 629.650000 ;
      RECT 1139.000000 628.350000 1149.500000 631.650000 ;
      RECT 386.500000 628.350000 389.000000 631.650000 ;
      RECT 372.500000 628.350000 373.500000 629.650000 ;
      RECT 357.500000 628.350000 358.500000 629.650000 ;
      RECT 0.000000 628.350000 349.500000 631.650000 ;
      RECT 1139.000000 627.650000 1158.500000 628.350000 ;
      RECT 372.500000 627.650000 389.000000 628.350000 ;
      RECT 0.000000 627.650000 358.500000 628.350000 ;
      RECT 1166.500000 626.350000 1186.000000 629.650000 ;
      RECT 1157.500000 626.350000 1158.500000 627.650000 ;
      RECT 372.500000 626.350000 373.500000 627.650000 ;
      RECT 357.500000 626.350000 358.500000 627.650000 ;
      RECT 1157.500000 625.650000 1186.000000 626.350000 ;
      RECT 357.500000 625.650000 373.500000 626.350000 ;
      RECT 1157.500000 624.350000 1158.500000 625.650000 ;
      RECT 1139.000000 624.350000 1149.500000 627.650000 ;
      RECT 386.500000 624.350000 389.000000 627.650000 ;
      RECT 372.500000 624.350000 373.500000 625.650000 ;
      RECT 357.500000 624.350000 358.500000 625.650000 ;
      RECT 0.000000 624.350000 349.500000 627.650000 ;
      RECT 1139.000000 623.650000 1158.500000 624.350000 ;
      RECT 372.500000 623.650000 389.000000 624.350000 ;
      RECT 0.000000 623.650000 358.500000 624.350000 ;
      RECT 1166.500000 622.350000 1186.000000 625.650000 ;
      RECT 1157.500000 622.350000 1158.500000 623.650000 ;
      RECT 372.500000 622.350000 373.500000 623.650000 ;
      RECT 357.500000 622.350000 358.500000 623.650000 ;
      RECT 1157.500000 621.650000 1186.000000 622.350000 ;
      RECT 357.500000 621.650000 373.500000 622.350000 ;
      RECT 1157.500000 620.350000 1158.500000 621.650000 ;
      RECT 1139.000000 620.350000 1149.500000 623.650000 ;
      RECT 386.500000 620.350000 389.000000 623.650000 ;
      RECT 372.500000 620.350000 373.500000 621.650000 ;
      RECT 357.500000 620.350000 358.500000 621.650000 ;
      RECT 0.000000 620.350000 349.500000 623.650000 ;
      RECT 1139.000000 619.650000 1158.500000 620.350000 ;
      RECT 372.500000 619.650000 389.000000 620.350000 ;
      RECT 0.000000 619.650000 358.500000 620.350000 ;
      RECT 1166.500000 618.350000 1186.000000 621.650000 ;
      RECT 1157.500000 618.350000 1158.500000 619.650000 ;
      RECT 372.500000 618.350000 373.500000 619.650000 ;
      RECT 357.500000 618.350000 358.500000 619.650000 ;
      RECT 1157.500000 617.650000 1186.000000 618.350000 ;
      RECT 357.500000 617.650000 373.500000 618.350000 ;
      RECT 1157.500000 616.350000 1158.500000 617.650000 ;
      RECT 1139.000000 616.350000 1149.500000 619.650000 ;
      RECT 386.500000 616.350000 389.000000 619.650000 ;
      RECT 372.500000 616.350000 373.500000 617.650000 ;
      RECT 357.500000 616.350000 358.500000 617.650000 ;
      RECT 0.000000 616.350000 349.500000 619.650000 ;
      RECT 1139.000000 615.650000 1158.500000 616.350000 ;
      RECT 372.500000 615.650000 389.000000 616.350000 ;
      RECT 0.000000 615.650000 358.500000 616.350000 ;
      RECT 1166.500000 614.350000 1186.000000 617.650000 ;
      RECT 1157.500000 614.350000 1158.500000 615.650000 ;
      RECT 372.500000 614.350000 373.500000 615.650000 ;
      RECT 357.500000 614.350000 358.500000 615.650000 ;
      RECT 1157.500000 613.650000 1186.000000 614.350000 ;
      RECT 357.500000 613.650000 373.500000 614.350000 ;
      RECT 1157.500000 612.350000 1158.500000 613.650000 ;
      RECT 1139.000000 612.350000 1149.500000 615.650000 ;
      RECT 386.500000 612.350000 389.000000 615.650000 ;
      RECT 372.500000 612.350000 373.500000 613.650000 ;
      RECT 357.500000 612.350000 358.500000 613.650000 ;
      RECT 0.000000 612.350000 349.500000 615.650000 ;
      RECT 1139.000000 611.650000 1158.500000 612.350000 ;
      RECT 372.500000 611.650000 389.000000 612.350000 ;
      RECT 0.000000 611.650000 358.500000 612.350000 ;
      RECT 1166.500000 610.350000 1186.000000 613.650000 ;
      RECT 1157.500000 610.350000 1158.500000 611.650000 ;
      RECT 372.500000 610.350000 373.500000 611.650000 ;
      RECT 357.500000 610.350000 358.500000 611.650000 ;
      RECT 1157.500000 609.650000 1186.000000 610.350000 ;
      RECT 357.500000 609.650000 373.500000 610.350000 ;
      RECT 1157.500000 608.350000 1158.500000 609.650000 ;
      RECT 1139.000000 608.350000 1149.500000 611.650000 ;
      RECT 386.500000 608.350000 389.000000 611.650000 ;
      RECT 372.500000 608.350000 373.500000 609.650000 ;
      RECT 357.500000 608.350000 358.500000 609.650000 ;
      RECT 0.000000 608.350000 349.500000 611.650000 ;
      RECT 1139.000000 607.650000 1158.500000 608.350000 ;
      RECT 372.500000 607.650000 389.000000 608.350000 ;
      RECT 0.000000 607.650000 358.500000 608.350000 ;
      RECT 1166.500000 606.350000 1186.000000 609.650000 ;
      RECT 1157.500000 606.350000 1158.500000 607.650000 ;
      RECT 372.500000 606.350000 373.500000 607.650000 ;
      RECT 357.500000 606.350000 358.500000 607.650000 ;
      RECT 1157.500000 605.650000 1186.000000 606.350000 ;
      RECT 357.500000 605.650000 373.500000 606.350000 ;
      RECT 1157.500000 604.350000 1158.500000 605.650000 ;
      RECT 1139.000000 604.350000 1149.500000 607.650000 ;
      RECT 386.500000 604.350000 389.000000 607.650000 ;
      RECT 372.500000 604.350000 373.500000 605.650000 ;
      RECT 357.500000 604.350000 358.500000 605.650000 ;
      RECT 0.000000 604.350000 349.500000 607.650000 ;
      RECT 1139.000000 603.650000 1158.500000 604.350000 ;
      RECT 372.500000 603.650000 389.000000 604.350000 ;
      RECT 0.000000 603.650000 358.500000 604.350000 ;
      RECT 1166.500000 602.350000 1186.000000 605.650000 ;
      RECT 1157.500000 602.350000 1158.500000 603.650000 ;
      RECT 372.500000 602.350000 373.500000 603.650000 ;
      RECT 357.500000 602.350000 358.500000 603.650000 ;
      RECT 1157.500000 601.650000 1186.000000 602.350000 ;
      RECT 357.500000 601.650000 373.500000 602.350000 ;
      RECT 1157.500000 600.350000 1158.500000 601.650000 ;
      RECT 1139.000000 600.350000 1149.500000 603.650000 ;
      RECT 386.500000 600.350000 389.000000 603.650000 ;
      RECT 372.500000 600.350000 373.500000 601.650000 ;
      RECT 357.500000 600.350000 358.500000 601.650000 ;
      RECT 0.000000 600.350000 349.500000 603.650000 ;
      RECT 1139.000000 599.650000 1158.500000 600.350000 ;
      RECT 372.500000 599.650000 389.000000 600.350000 ;
      RECT 0.000000 599.650000 358.500000 600.350000 ;
      RECT 1166.500000 598.350000 1186.000000 601.650000 ;
      RECT 1157.500000 598.350000 1158.500000 599.650000 ;
      RECT 372.500000 598.350000 373.500000 599.650000 ;
      RECT 357.500000 598.350000 358.500000 599.650000 ;
      RECT 1157.500000 597.650000 1186.000000 598.350000 ;
      RECT 357.500000 597.650000 373.500000 598.350000 ;
      RECT 1157.500000 596.350000 1158.500000 597.650000 ;
      RECT 1139.000000 596.350000 1149.500000 599.650000 ;
      RECT 386.500000 596.350000 389.000000 599.650000 ;
      RECT 372.500000 596.350000 373.500000 597.650000 ;
      RECT 357.500000 596.350000 358.500000 597.650000 ;
      RECT 0.000000 596.350000 349.500000 599.650000 ;
      RECT 1139.000000 595.650000 1158.500000 596.350000 ;
      RECT 372.500000 595.650000 389.000000 596.350000 ;
      RECT 0.000000 595.650000 358.500000 596.350000 ;
      RECT 1166.500000 594.350000 1186.000000 597.650000 ;
      RECT 1157.500000 594.350000 1158.500000 595.650000 ;
      RECT 372.500000 594.350000 373.500000 595.650000 ;
      RECT 357.500000 594.350000 358.500000 595.650000 ;
      RECT 1157.500000 593.650000 1186.000000 594.350000 ;
      RECT 357.500000 593.650000 373.500000 594.350000 ;
      RECT 1157.500000 592.350000 1158.500000 593.650000 ;
      RECT 1139.000000 592.350000 1149.500000 595.650000 ;
      RECT 386.500000 592.350000 389.000000 595.650000 ;
      RECT 372.500000 592.350000 373.500000 593.650000 ;
      RECT 357.500000 592.350000 358.500000 593.650000 ;
      RECT 0.000000 592.350000 349.500000 595.650000 ;
      RECT 1139.000000 591.650000 1158.500000 592.350000 ;
      RECT 372.500000 591.650000 389.000000 592.350000 ;
      RECT 0.000000 591.650000 358.500000 592.350000 ;
      RECT 1166.500000 590.350000 1186.000000 593.650000 ;
      RECT 1157.500000 590.350000 1158.500000 591.650000 ;
      RECT 372.500000 590.350000 373.500000 591.650000 ;
      RECT 357.500000 590.350000 358.500000 591.650000 ;
      RECT 1157.500000 589.650000 1186.000000 590.350000 ;
      RECT 357.500000 589.650000 373.500000 590.350000 ;
      RECT 1157.500000 588.350000 1158.500000 589.650000 ;
      RECT 1139.000000 588.350000 1149.500000 591.650000 ;
      RECT 386.500000 588.350000 389.000000 591.650000 ;
      RECT 372.500000 588.350000 373.500000 589.650000 ;
      RECT 357.500000 588.350000 358.500000 589.650000 ;
      RECT 0.000000 588.350000 349.500000 591.650000 ;
      RECT 1139.000000 587.650000 1158.500000 588.350000 ;
      RECT 372.500000 587.650000 389.000000 588.350000 ;
      RECT 0.000000 587.650000 358.500000 588.350000 ;
      RECT 1166.500000 586.350000 1186.000000 589.650000 ;
      RECT 1157.500000 586.350000 1158.500000 587.650000 ;
      RECT 372.500000 586.350000 373.500000 587.650000 ;
      RECT 357.500000 586.350000 358.500000 587.650000 ;
      RECT 1157.500000 585.650000 1186.000000 586.350000 ;
      RECT 357.500000 585.650000 373.500000 586.350000 ;
      RECT 1157.500000 584.350000 1158.500000 585.650000 ;
      RECT 1139.000000 584.350000 1149.500000 587.650000 ;
      RECT 386.500000 584.350000 389.000000 587.650000 ;
      RECT 372.500000 584.350000 373.500000 585.650000 ;
      RECT 357.500000 584.350000 358.500000 585.650000 ;
      RECT 0.000000 584.350000 349.500000 587.650000 ;
      RECT 1139.000000 583.650000 1158.500000 584.350000 ;
      RECT 372.500000 583.650000 389.000000 584.350000 ;
      RECT 0.000000 583.650000 358.500000 584.350000 ;
      RECT 1166.500000 582.350000 1186.000000 585.650000 ;
      RECT 1157.500000 582.350000 1158.500000 583.650000 ;
      RECT 372.500000 582.350000 373.500000 583.650000 ;
      RECT 357.500000 582.350000 358.500000 583.650000 ;
      RECT 1157.500000 581.650000 1186.000000 582.350000 ;
      RECT 357.500000 581.650000 373.500000 582.350000 ;
      RECT 1157.500000 580.350000 1158.500000 581.650000 ;
      RECT 1139.000000 580.350000 1149.500000 583.650000 ;
      RECT 386.500000 580.350000 389.000000 583.650000 ;
      RECT 372.500000 580.350000 373.500000 581.650000 ;
      RECT 357.500000 580.350000 358.500000 581.650000 ;
      RECT 0.000000 580.350000 349.500000 583.650000 ;
      RECT 1139.000000 579.650000 1158.500000 580.350000 ;
      RECT 372.500000 579.650000 389.000000 580.350000 ;
      RECT 0.000000 579.650000 358.500000 580.350000 ;
      RECT 1166.500000 578.350000 1186.000000 581.650000 ;
      RECT 1157.500000 578.350000 1158.500000 579.650000 ;
      RECT 372.500000 578.350000 373.500000 579.650000 ;
      RECT 357.500000 578.350000 358.500000 579.650000 ;
      RECT 1157.500000 577.650000 1186.000000 578.350000 ;
      RECT 357.500000 577.650000 373.500000 578.350000 ;
      RECT 1157.500000 576.350000 1158.500000 577.650000 ;
      RECT 1139.000000 576.350000 1149.500000 579.650000 ;
      RECT 386.500000 576.350000 389.000000 579.650000 ;
      RECT 372.500000 576.350000 373.500000 577.650000 ;
      RECT 357.500000 576.350000 358.500000 577.650000 ;
      RECT 0.000000 576.350000 349.500000 579.650000 ;
      RECT 1139.000000 575.650000 1158.500000 576.350000 ;
      RECT 372.500000 575.650000 389.000000 576.350000 ;
      RECT 0.000000 575.650000 358.500000 576.350000 ;
      RECT 1166.500000 574.350000 1186.000000 577.650000 ;
      RECT 1157.500000 574.350000 1158.500000 575.650000 ;
      RECT 372.500000 574.350000 373.500000 575.650000 ;
      RECT 357.500000 574.350000 358.500000 575.650000 ;
      RECT 1157.500000 573.650000 1186.000000 574.350000 ;
      RECT 357.500000 573.650000 373.500000 574.350000 ;
      RECT 1157.500000 572.350000 1158.500000 573.650000 ;
      RECT 1139.000000 572.350000 1149.500000 575.650000 ;
      RECT 386.500000 572.350000 389.000000 575.650000 ;
      RECT 372.500000 572.350000 373.500000 573.650000 ;
      RECT 357.500000 572.350000 358.500000 573.650000 ;
      RECT 0.000000 572.350000 349.500000 575.650000 ;
      RECT 1139.000000 571.650000 1158.500000 572.350000 ;
      RECT 372.500000 571.650000 389.000000 572.350000 ;
      RECT 0.000000 571.650000 358.500000 572.350000 ;
      RECT 1166.500000 570.350000 1186.000000 573.650000 ;
      RECT 1157.500000 570.350000 1158.500000 571.650000 ;
      RECT 372.500000 570.350000 373.500000 571.650000 ;
      RECT 357.500000 570.350000 358.500000 571.650000 ;
      RECT 1157.500000 569.650000 1186.000000 570.350000 ;
      RECT 357.500000 569.650000 373.500000 570.350000 ;
      RECT 1157.500000 568.350000 1158.500000 569.650000 ;
      RECT 1139.000000 568.350000 1149.500000 571.650000 ;
      RECT 386.500000 568.350000 389.000000 571.650000 ;
      RECT 372.500000 568.350000 373.500000 569.650000 ;
      RECT 357.500000 568.350000 358.500000 569.650000 ;
      RECT 0.000000 568.350000 349.500000 571.650000 ;
      RECT 1139.000000 567.650000 1158.500000 568.350000 ;
      RECT 372.500000 567.650000 389.000000 568.350000 ;
      RECT 0.000000 567.650000 358.500000 568.350000 ;
      RECT 1166.500000 566.350000 1186.000000 569.650000 ;
      RECT 1157.500000 566.350000 1158.500000 567.650000 ;
      RECT 372.500000 566.350000 373.500000 567.650000 ;
      RECT 357.500000 566.350000 358.500000 567.650000 ;
      RECT 1157.500000 565.650000 1186.000000 566.350000 ;
      RECT 357.500000 565.650000 373.500000 566.350000 ;
      RECT 1157.500000 564.350000 1158.500000 565.650000 ;
      RECT 1139.000000 564.350000 1149.500000 567.650000 ;
      RECT 386.500000 564.350000 389.000000 567.650000 ;
      RECT 372.500000 564.350000 373.500000 565.650000 ;
      RECT 357.500000 564.350000 358.500000 565.650000 ;
      RECT 0.000000 564.350000 349.500000 567.650000 ;
      RECT 1139.000000 563.650000 1158.500000 564.350000 ;
      RECT 372.500000 563.650000 389.000000 564.350000 ;
      RECT 0.000000 563.650000 358.500000 564.350000 ;
      RECT 1166.500000 562.350000 1186.000000 565.650000 ;
      RECT 1157.500000 562.350000 1158.500000 563.650000 ;
      RECT 372.500000 562.350000 373.500000 563.650000 ;
      RECT 357.500000 562.350000 358.500000 563.650000 ;
      RECT 1157.500000 561.650000 1186.000000 562.350000 ;
      RECT 357.500000 561.650000 373.500000 562.350000 ;
      RECT 1157.500000 560.350000 1158.500000 561.650000 ;
      RECT 1139.000000 560.350000 1149.500000 563.650000 ;
      RECT 386.500000 560.350000 389.000000 563.650000 ;
      RECT 372.500000 560.350000 373.500000 561.650000 ;
      RECT 357.500000 560.350000 358.500000 561.650000 ;
      RECT 0.000000 560.350000 349.500000 563.650000 ;
      RECT 1139.000000 559.650000 1158.500000 560.350000 ;
      RECT 372.500000 559.650000 389.000000 560.350000 ;
      RECT 0.000000 559.650000 358.500000 560.350000 ;
      RECT 1166.500000 558.350000 1186.000000 561.650000 ;
      RECT 1157.500000 558.350000 1158.500000 559.650000 ;
      RECT 372.500000 558.350000 373.500000 559.650000 ;
      RECT 357.500000 558.350000 358.500000 559.650000 ;
      RECT 1157.500000 557.650000 1186.000000 558.350000 ;
      RECT 357.500000 557.650000 373.500000 558.350000 ;
      RECT 1157.500000 556.350000 1158.500000 557.650000 ;
      RECT 1139.000000 556.350000 1149.500000 559.650000 ;
      RECT 386.500000 556.350000 389.000000 559.650000 ;
      RECT 372.500000 556.350000 373.500000 557.650000 ;
      RECT 357.500000 556.350000 358.500000 557.650000 ;
      RECT 0.000000 556.350000 349.500000 559.650000 ;
      RECT 1139.000000 555.650000 1158.500000 556.350000 ;
      RECT 372.500000 555.650000 389.000000 556.350000 ;
      RECT 0.000000 555.650000 358.500000 556.350000 ;
      RECT 1166.500000 554.350000 1186.000000 557.650000 ;
      RECT 1157.500000 554.350000 1158.500000 555.650000 ;
      RECT 372.500000 554.350000 373.500000 555.650000 ;
      RECT 357.500000 554.350000 358.500000 555.650000 ;
      RECT 1157.500000 553.650000 1186.000000 554.350000 ;
      RECT 357.500000 553.650000 373.500000 554.350000 ;
      RECT 1157.500000 552.350000 1158.500000 553.650000 ;
      RECT 1139.000000 552.350000 1149.500000 555.650000 ;
      RECT 386.500000 552.350000 389.000000 555.650000 ;
      RECT 372.500000 552.350000 373.500000 553.650000 ;
      RECT 357.500000 552.350000 358.500000 553.650000 ;
      RECT 0.000000 552.350000 349.500000 555.650000 ;
      RECT 1139.000000 551.650000 1158.500000 552.350000 ;
      RECT 372.500000 551.650000 389.000000 552.350000 ;
      RECT 0.000000 551.650000 358.500000 552.350000 ;
      RECT 1166.500000 550.350000 1186.000000 553.650000 ;
      RECT 1157.500000 550.350000 1158.500000 551.650000 ;
      RECT 372.500000 550.350000 373.500000 551.650000 ;
      RECT 357.500000 550.350000 358.500000 551.650000 ;
      RECT 1157.500000 549.650000 1186.000000 550.350000 ;
      RECT 357.500000 549.650000 373.500000 550.350000 ;
      RECT 1157.500000 548.350000 1158.500000 549.650000 ;
      RECT 1139.000000 548.350000 1149.500000 551.650000 ;
      RECT 386.500000 548.350000 389.000000 551.650000 ;
      RECT 372.500000 548.350000 373.500000 549.650000 ;
      RECT 357.500000 548.350000 358.500000 549.650000 ;
      RECT 0.000000 548.350000 349.500000 551.650000 ;
      RECT 1139.000000 547.650000 1158.500000 548.350000 ;
      RECT 372.500000 547.650000 389.000000 548.350000 ;
      RECT 0.000000 547.650000 358.500000 548.350000 ;
      RECT 1166.500000 546.350000 1186.000000 549.650000 ;
      RECT 1157.500000 546.350000 1158.500000 547.650000 ;
      RECT 372.500000 546.350000 373.500000 547.650000 ;
      RECT 357.500000 546.350000 358.500000 547.650000 ;
      RECT 1157.500000 545.650000 1186.000000 546.350000 ;
      RECT 357.500000 545.650000 373.500000 546.350000 ;
      RECT 1157.500000 544.350000 1158.500000 545.650000 ;
      RECT 1139.000000 544.350000 1149.500000 547.650000 ;
      RECT 386.500000 544.350000 389.000000 547.650000 ;
      RECT 372.500000 544.350000 373.500000 545.650000 ;
      RECT 357.500000 544.350000 358.500000 545.650000 ;
      RECT 0.000000 544.350000 349.500000 547.650000 ;
      RECT 1139.000000 543.650000 1158.500000 544.350000 ;
      RECT 372.500000 543.650000 389.000000 544.350000 ;
      RECT 0.000000 543.650000 358.500000 544.350000 ;
      RECT 1166.500000 542.350000 1186.000000 545.650000 ;
      RECT 1157.500000 542.350000 1158.500000 543.650000 ;
      RECT 372.500000 542.350000 373.500000 543.650000 ;
      RECT 357.500000 542.350000 358.500000 543.650000 ;
      RECT 1157.500000 541.650000 1186.000000 542.350000 ;
      RECT 357.500000 541.650000 373.500000 542.350000 ;
      RECT 1157.500000 540.350000 1158.500000 541.650000 ;
      RECT 1139.000000 540.350000 1149.500000 543.650000 ;
      RECT 386.500000 540.350000 389.000000 543.650000 ;
      RECT 372.500000 540.350000 373.500000 541.650000 ;
      RECT 357.500000 540.350000 358.500000 541.650000 ;
      RECT 0.000000 540.350000 349.500000 543.650000 ;
      RECT 1139.000000 539.650000 1158.500000 540.350000 ;
      RECT 372.500000 539.650000 389.000000 540.350000 ;
      RECT 0.000000 539.650000 358.500000 540.350000 ;
      RECT 1166.500000 538.350000 1186.000000 541.650000 ;
      RECT 1157.500000 538.350000 1158.500000 539.650000 ;
      RECT 372.500000 538.350000 373.500000 539.650000 ;
      RECT 357.500000 538.350000 358.500000 539.650000 ;
      RECT 1157.500000 537.650000 1186.000000 538.350000 ;
      RECT 357.500000 537.650000 373.500000 538.350000 ;
      RECT 1157.500000 536.350000 1158.500000 537.650000 ;
      RECT 1139.000000 536.350000 1149.500000 539.650000 ;
      RECT 386.500000 536.350000 389.000000 539.650000 ;
      RECT 372.500000 536.350000 373.500000 537.650000 ;
      RECT 357.500000 536.350000 358.500000 537.650000 ;
      RECT 0.000000 536.350000 349.500000 539.650000 ;
      RECT 1139.000000 535.650000 1158.500000 536.350000 ;
      RECT 372.500000 535.650000 389.000000 536.350000 ;
      RECT 0.000000 535.650000 358.500000 536.350000 ;
      RECT 1166.500000 534.350000 1186.000000 537.650000 ;
      RECT 1157.500000 534.350000 1158.500000 535.650000 ;
      RECT 372.500000 534.350000 373.500000 535.650000 ;
      RECT 357.500000 534.350000 358.500000 535.650000 ;
      RECT 1157.500000 533.650000 1186.000000 534.350000 ;
      RECT 357.500000 533.650000 373.500000 534.350000 ;
      RECT 1157.500000 532.350000 1158.500000 533.650000 ;
      RECT 1139.000000 532.350000 1149.500000 535.650000 ;
      RECT 386.500000 532.350000 389.000000 535.650000 ;
      RECT 372.500000 532.350000 373.500000 533.650000 ;
      RECT 357.500000 532.350000 358.500000 533.650000 ;
      RECT 0.000000 532.350000 349.500000 535.650000 ;
      RECT 1139.000000 531.650000 1158.500000 532.350000 ;
      RECT 372.500000 531.650000 389.000000 532.350000 ;
      RECT 0.000000 531.650000 358.500000 532.350000 ;
      RECT 1166.500000 530.350000 1186.000000 533.650000 ;
      RECT 1157.500000 530.350000 1158.500000 531.650000 ;
      RECT 372.500000 530.350000 373.500000 531.650000 ;
      RECT 357.500000 530.350000 358.500000 531.650000 ;
      RECT 1157.500000 529.650000 1186.000000 530.350000 ;
      RECT 357.500000 529.650000 373.500000 530.350000 ;
      RECT 1157.500000 528.350000 1158.500000 529.650000 ;
      RECT 1139.000000 528.350000 1149.500000 531.650000 ;
      RECT 386.500000 528.350000 389.000000 531.650000 ;
      RECT 372.500000 528.350000 373.500000 529.650000 ;
      RECT 357.500000 528.350000 358.500000 529.650000 ;
      RECT 0.000000 528.350000 349.500000 531.650000 ;
      RECT 1139.000000 527.650000 1158.500000 528.350000 ;
      RECT 372.500000 527.650000 389.000000 528.350000 ;
      RECT 0.000000 527.650000 358.500000 528.350000 ;
      RECT 1166.500000 526.350000 1186.000000 529.650000 ;
      RECT 1157.500000 526.350000 1158.500000 527.650000 ;
      RECT 372.500000 526.350000 373.500000 527.650000 ;
      RECT 357.500000 526.350000 358.500000 527.650000 ;
      RECT 1157.500000 525.650000 1186.000000 526.350000 ;
      RECT 357.500000 525.650000 373.500000 526.350000 ;
      RECT 1157.500000 524.350000 1158.500000 525.650000 ;
      RECT 1139.000000 524.350000 1149.500000 527.650000 ;
      RECT 386.500000 524.350000 389.000000 527.650000 ;
      RECT 372.500000 524.350000 373.500000 525.650000 ;
      RECT 357.500000 524.350000 358.500000 525.650000 ;
      RECT 0.000000 524.350000 349.500000 527.650000 ;
      RECT 1139.000000 523.650000 1158.500000 524.350000 ;
      RECT 372.500000 523.650000 389.000000 524.350000 ;
      RECT 0.000000 523.650000 358.500000 524.350000 ;
      RECT 1166.500000 522.350000 1186.000000 525.650000 ;
      RECT 1157.500000 522.350000 1158.500000 523.650000 ;
      RECT 372.500000 522.350000 373.500000 523.650000 ;
      RECT 357.500000 522.350000 358.500000 523.650000 ;
      RECT 1157.500000 521.650000 1186.000000 522.350000 ;
      RECT 357.500000 521.650000 373.500000 522.350000 ;
      RECT 1157.500000 520.350000 1158.500000 521.650000 ;
      RECT 1139.000000 520.350000 1149.500000 523.650000 ;
      RECT 386.500000 520.350000 389.000000 523.650000 ;
      RECT 372.500000 520.350000 373.500000 521.650000 ;
      RECT 357.500000 520.350000 358.500000 521.650000 ;
      RECT 0.000000 520.350000 349.500000 523.650000 ;
      RECT 1139.000000 519.650000 1158.500000 520.350000 ;
      RECT 372.500000 519.650000 389.000000 520.350000 ;
      RECT 0.000000 519.650000 358.500000 520.350000 ;
      RECT 1166.500000 518.350000 1186.000000 521.650000 ;
      RECT 1157.500000 518.350000 1158.500000 519.650000 ;
      RECT 372.500000 518.350000 373.500000 519.650000 ;
      RECT 357.500000 518.350000 358.500000 519.650000 ;
      RECT 1157.500000 517.650000 1186.000000 518.350000 ;
      RECT 357.500000 517.650000 373.500000 518.350000 ;
      RECT 307.500000 517.650000 349.500000 519.650000 ;
      RECT 0.000000 517.650000 299.500000 519.650000 ;
      RECT 1157.500000 516.350000 1158.500000 517.650000 ;
      RECT 1139.000000 516.350000 1149.500000 519.650000 ;
      RECT 386.500000 516.350000 389.000000 519.650000 ;
      RECT 372.500000 516.350000 373.500000 517.650000 ;
      RECT 357.500000 516.350000 358.500000 517.650000 ;
      RECT 316.500000 516.350000 349.500000 517.650000 ;
      RECT 307.500000 516.350000 308.500000 517.650000 ;
      RECT 266.500000 516.350000 299.500000 517.650000 ;
      RECT 1139.000000 515.650000 1158.500000 516.350000 ;
      RECT 372.500000 515.650000 389.000000 516.350000 ;
      RECT 316.500000 515.650000 358.500000 516.350000 ;
      RECT 266.500000 515.650000 308.500000 516.350000 ;
      RECT 216.500000 515.650000 258.500000 517.650000 ;
      RECT 166.500000 515.650000 208.500000 517.650000 ;
      RECT 116.500000 515.650000 158.500000 517.650000 ;
      RECT 66.500000 515.650000 108.500000 517.650000 ;
      RECT 29.500000 515.650000 58.500000 517.650000 ;
      RECT 0.000000 515.650000 16.500000 517.650000 ;
      RECT 1166.500000 514.350000 1186.000000 517.650000 ;
      RECT 1157.500000 514.350000 1158.500000 515.650000 ;
      RECT 372.500000 514.350000 373.500000 515.650000 ;
      RECT 357.500000 514.350000 358.500000 515.650000 ;
      RECT 316.500000 514.350000 349.500000 515.650000 ;
      RECT 307.500000 514.350000 308.500000 515.650000 ;
      RECT 266.500000 514.350000 299.500000 515.650000 ;
      RECT 257.500000 514.350000 258.500000 515.650000 ;
      RECT 216.500000 514.350000 249.500000 515.650000 ;
      RECT 207.500000 514.350000 208.500000 515.650000 ;
      RECT 166.500000 514.350000 199.500000 515.650000 ;
      RECT 157.500000 514.350000 158.500000 515.650000 ;
      RECT 116.500000 514.350000 149.500000 515.650000 ;
      RECT 107.500000 514.350000 108.500000 515.650000 ;
      RECT 66.500000 514.350000 99.500000 515.650000 ;
      RECT 57.500000 514.350000 58.500000 515.650000 ;
      RECT 29.500000 514.350000 49.500000 515.650000 ;
      RECT 15.500000 514.350000 16.500000 515.650000 ;
      RECT 1157.500000 513.650000 1186.000000 514.350000 ;
      RECT 357.500000 513.650000 373.500000 514.350000 ;
      RECT 307.500000 513.650000 349.500000 514.350000 ;
      RECT 257.500000 513.650000 299.500000 514.350000 ;
      RECT 207.500000 513.650000 249.500000 514.350000 ;
      RECT 157.500000 513.650000 199.500000 514.350000 ;
      RECT 107.500000 513.650000 149.500000 514.350000 ;
      RECT 57.500000 513.650000 99.500000 514.350000 ;
      RECT 15.500000 513.650000 49.500000 514.350000 ;
      RECT 1157.500000 512.350000 1158.500000 513.650000 ;
      RECT 1139.000000 512.350000 1149.500000 515.650000 ;
      RECT 386.500000 512.350000 389.000000 515.650000 ;
      RECT 372.500000 512.350000 373.500000 513.650000 ;
      RECT 357.500000 512.350000 358.500000 513.650000 ;
      RECT 316.500000 512.350000 349.500000 513.650000 ;
      RECT 307.500000 512.350000 308.500000 513.650000 ;
      RECT 266.500000 512.350000 299.500000 513.650000 ;
      RECT 257.500000 512.350000 258.500000 513.650000 ;
      RECT 216.500000 512.350000 249.500000 513.650000 ;
      RECT 207.500000 512.350000 208.500000 513.650000 ;
      RECT 166.500000 512.350000 199.500000 513.650000 ;
      RECT 157.500000 512.350000 158.500000 513.650000 ;
      RECT 116.500000 512.350000 149.500000 513.650000 ;
      RECT 107.500000 512.350000 108.500000 513.650000 ;
      RECT 66.500000 512.350000 99.500000 513.650000 ;
      RECT 57.500000 512.350000 58.500000 513.650000 ;
      RECT 29.500000 512.350000 49.500000 513.650000 ;
      RECT 15.500000 512.350000 16.500000 513.650000 ;
      RECT 0.000000 512.350000 2.500000 515.650000 ;
      RECT 1139.000000 511.650000 1158.500000 512.350000 ;
      RECT 372.500000 511.650000 389.000000 512.350000 ;
      RECT 316.500000 511.650000 358.500000 512.350000 ;
      RECT 266.500000 511.650000 308.500000 512.350000 ;
      RECT 216.500000 511.650000 258.500000 512.350000 ;
      RECT 166.500000 511.650000 208.500000 512.350000 ;
      RECT 116.500000 511.650000 158.500000 512.350000 ;
      RECT 66.500000 511.650000 108.500000 512.350000 ;
      RECT 29.500000 511.650000 58.500000 512.350000 ;
      RECT 0.000000 511.650000 16.500000 512.350000 ;
      RECT 1166.500000 510.350000 1186.000000 513.650000 ;
      RECT 1157.500000 510.350000 1158.500000 511.650000 ;
      RECT 372.500000 510.350000 373.500000 511.650000 ;
      RECT 357.500000 510.350000 358.500000 511.650000 ;
      RECT 316.500000 510.350000 349.500000 511.650000 ;
      RECT 307.500000 510.350000 308.500000 511.650000 ;
      RECT 266.500000 510.350000 299.500000 511.650000 ;
      RECT 257.500000 510.350000 258.500000 511.650000 ;
      RECT 216.500000 510.350000 249.500000 511.650000 ;
      RECT 207.500000 510.350000 208.500000 511.650000 ;
      RECT 166.500000 510.350000 199.500000 511.650000 ;
      RECT 157.500000 510.350000 158.500000 511.650000 ;
      RECT 116.500000 510.350000 149.500000 511.650000 ;
      RECT 107.500000 510.350000 108.500000 511.650000 ;
      RECT 66.500000 510.350000 99.500000 511.650000 ;
      RECT 57.500000 510.350000 58.500000 511.650000 ;
      RECT 29.500000 510.350000 49.500000 511.650000 ;
      RECT 15.500000 510.350000 16.500000 511.650000 ;
      RECT 1157.500000 509.650000 1186.000000 510.350000 ;
      RECT 357.500000 509.650000 373.500000 510.350000 ;
      RECT 307.500000 509.650000 349.500000 510.350000 ;
      RECT 257.500000 509.650000 299.500000 510.350000 ;
      RECT 207.500000 509.650000 249.500000 510.350000 ;
      RECT 157.500000 509.650000 199.500000 510.350000 ;
      RECT 107.500000 509.650000 149.500000 510.350000 ;
      RECT 57.500000 509.650000 99.500000 510.350000 ;
      RECT 15.500000 509.650000 49.500000 510.350000 ;
      RECT 1157.500000 508.350000 1158.500000 509.650000 ;
      RECT 1139.000000 508.350000 1149.500000 511.650000 ;
      RECT 386.500000 508.350000 389.000000 511.650000 ;
      RECT 372.500000 508.350000 373.500000 509.650000 ;
      RECT 357.500000 508.350000 358.500000 509.650000 ;
      RECT 316.500000 508.350000 349.500000 509.650000 ;
      RECT 307.500000 508.350000 308.500000 509.650000 ;
      RECT 266.500000 508.350000 299.500000 509.650000 ;
      RECT 257.500000 508.350000 258.500000 509.650000 ;
      RECT 216.500000 508.350000 249.500000 509.650000 ;
      RECT 207.500000 508.350000 208.500000 509.650000 ;
      RECT 166.500000 508.350000 199.500000 509.650000 ;
      RECT 157.500000 508.350000 158.500000 509.650000 ;
      RECT 116.500000 508.350000 149.500000 509.650000 ;
      RECT 107.500000 508.350000 108.500000 509.650000 ;
      RECT 66.500000 508.350000 99.500000 509.650000 ;
      RECT 57.500000 508.350000 58.500000 509.650000 ;
      RECT 29.500000 508.350000 49.500000 509.650000 ;
      RECT 15.500000 508.350000 16.500000 509.650000 ;
      RECT 0.000000 508.350000 2.500000 511.650000 ;
      RECT 1139.000000 507.650000 1158.500000 508.350000 ;
      RECT 372.500000 507.650000 389.000000 508.350000 ;
      RECT 316.500000 507.650000 358.500000 508.350000 ;
      RECT 266.500000 507.650000 308.500000 508.350000 ;
      RECT 216.500000 507.650000 258.500000 508.350000 ;
      RECT 166.500000 507.650000 208.500000 508.350000 ;
      RECT 116.500000 507.650000 158.500000 508.350000 ;
      RECT 66.500000 507.650000 108.500000 508.350000 ;
      RECT 29.500000 507.650000 58.500000 508.350000 ;
      RECT 0.000000 507.650000 16.500000 508.350000 ;
      RECT 1166.500000 506.350000 1186.000000 509.650000 ;
      RECT 1157.500000 506.350000 1158.500000 507.650000 ;
      RECT 372.500000 506.350000 373.500000 507.650000 ;
      RECT 357.500000 506.350000 358.500000 507.650000 ;
      RECT 316.500000 506.350000 349.500000 507.650000 ;
      RECT 307.500000 506.350000 308.500000 507.650000 ;
      RECT 266.500000 506.350000 299.500000 507.650000 ;
      RECT 257.500000 506.350000 258.500000 507.650000 ;
      RECT 216.500000 506.350000 249.500000 507.650000 ;
      RECT 207.500000 506.350000 208.500000 507.650000 ;
      RECT 166.500000 506.350000 199.500000 507.650000 ;
      RECT 157.500000 506.350000 158.500000 507.650000 ;
      RECT 116.500000 506.350000 149.500000 507.650000 ;
      RECT 107.500000 506.350000 108.500000 507.650000 ;
      RECT 66.500000 506.350000 99.500000 507.650000 ;
      RECT 57.500000 506.350000 58.500000 507.650000 ;
      RECT 29.500000 506.350000 49.500000 507.650000 ;
      RECT 15.500000 506.350000 16.500000 507.650000 ;
      RECT 386.500000 506.000000 389.000000 507.650000 ;
      RECT 1157.500000 505.650000 1186.000000 506.350000 ;
      RECT 386.500000 505.650000 739.000000 506.000000 ;
      RECT 357.500000 505.650000 373.500000 506.350000 ;
      RECT 307.500000 505.650000 349.500000 506.350000 ;
      RECT 257.500000 505.650000 299.500000 506.350000 ;
      RECT 207.500000 505.650000 249.500000 506.350000 ;
      RECT 157.500000 505.650000 199.500000 506.350000 ;
      RECT 107.500000 505.650000 149.500000 506.350000 ;
      RECT 57.500000 505.650000 99.500000 506.350000 ;
      RECT 15.500000 505.650000 49.500000 506.350000 ;
      RECT 1157.500000 504.350000 1158.500000 505.650000 ;
      RECT 1139.000000 504.350000 1149.500000 507.650000 ;
      RECT 386.500000 504.350000 408.500000 505.650000 ;
      RECT 372.500000 504.350000 373.500000 505.650000 ;
      RECT 357.500000 504.350000 358.500000 505.650000 ;
      RECT 316.500000 504.350000 349.500000 505.650000 ;
      RECT 307.500000 504.350000 308.500000 505.650000 ;
      RECT 266.500000 504.350000 299.500000 505.650000 ;
      RECT 257.500000 504.350000 258.500000 505.650000 ;
      RECT 216.500000 504.350000 249.500000 505.650000 ;
      RECT 207.500000 504.350000 208.500000 505.650000 ;
      RECT 166.500000 504.350000 199.500000 505.650000 ;
      RECT 157.500000 504.350000 158.500000 505.650000 ;
      RECT 116.500000 504.350000 149.500000 505.650000 ;
      RECT 107.500000 504.350000 108.500000 505.650000 ;
      RECT 66.500000 504.350000 99.500000 505.650000 ;
      RECT 57.500000 504.350000 58.500000 505.650000 ;
      RECT 29.500000 504.350000 49.500000 505.650000 ;
      RECT 15.500000 504.350000 16.500000 505.650000 ;
      RECT 0.000000 504.350000 2.500000 507.650000 ;
      RECT 1139.000000 503.650000 1158.500000 504.350000 ;
      RECT 716.500000 503.650000 739.000000 505.650000 ;
      RECT 666.500000 503.650000 708.500000 505.650000 ;
      RECT 616.500000 503.650000 658.500000 505.650000 ;
      RECT 566.500000 503.650000 608.500000 505.650000 ;
      RECT 516.500000 503.650000 558.500000 505.650000 ;
      RECT 466.500000 503.650000 508.500000 505.650000 ;
      RECT 416.500000 503.650000 458.500000 505.650000 ;
      RECT 372.500000 503.650000 408.500000 504.350000 ;
      RECT 316.500000 503.650000 358.500000 504.350000 ;
      RECT 266.500000 503.650000 308.500000 504.350000 ;
      RECT 216.500000 503.650000 258.500000 504.350000 ;
      RECT 166.500000 503.650000 208.500000 504.350000 ;
      RECT 116.500000 503.650000 158.500000 504.350000 ;
      RECT 66.500000 503.650000 108.500000 504.350000 ;
      RECT 29.500000 503.650000 58.500000 504.350000 ;
      RECT 0.000000 503.650000 16.500000 504.350000 ;
      RECT 1166.500000 502.350000 1186.000000 505.650000 ;
      RECT 1157.500000 502.350000 1158.500000 503.650000 ;
      RECT 716.500000 502.350000 723.500000 503.650000 ;
      RECT 707.500000 502.350000 708.500000 503.650000 ;
      RECT 666.500000 502.350000 699.500000 503.650000 ;
      RECT 657.500000 502.350000 658.500000 503.650000 ;
      RECT 616.500000 502.350000 649.500000 503.650000 ;
      RECT 607.500000 502.350000 608.500000 503.650000 ;
      RECT 566.500000 502.350000 599.500000 503.650000 ;
      RECT 557.500000 502.350000 558.500000 503.650000 ;
      RECT 516.500000 502.350000 549.500000 503.650000 ;
      RECT 507.500000 502.350000 508.500000 503.650000 ;
      RECT 466.500000 502.350000 499.500000 503.650000 ;
      RECT 457.500000 502.350000 458.500000 503.650000 ;
      RECT 416.500000 502.350000 449.500000 503.650000 ;
      RECT 407.500000 502.350000 408.500000 503.650000 ;
      RECT 372.500000 502.350000 373.500000 503.650000 ;
      RECT 357.500000 502.350000 358.500000 503.650000 ;
      RECT 316.500000 502.350000 349.500000 503.650000 ;
      RECT 307.500000 502.350000 308.500000 503.650000 ;
      RECT 266.500000 502.350000 299.500000 503.650000 ;
      RECT 257.500000 502.350000 258.500000 503.650000 ;
      RECT 216.500000 502.350000 249.500000 503.650000 ;
      RECT 207.500000 502.350000 208.500000 503.650000 ;
      RECT 166.500000 502.350000 199.500000 503.650000 ;
      RECT 157.500000 502.350000 158.500000 503.650000 ;
      RECT 116.500000 502.350000 149.500000 503.650000 ;
      RECT 107.500000 502.350000 108.500000 503.650000 ;
      RECT 66.500000 502.350000 99.500000 503.650000 ;
      RECT 57.500000 502.350000 58.500000 503.650000 ;
      RECT 29.500000 502.350000 49.500000 503.650000 ;
      RECT 15.500000 502.350000 16.500000 503.650000 ;
      RECT 1157.500000 501.650000 1186.000000 502.350000 ;
      RECT 707.500000 501.650000 723.500000 502.350000 ;
      RECT 657.500000 501.650000 699.500000 502.350000 ;
      RECT 607.500000 501.650000 649.500000 502.350000 ;
      RECT 557.500000 501.650000 599.500000 502.350000 ;
      RECT 507.500000 501.650000 549.500000 502.350000 ;
      RECT 457.500000 501.650000 499.500000 502.350000 ;
      RECT 407.500000 501.650000 449.500000 502.350000 ;
      RECT 357.500000 501.650000 373.500000 502.350000 ;
      RECT 307.500000 501.650000 349.500000 502.350000 ;
      RECT 257.500000 501.650000 299.500000 502.350000 ;
      RECT 207.500000 501.650000 249.500000 502.350000 ;
      RECT 157.500000 501.650000 199.500000 502.350000 ;
      RECT 107.500000 501.650000 149.500000 502.350000 ;
      RECT 57.500000 501.650000 99.500000 502.350000 ;
      RECT 15.500000 501.650000 49.500000 502.350000 ;
      RECT 1157.500000 500.350000 1158.500000 501.650000 ;
      RECT 1139.000000 500.350000 1149.500000 503.650000 ;
      RECT 736.500000 500.350000 739.000000 503.650000 ;
      RECT 716.500000 500.350000 723.500000 501.650000 ;
      RECT 707.500000 500.350000 708.500000 501.650000 ;
      RECT 666.500000 500.350000 699.500000 501.650000 ;
      RECT 657.500000 500.350000 658.500000 501.650000 ;
      RECT 616.500000 500.350000 649.500000 501.650000 ;
      RECT 607.500000 500.350000 608.500000 501.650000 ;
      RECT 566.500000 500.350000 599.500000 501.650000 ;
      RECT 557.500000 500.350000 558.500000 501.650000 ;
      RECT 516.500000 500.350000 549.500000 501.650000 ;
      RECT 507.500000 500.350000 508.500000 501.650000 ;
      RECT 466.500000 500.350000 499.500000 501.650000 ;
      RECT 457.500000 500.350000 458.500000 501.650000 ;
      RECT 416.500000 500.350000 449.500000 501.650000 ;
      RECT 407.500000 500.350000 408.500000 501.650000 ;
      RECT 386.500000 500.350000 399.500000 503.650000 ;
      RECT 372.500000 500.350000 373.500000 501.650000 ;
      RECT 357.500000 500.350000 358.500000 501.650000 ;
      RECT 316.500000 500.350000 349.500000 501.650000 ;
      RECT 307.500000 500.350000 308.500000 501.650000 ;
      RECT 266.500000 500.350000 299.500000 501.650000 ;
      RECT 257.500000 500.350000 258.500000 501.650000 ;
      RECT 216.500000 500.350000 249.500000 501.650000 ;
      RECT 207.500000 500.350000 208.500000 501.650000 ;
      RECT 166.500000 500.350000 199.500000 501.650000 ;
      RECT 157.500000 500.350000 158.500000 501.650000 ;
      RECT 116.500000 500.350000 149.500000 501.650000 ;
      RECT 107.500000 500.350000 108.500000 501.650000 ;
      RECT 66.500000 500.350000 99.500000 501.650000 ;
      RECT 57.500000 500.350000 58.500000 501.650000 ;
      RECT 29.500000 500.350000 49.500000 501.650000 ;
      RECT 15.500000 500.350000 16.500000 501.650000 ;
      RECT 0.000000 500.350000 2.500000 503.650000 ;
      RECT 1139.000000 499.650000 1158.500000 500.350000 ;
      RECT 716.500000 499.650000 739.000000 500.350000 ;
      RECT 666.500000 499.650000 708.500000 500.350000 ;
      RECT 616.500000 499.650000 658.500000 500.350000 ;
      RECT 566.500000 499.650000 608.500000 500.350000 ;
      RECT 516.500000 499.650000 558.500000 500.350000 ;
      RECT 466.500000 499.650000 508.500000 500.350000 ;
      RECT 416.500000 499.650000 458.500000 500.350000 ;
      RECT 372.500000 499.650000 408.500000 500.350000 ;
      RECT 316.500000 499.650000 358.500000 500.350000 ;
      RECT 266.500000 499.650000 308.500000 500.350000 ;
      RECT 216.500000 499.650000 258.500000 500.350000 ;
      RECT 166.500000 499.650000 208.500000 500.350000 ;
      RECT 116.500000 499.650000 158.500000 500.350000 ;
      RECT 66.500000 499.650000 108.500000 500.350000 ;
      RECT 29.500000 499.650000 58.500000 500.350000 ;
      RECT 0.000000 499.650000 16.500000 500.350000 ;
      RECT 1166.500000 498.350000 1186.000000 501.650000 ;
      RECT 1157.500000 498.350000 1158.500000 499.650000 ;
      RECT 716.500000 498.350000 723.500000 499.650000 ;
      RECT 707.500000 498.350000 708.500000 499.650000 ;
      RECT 666.500000 498.350000 699.500000 499.650000 ;
      RECT 657.500000 498.350000 658.500000 499.650000 ;
      RECT 616.500000 498.350000 649.500000 499.650000 ;
      RECT 607.500000 498.350000 608.500000 499.650000 ;
      RECT 566.500000 498.350000 599.500000 499.650000 ;
      RECT 557.500000 498.350000 558.500000 499.650000 ;
      RECT 516.500000 498.350000 549.500000 499.650000 ;
      RECT 507.500000 498.350000 508.500000 499.650000 ;
      RECT 466.500000 498.350000 499.500000 499.650000 ;
      RECT 457.500000 498.350000 458.500000 499.650000 ;
      RECT 416.500000 498.350000 449.500000 499.650000 ;
      RECT 407.500000 498.350000 408.500000 499.650000 ;
      RECT 372.500000 498.350000 373.500000 499.650000 ;
      RECT 357.500000 498.350000 358.500000 499.650000 ;
      RECT 316.500000 498.350000 349.500000 499.650000 ;
      RECT 307.500000 498.350000 308.500000 499.650000 ;
      RECT 266.500000 498.350000 299.500000 499.650000 ;
      RECT 257.500000 498.350000 258.500000 499.650000 ;
      RECT 216.500000 498.350000 249.500000 499.650000 ;
      RECT 207.500000 498.350000 208.500000 499.650000 ;
      RECT 166.500000 498.350000 199.500000 499.650000 ;
      RECT 157.500000 498.350000 158.500000 499.650000 ;
      RECT 116.500000 498.350000 149.500000 499.650000 ;
      RECT 107.500000 498.350000 108.500000 499.650000 ;
      RECT 66.500000 498.350000 99.500000 499.650000 ;
      RECT 57.500000 498.350000 58.500000 499.650000 ;
      RECT 29.500000 498.350000 49.500000 499.650000 ;
      RECT 15.500000 498.350000 16.500000 499.650000 ;
      RECT 1157.500000 497.650000 1186.000000 498.350000 ;
      RECT 707.500000 497.650000 723.500000 498.350000 ;
      RECT 657.500000 497.650000 699.500000 498.350000 ;
      RECT 607.500000 497.650000 649.500000 498.350000 ;
      RECT 557.500000 497.650000 599.500000 498.350000 ;
      RECT 507.500000 497.650000 549.500000 498.350000 ;
      RECT 457.500000 497.650000 499.500000 498.350000 ;
      RECT 407.500000 497.650000 449.500000 498.350000 ;
      RECT 357.500000 497.650000 373.500000 498.350000 ;
      RECT 307.500000 497.650000 349.500000 498.350000 ;
      RECT 257.500000 497.650000 299.500000 498.350000 ;
      RECT 207.500000 497.650000 249.500000 498.350000 ;
      RECT 157.500000 497.650000 199.500000 498.350000 ;
      RECT 107.500000 497.650000 149.500000 498.350000 ;
      RECT 57.500000 497.650000 99.500000 498.350000 ;
      RECT 15.500000 497.650000 49.500000 498.350000 ;
      RECT 1157.500000 496.350000 1158.500000 497.650000 ;
      RECT 1139.000000 496.350000 1149.500000 499.650000 ;
      RECT 736.500000 496.350000 739.000000 499.650000 ;
      RECT 716.500000 496.350000 723.500000 497.650000 ;
      RECT 707.500000 496.350000 708.500000 497.650000 ;
      RECT 666.500000 496.350000 699.500000 497.650000 ;
      RECT 657.500000 496.350000 658.500000 497.650000 ;
      RECT 616.500000 496.350000 649.500000 497.650000 ;
      RECT 607.500000 496.350000 608.500000 497.650000 ;
      RECT 566.500000 496.350000 599.500000 497.650000 ;
      RECT 557.500000 496.350000 558.500000 497.650000 ;
      RECT 516.500000 496.350000 549.500000 497.650000 ;
      RECT 507.500000 496.350000 508.500000 497.650000 ;
      RECT 466.500000 496.350000 499.500000 497.650000 ;
      RECT 457.500000 496.350000 458.500000 497.650000 ;
      RECT 416.500000 496.350000 449.500000 497.650000 ;
      RECT 407.500000 496.350000 408.500000 497.650000 ;
      RECT 386.500000 496.350000 399.500000 499.650000 ;
      RECT 372.500000 496.350000 373.500000 497.650000 ;
      RECT 357.500000 496.350000 358.500000 497.650000 ;
      RECT 316.500000 496.350000 349.500000 497.650000 ;
      RECT 307.500000 496.350000 308.500000 497.650000 ;
      RECT 266.500000 496.350000 299.500000 497.650000 ;
      RECT 257.500000 496.350000 258.500000 497.650000 ;
      RECT 216.500000 496.350000 249.500000 497.650000 ;
      RECT 207.500000 496.350000 208.500000 497.650000 ;
      RECT 166.500000 496.350000 199.500000 497.650000 ;
      RECT 157.500000 496.350000 158.500000 497.650000 ;
      RECT 116.500000 496.350000 149.500000 497.650000 ;
      RECT 107.500000 496.350000 108.500000 497.650000 ;
      RECT 66.500000 496.350000 99.500000 497.650000 ;
      RECT 57.500000 496.350000 58.500000 497.650000 ;
      RECT 29.500000 496.350000 49.500000 497.650000 ;
      RECT 15.500000 496.350000 16.500000 497.650000 ;
      RECT 0.000000 496.350000 2.500000 499.650000 ;
      RECT 1139.000000 495.650000 1158.500000 496.350000 ;
      RECT 716.500000 495.650000 739.000000 496.350000 ;
      RECT 666.500000 495.650000 708.500000 496.350000 ;
      RECT 616.500000 495.650000 658.500000 496.350000 ;
      RECT 566.500000 495.650000 608.500000 496.350000 ;
      RECT 516.500000 495.650000 558.500000 496.350000 ;
      RECT 466.500000 495.650000 508.500000 496.350000 ;
      RECT 416.500000 495.650000 458.500000 496.350000 ;
      RECT 372.500000 495.650000 408.500000 496.350000 ;
      RECT 316.500000 495.650000 358.500000 496.350000 ;
      RECT 266.500000 495.650000 308.500000 496.350000 ;
      RECT 216.500000 495.650000 258.500000 496.350000 ;
      RECT 166.500000 495.650000 208.500000 496.350000 ;
      RECT 116.500000 495.650000 158.500000 496.350000 ;
      RECT 66.500000 495.650000 108.500000 496.350000 ;
      RECT 29.500000 495.650000 58.500000 496.350000 ;
      RECT 0.000000 495.650000 16.500000 496.350000 ;
      RECT 1166.500000 494.350000 1186.000000 497.650000 ;
      RECT 1157.500000 494.350000 1158.500000 495.650000 ;
      RECT 716.500000 494.350000 723.500000 495.650000 ;
      RECT 707.500000 494.350000 708.500000 495.650000 ;
      RECT 666.500000 494.350000 699.500000 495.650000 ;
      RECT 657.500000 494.350000 658.500000 495.650000 ;
      RECT 616.500000 494.350000 649.500000 495.650000 ;
      RECT 607.500000 494.350000 608.500000 495.650000 ;
      RECT 566.500000 494.350000 599.500000 495.650000 ;
      RECT 557.500000 494.350000 558.500000 495.650000 ;
      RECT 516.500000 494.350000 549.500000 495.650000 ;
      RECT 507.500000 494.350000 508.500000 495.650000 ;
      RECT 466.500000 494.350000 499.500000 495.650000 ;
      RECT 457.500000 494.350000 458.500000 495.650000 ;
      RECT 416.500000 494.350000 449.500000 495.650000 ;
      RECT 407.500000 494.350000 408.500000 495.650000 ;
      RECT 372.500000 494.350000 373.500000 495.650000 ;
      RECT 357.500000 494.350000 358.500000 495.650000 ;
      RECT 316.500000 494.350000 349.500000 495.650000 ;
      RECT 307.500000 494.350000 308.500000 495.650000 ;
      RECT 266.500000 494.350000 299.500000 495.650000 ;
      RECT 257.500000 494.350000 258.500000 495.650000 ;
      RECT 216.500000 494.350000 249.500000 495.650000 ;
      RECT 207.500000 494.350000 208.500000 495.650000 ;
      RECT 166.500000 494.350000 199.500000 495.650000 ;
      RECT 157.500000 494.350000 158.500000 495.650000 ;
      RECT 116.500000 494.350000 149.500000 495.650000 ;
      RECT 107.500000 494.350000 108.500000 495.650000 ;
      RECT 66.500000 494.350000 99.500000 495.650000 ;
      RECT 57.500000 494.350000 58.500000 495.650000 ;
      RECT 29.500000 494.350000 49.500000 495.650000 ;
      RECT 15.500000 494.350000 16.500000 495.650000 ;
      RECT 1157.500000 493.650000 1186.000000 494.350000 ;
      RECT 707.500000 493.650000 723.500000 494.350000 ;
      RECT 657.500000 493.650000 699.500000 494.350000 ;
      RECT 607.500000 493.650000 649.500000 494.350000 ;
      RECT 557.500000 493.650000 599.500000 494.350000 ;
      RECT 507.500000 493.650000 549.500000 494.350000 ;
      RECT 457.500000 493.650000 499.500000 494.350000 ;
      RECT 407.500000 493.650000 449.500000 494.350000 ;
      RECT 357.500000 493.650000 373.500000 494.350000 ;
      RECT 307.500000 493.650000 349.500000 494.350000 ;
      RECT 257.500000 493.650000 299.500000 494.350000 ;
      RECT 207.500000 493.650000 249.500000 494.350000 ;
      RECT 157.500000 493.650000 199.500000 494.350000 ;
      RECT 107.500000 493.650000 149.500000 494.350000 ;
      RECT 57.500000 493.650000 99.500000 494.350000 ;
      RECT 15.500000 493.650000 49.500000 494.350000 ;
      RECT 1157.500000 492.350000 1158.500000 493.650000 ;
      RECT 1139.000000 492.350000 1149.500000 495.650000 ;
      RECT 736.500000 492.350000 739.000000 495.650000 ;
      RECT 716.500000 492.350000 723.500000 493.650000 ;
      RECT 707.500000 492.350000 708.500000 493.650000 ;
      RECT 666.500000 492.350000 699.500000 493.650000 ;
      RECT 657.500000 492.350000 658.500000 493.650000 ;
      RECT 616.500000 492.350000 649.500000 493.650000 ;
      RECT 607.500000 492.350000 608.500000 493.650000 ;
      RECT 566.500000 492.350000 599.500000 493.650000 ;
      RECT 557.500000 492.350000 558.500000 493.650000 ;
      RECT 516.500000 492.350000 549.500000 493.650000 ;
      RECT 507.500000 492.350000 508.500000 493.650000 ;
      RECT 466.500000 492.350000 499.500000 493.650000 ;
      RECT 457.500000 492.350000 458.500000 493.650000 ;
      RECT 416.500000 492.350000 449.500000 493.650000 ;
      RECT 407.500000 492.350000 408.500000 493.650000 ;
      RECT 386.500000 492.350000 399.500000 495.650000 ;
      RECT 372.500000 492.350000 373.500000 493.650000 ;
      RECT 357.500000 492.350000 358.500000 493.650000 ;
      RECT 316.500000 492.350000 349.500000 493.650000 ;
      RECT 307.500000 492.350000 308.500000 493.650000 ;
      RECT 266.500000 492.350000 299.500000 493.650000 ;
      RECT 257.500000 492.350000 258.500000 493.650000 ;
      RECT 216.500000 492.350000 249.500000 493.650000 ;
      RECT 207.500000 492.350000 208.500000 493.650000 ;
      RECT 166.500000 492.350000 199.500000 493.650000 ;
      RECT 157.500000 492.350000 158.500000 493.650000 ;
      RECT 116.500000 492.350000 149.500000 493.650000 ;
      RECT 107.500000 492.350000 108.500000 493.650000 ;
      RECT 66.500000 492.350000 99.500000 493.650000 ;
      RECT 57.500000 492.350000 58.500000 493.650000 ;
      RECT 29.500000 492.350000 49.500000 493.650000 ;
      RECT 15.500000 492.350000 16.500000 493.650000 ;
      RECT 0.000000 492.350000 2.500000 495.650000 ;
      RECT 1139.000000 491.650000 1158.500000 492.350000 ;
      RECT 716.500000 491.650000 739.000000 492.350000 ;
      RECT 666.500000 491.650000 708.500000 492.350000 ;
      RECT 616.500000 491.650000 658.500000 492.350000 ;
      RECT 566.500000 491.650000 608.500000 492.350000 ;
      RECT 516.500000 491.650000 558.500000 492.350000 ;
      RECT 466.500000 491.650000 508.500000 492.350000 ;
      RECT 416.500000 491.650000 458.500000 492.350000 ;
      RECT 372.500000 491.650000 408.500000 492.350000 ;
      RECT 316.500000 491.650000 358.500000 492.350000 ;
      RECT 266.500000 491.650000 308.500000 492.350000 ;
      RECT 216.500000 491.650000 258.500000 492.350000 ;
      RECT 166.500000 491.650000 208.500000 492.350000 ;
      RECT 116.500000 491.650000 158.500000 492.350000 ;
      RECT 66.500000 491.650000 108.500000 492.350000 ;
      RECT 29.500000 491.650000 58.500000 492.350000 ;
      RECT 0.000000 491.650000 16.500000 492.350000 ;
      RECT 1166.500000 490.350000 1186.000000 493.650000 ;
      RECT 1157.500000 490.350000 1158.500000 491.650000 ;
      RECT 716.500000 490.350000 723.500000 491.650000 ;
      RECT 707.500000 490.350000 708.500000 491.650000 ;
      RECT 666.500000 490.350000 699.500000 491.650000 ;
      RECT 657.500000 490.350000 658.500000 491.650000 ;
      RECT 616.500000 490.350000 649.500000 491.650000 ;
      RECT 607.500000 490.350000 608.500000 491.650000 ;
      RECT 566.500000 490.350000 599.500000 491.650000 ;
      RECT 557.500000 490.350000 558.500000 491.650000 ;
      RECT 516.500000 490.350000 549.500000 491.650000 ;
      RECT 507.500000 490.350000 508.500000 491.650000 ;
      RECT 466.500000 490.350000 499.500000 491.650000 ;
      RECT 457.500000 490.350000 458.500000 491.650000 ;
      RECT 416.500000 490.350000 449.500000 491.650000 ;
      RECT 407.500000 490.350000 408.500000 491.650000 ;
      RECT 372.500000 490.350000 399.500000 491.650000 ;
      RECT 357.500000 490.350000 358.500000 491.650000 ;
      RECT 316.500000 490.350000 349.500000 491.650000 ;
      RECT 307.500000 490.350000 308.500000 491.650000 ;
      RECT 266.500000 490.350000 299.500000 491.650000 ;
      RECT 257.500000 490.350000 258.500000 491.650000 ;
      RECT 216.500000 490.350000 249.500000 491.650000 ;
      RECT 207.500000 490.350000 208.500000 491.650000 ;
      RECT 166.500000 490.350000 199.500000 491.650000 ;
      RECT 157.500000 490.350000 158.500000 491.650000 ;
      RECT 116.500000 490.350000 149.500000 491.650000 ;
      RECT 107.500000 490.350000 108.500000 491.650000 ;
      RECT 66.500000 490.350000 99.500000 491.650000 ;
      RECT 57.500000 490.350000 58.500000 491.650000 ;
      RECT 29.500000 490.350000 49.500000 491.650000 ;
      RECT 15.500000 490.350000 16.500000 491.650000 ;
      RECT 1157.500000 489.650000 1186.000000 490.350000 ;
      RECT 707.500000 489.650000 723.500000 490.350000 ;
      RECT 657.500000 489.650000 699.500000 490.350000 ;
      RECT 607.500000 489.650000 649.500000 490.350000 ;
      RECT 557.500000 489.650000 599.500000 490.350000 ;
      RECT 507.500000 489.650000 549.500000 490.350000 ;
      RECT 457.500000 489.650000 499.500000 490.350000 ;
      RECT 407.500000 489.650000 449.500000 490.350000 ;
      RECT 357.500000 489.650000 399.500000 490.350000 ;
      RECT 307.500000 489.650000 349.500000 490.350000 ;
      RECT 257.500000 489.650000 299.500000 490.350000 ;
      RECT 207.500000 489.650000 249.500000 490.350000 ;
      RECT 157.500000 489.650000 199.500000 490.350000 ;
      RECT 107.500000 489.650000 149.500000 490.350000 ;
      RECT 57.500000 489.650000 99.500000 490.350000 ;
      RECT 15.500000 489.650000 49.500000 490.350000 ;
      RECT 1157.500000 488.350000 1158.500000 489.650000 ;
      RECT 1139.000000 488.350000 1149.500000 491.650000 ;
      RECT 736.500000 488.350000 739.000000 491.650000 ;
      RECT 722.500000 488.350000 723.500000 489.650000 ;
      RECT 707.500000 488.350000 708.500000 489.650000 ;
      RECT 666.500000 488.350000 699.500000 489.650000 ;
      RECT 657.500000 488.350000 658.500000 489.650000 ;
      RECT 616.500000 488.350000 649.500000 489.650000 ;
      RECT 607.500000 488.350000 608.500000 489.650000 ;
      RECT 566.500000 488.350000 599.500000 489.650000 ;
      RECT 557.500000 488.350000 558.500000 489.650000 ;
      RECT 516.500000 488.350000 549.500000 489.650000 ;
      RECT 507.500000 488.350000 508.500000 489.650000 ;
      RECT 466.500000 488.350000 499.500000 489.650000 ;
      RECT 457.500000 488.350000 458.500000 489.650000 ;
      RECT 416.500000 488.350000 449.500000 489.650000 ;
      RECT 407.500000 488.350000 408.500000 489.650000 ;
      RECT 372.500000 488.350000 399.500000 489.650000 ;
      RECT 357.500000 488.350000 359.500000 489.650000 ;
      RECT 316.500000 488.350000 349.500000 489.650000 ;
      RECT 307.500000 488.350000 308.500000 489.650000 ;
      RECT 266.500000 488.350000 299.500000 489.650000 ;
      RECT 257.500000 488.350000 258.500000 489.650000 ;
      RECT 216.500000 488.350000 249.500000 489.650000 ;
      RECT 207.500000 488.350000 208.500000 489.650000 ;
      RECT 166.500000 488.350000 199.500000 489.650000 ;
      RECT 157.500000 488.350000 158.500000 489.650000 ;
      RECT 116.500000 488.350000 149.500000 489.650000 ;
      RECT 107.500000 488.350000 108.500000 489.650000 ;
      RECT 66.500000 488.350000 99.500000 489.650000 ;
      RECT 57.500000 488.350000 58.500000 489.650000 ;
      RECT 29.500000 488.350000 49.500000 489.650000 ;
      RECT 15.500000 488.350000 16.500000 489.650000 ;
      RECT 0.000000 488.350000 2.500000 491.650000 ;
      RECT 1139.000000 487.650000 1158.500000 488.350000 ;
      RECT 722.500000 487.650000 739.000000 488.350000 ;
      RECT 666.500000 487.650000 708.500000 488.350000 ;
      RECT 616.500000 487.650000 658.500000 488.350000 ;
      RECT 566.500000 487.650000 608.500000 488.350000 ;
      RECT 516.500000 487.650000 558.500000 488.350000 ;
      RECT 466.500000 487.650000 508.500000 488.350000 ;
      RECT 416.500000 487.650000 458.500000 488.350000 ;
      RECT 372.500000 487.650000 408.500000 488.350000 ;
      RECT 316.500000 487.650000 359.500000 488.350000 ;
      RECT 266.500000 487.650000 308.500000 488.350000 ;
      RECT 216.500000 487.650000 258.500000 488.350000 ;
      RECT 166.500000 487.650000 208.500000 488.350000 ;
      RECT 116.500000 487.650000 158.500000 488.350000 ;
      RECT 66.500000 487.650000 108.500000 488.350000 ;
      RECT 29.500000 487.650000 58.500000 488.350000 ;
      RECT 0.000000 487.650000 16.500000 488.350000 ;
      RECT 1166.500000 486.350000 1186.000000 489.650000 ;
      RECT 1157.500000 486.350000 1158.500000 487.650000 ;
      RECT 722.500000 486.350000 723.500000 487.650000 ;
      RECT 707.500000 486.350000 708.500000 487.650000 ;
      RECT 666.500000 486.350000 699.500000 487.650000 ;
      RECT 657.500000 486.350000 658.500000 487.650000 ;
      RECT 616.500000 486.350000 649.500000 487.650000 ;
      RECT 607.500000 486.350000 608.500000 487.650000 ;
      RECT 566.500000 486.350000 599.500000 487.650000 ;
      RECT 557.500000 486.350000 558.500000 487.650000 ;
      RECT 516.500000 486.350000 549.500000 487.650000 ;
      RECT 507.500000 486.350000 508.500000 487.650000 ;
      RECT 466.500000 486.350000 499.500000 487.650000 ;
      RECT 457.500000 486.350000 458.500000 487.650000 ;
      RECT 416.500000 486.350000 449.500000 487.650000 ;
      RECT 407.500000 486.350000 408.500000 487.650000 ;
      RECT 372.500000 486.350000 399.500000 487.650000 ;
      RECT 357.500000 486.350000 359.500000 487.650000 ;
      RECT 316.500000 486.350000 349.500000 487.650000 ;
      RECT 307.500000 486.350000 308.500000 487.650000 ;
      RECT 266.500000 486.350000 299.500000 487.650000 ;
      RECT 257.500000 486.350000 258.500000 487.650000 ;
      RECT 216.500000 486.350000 249.500000 487.650000 ;
      RECT 207.500000 486.350000 208.500000 487.650000 ;
      RECT 166.500000 486.350000 199.500000 487.650000 ;
      RECT 157.500000 486.350000 158.500000 487.650000 ;
      RECT 116.500000 486.350000 149.500000 487.650000 ;
      RECT 107.500000 486.350000 108.500000 487.650000 ;
      RECT 66.500000 486.350000 99.500000 487.650000 ;
      RECT 57.500000 486.350000 58.500000 487.650000 ;
      RECT 29.500000 486.350000 49.500000 487.650000 ;
      RECT 15.500000 486.350000 16.500000 487.650000 ;
      RECT 1157.500000 485.650000 1186.000000 486.350000 ;
      RECT 707.500000 485.650000 723.500000 486.350000 ;
      RECT 657.500000 485.650000 699.500000 486.350000 ;
      RECT 607.500000 485.650000 649.500000 486.350000 ;
      RECT 557.500000 485.650000 599.500000 486.350000 ;
      RECT 507.500000 485.650000 549.500000 486.350000 ;
      RECT 457.500000 485.650000 499.500000 486.350000 ;
      RECT 407.500000 485.650000 449.500000 486.350000 ;
      RECT 357.500000 485.650000 399.500000 486.350000 ;
      RECT 307.500000 485.650000 349.500000 486.350000 ;
      RECT 257.500000 485.650000 299.500000 486.350000 ;
      RECT 207.500000 485.650000 249.500000 486.350000 ;
      RECT 157.500000 485.650000 199.500000 486.350000 ;
      RECT 107.500000 485.650000 149.500000 486.350000 ;
      RECT 57.500000 485.650000 99.500000 486.350000 ;
      RECT 15.500000 485.650000 49.500000 486.350000 ;
      RECT 1157.500000 484.350000 1158.500000 485.650000 ;
      RECT 1139.000000 484.350000 1149.500000 487.650000 ;
      RECT 736.500000 484.350000 739.000000 487.650000 ;
      RECT 722.500000 484.350000 723.500000 485.650000 ;
      RECT 707.500000 484.350000 708.500000 485.650000 ;
      RECT 666.500000 484.350000 699.500000 485.650000 ;
      RECT 657.500000 484.350000 658.500000 485.650000 ;
      RECT 616.500000 484.350000 649.500000 485.650000 ;
      RECT 607.500000 484.350000 608.500000 485.650000 ;
      RECT 566.500000 484.350000 599.500000 485.650000 ;
      RECT 557.500000 484.350000 558.500000 485.650000 ;
      RECT 516.500000 484.350000 549.500000 485.650000 ;
      RECT 507.500000 484.350000 508.500000 485.650000 ;
      RECT 466.500000 484.350000 499.500000 485.650000 ;
      RECT 457.500000 484.350000 458.500000 485.650000 ;
      RECT 416.500000 484.350000 449.500000 485.650000 ;
      RECT 407.500000 484.350000 408.500000 485.650000 ;
      RECT 372.500000 484.350000 399.500000 485.650000 ;
      RECT 357.500000 484.350000 359.500000 485.650000 ;
      RECT 316.500000 484.350000 349.500000 485.650000 ;
      RECT 307.500000 484.350000 308.500000 485.650000 ;
      RECT 266.500000 484.350000 299.500000 485.650000 ;
      RECT 257.500000 484.350000 258.500000 485.650000 ;
      RECT 216.500000 484.350000 249.500000 485.650000 ;
      RECT 207.500000 484.350000 208.500000 485.650000 ;
      RECT 166.500000 484.350000 199.500000 485.650000 ;
      RECT 157.500000 484.350000 158.500000 485.650000 ;
      RECT 116.500000 484.350000 149.500000 485.650000 ;
      RECT 107.500000 484.350000 108.500000 485.650000 ;
      RECT 66.500000 484.350000 99.500000 485.650000 ;
      RECT 57.500000 484.350000 58.500000 485.650000 ;
      RECT 29.500000 484.350000 49.500000 485.650000 ;
      RECT 15.500000 484.350000 16.500000 485.650000 ;
      RECT 0.000000 484.350000 2.500000 487.650000 ;
      RECT 1139.000000 483.650000 1158.500000 484.350000 ;
      RECT 722.500000 483.650000 739.000000 484.350000 ;
      RECT 666.500000 483.650000 708.500000 484.350000 ;
      RECT 616.500000 483.650000 658.500000 484.350000 ;
      RECT 566.500000 483.650000 608.500000 484.350000 ;
      RECT 516.500000 483.650000 558.500000 484.350000 ;
      RECT 466.500000 483.650000 508.500000 484.350000 ;
      RECT 416.500000 483.650000 458.500000 484.350000 ;
      RECT 372.500000 483.650000 408.500000 484.350000 ;
      RECT 316.500000 483.650000 359.500000 484.350000 ;
      RECT 266.500000 483.650000 308.500000 484.350000 ;
      RECT 216.500000 483.650000 258.500000 484.350000 ;
      RECT 166.500000 483.650000 208.500000 484.350000 ;
      RECT 116.500000 483.650000 158.500000 484.350000 ;
      RECT 66.500000 483.650000 108.500000 484.350000 ;
      RECT 29.500000 483.650000 58.500000 484.350000 ;
      RECT 0.000000 483.650000 16.500000 484.350000 ;
      RECT 1166.500000 482.350000 1186.000000 485.650000 ;
      RECT 1157.500000 482.350000 1158.500000 483.650000 ;
      RECT 722.500000 482.350000 723.500000 483.650000 ;
      RECT 707.500000 482.350000 708.500000 483.650000 ;
      RECT 666.500000 482.350000 699.500000 483.650000 ;
      RECT 657.500000 482.350000 658.500000 483.650000 ;
      RECT 616.500000 482.350000 649.500000 483.650000 ;
      RECT 607.500000 482.350000 608.500000 483.650000 ;
      RECT 566.500000 482.350000 599.500000 483.650000 ;
      RECT 557.500000 482.350000 558.500000 483.650000 ;
      RECT 516.500000 482.350000 549.500000 483.650000 ;
      RECT 507.500000 482.350000 508.500000 483.650000 ;
      RECT 466.500000 482.350000 499.500000 483.650000 ;
      RECT 457.500000 482.350000 458.500000 483.650000 ;
      RECT 416.500000 482.350000 449.500000 483.650000 ;
      RECT 407.500000 482.350000 408.500000 483.650000 ;
      RECT 372.500000 482.350000 399.500000 483.650000 ;
      RECT 357.500000 482.350000 359.500000 483.650000 ;
      RECT 316.500000 482.350000 349.500000 483.650000 ;
      RECT 307.500000 482.350000 308.500000 483.650000 ;
      RECT 266.500000 482.350000 299.500000 483.650000 ;
      RECT 257.500000 482.350000 258.500000 483.650000 ;
      RECT 216.500000 482.350000 249.500000 483.650000 ;
      RECT 207.500000 482.350000 208.500000 483.650000 ;
      RECT 166.500000 482.350000 199.500000 483.650000 ;
      RECT 157.500000 482.350000 158.500000 483.650000 ;
      RECT 116.500000 482.350000 149.500000 483.650000 ;
      RECT 107.500000 482.350000 108.500000 483.650000 ;
      RECT 66.500000 482.350000 99.500000 483.650000 ;
      RECT 57.500000 482.350000 58.500000 483.650000 ;
      RECT 29.500000 482.350000 49.500000 483.650000 ;
      RECT 15.500000 482.350000 16.500000 483.650000 ;
      RECT 1157.500000 481.650000 1186.000000 482.350000 ;
      RECT 707.500000 481.650000 723.500000 482.350000 ;
      RECT 657.500000 481.650000 699.500000 482.350000 ;
      RECT 607.500000 481.650000 649.500000 482.350000 ;
      RECT 557.500000 481.650000 599.500000 482.350000 ;
      RECT 507.500000 481.650000 549.500000 482.350000 ;
      RECT 457.500000 481.650000 499.500000 482.350000 ;
      RECT 407.500000 481.650000 449.500000 482.350000 ;
      RECT 357.500000 481.650000 399.500000 482.350000 ;
      RECT 307.500000 481.650000 349.500000 482.350000 ;
      RECT 257.500000 481.650000 299.500000 482.350000 ;
      RECT 207.500000 481.650000 249.500000 482.350000 ;
      RECT 157.500000 481.650000 199.500000 482.350000 ;
      RECT 107.500000 481.650000 149.500000 482.350000 ;
      RECT 57.500000 481.650000 99.500000 482.350000 ;
      RECT 15.500000 481.650000 49.500000 482.350000 ;
      RECT 1157.500000 480.350000 1158.500000 481.650000 ;
      RECT 1139.000000 480.350000 1149.500000 483.650000 ;
      RECT 736.500000 480.350000 739.000000 483.650000 ;
      RECT 722.500000 480.350000 723.500000 481.650000 ;
      RECT 707.500000 480.350000 708.500000 481.650000 ;
      RECT 666.500000 480.350000 699.500000 481.650000 ;
      RECT 657.500000 480.350000 658.500000 481.650000 ;
      RECT 616.500000 480.350000 649.500000 481.650000 ;
      RECT 607.500000 480.350000 608.500000 481.650000 ;
      RECT 566.500000 480.350000 599.500000 481.650000 ;
      RECT 557.500000 480.350000 558.500000 481.650000 ;
      RECT 516.500000 480.350000 549.500000 481.650000 ;
      RECT 507.500000 480.350000 508.500000 481.650000 ;
      RECT 466.500000 480.350000 499.500000 481.650000 ;
      RECT 457.500000 480.350000 458.500000 481.650000 ;
      RECT 416.500000 480.350000 449.500000 481.650000 ;
      RECT 407.500000 480.350000 408.500000 481.650000 ;
      RECT 372.500000 480.350000 399.500000 481.650000 ;
      RECT 357.500000 480.350000 359.500000 481.650000 ;
      RECT 316.500000 480.350000 349.500000 481.650000 ;
      RECT 307.500000 480.350000 308.500000 481.650000 ;
      RECT 266.500000 480.350000 299.500000 481.650000 ;
      RECT 257.500000 480.350000 258.500000 481.650000 ;
      RECT 216.500000 480.350000 249.500000 481.650000 ;
      RECT 207.500000 480.350000 208.500000 481.650000 ;
      RECT 166.500000 480.350000 199.500000 481.650000 ;
      RECT 157.500000 480.350000 158.500000 481.650000 ;
      RECT 116.500000 480.350000 149.500000 481.650000 ;
      RECT 107.500000 480.350000 108.500000 481.650000 ;
      RECT 66.500000 480.350000 99.500000 481.650000 ;
      RECT 57.500000 480.350000 58.500000 481.650000 ;
      RECT 29.500000 480.350000 49.500000 481.650000 ;
      RECT 15.500000 480.350000 16.500000 481.650000 ;
      RECT 0.000000 480.350000 2.500000 483.650000 ;
      RECT 1139.000000 479.650000 1158.500000 480.350000 ;
      RECT 722.500000 479.650000 739.000000 480.350000 ;
      RECT 666.500000 479.650000 708.500000 480.350000 ;
      RECT 616.500000 479.650000 658.500000 480.350000 ;
      RECT 566.500000 479.650000 608.500000 480.350000 ;
      RECT 516.500000 479.650000 558.500000 480.350000 ;
      RECT 466.500000 479.650000 508.500000 480.350000 ;
      RECT 416.500000 479.650000 458.500000 480.350000 ;
      RECT 372.500000 479.650000 408.500000 480.350000 ;
      RECT 316.500000 479.650000 359.500000 480.350000 ;
      RECT 266.500000 479.650000 308.500000 480.350000 ;
      RECT 216.500000 479.650000 258.500000 480.350000 ;
      RECT 166.500000 479.650000 208.500000 480.350000 ;
      RECT 116.500000 479.650000 158.500000 480.350000 ;
      RECT 66.500000 479.650000 108.500000 480.350000 ;
      RECT 29.500000 479.650000 58.500000 480.350000 ;
      RECT 0.000000 479.650000 16.500000 480.350000 ;
      RECT 1166.500000 478.350000 1186.000000 481.650000 ;
      RECT 1157.500000 478.350000 1158.500000 479.650000 ;
      RECT 722.500000 478.350000 723.500000 479.650000 ;
      RECT 707.500000 478.350000 708.500000 479.650000 ;
      RECT 666.500000 478.350000 699.500000 479.650000 ;
      RECT 657.500000 478.350000 658.500000 479.650000 ;
      RECT 616.500000 478.350000 649.500000 479.650000 ;
      RECT 607.500000 478.350000 608.500000 479.650000 ;
      RECT 566.500000 478.350000 599.500000 479.650000 ;
      RECT 557.500000 478.350000 558.500000 479.650000 ;
      RECT 516.500000 478.350000 549.500000 479.650000 ;
      RECT 507.500000 478.350000 508.500000 479.650000 ;
      RECT 466.500000 478.350000 499.500000 479.650000 ;
      RECT 457.500000 478.350000 458.500000 479.650000 ;
      RECT 416.500000 478.350000 449.500000 479.650000 ;
      RECT 407.500000 478.350000 408.500000 479.650000 ;
      RECT 372.500000 478.350000 399.500000 479.650000 ;
      RECT 357.500000 478.350000 359.500000 479.650000 ;
      RECT 316.500000 478.350000 349.500000 479.650000 ;
      RECT 307.500000 478.350000 308.500000 479.650000 ;
      RECT 266.500000 478.350000 299.500000 479.650000 ;
      RECT 257.500000 478.350000 258.500000 479.650000 ;
      RECT 216.500000 478.350000 249.500000 479.650000 ;
      RECT 207.500000 478.350000 208.500000 479.650000 ;
      RECT 166.500000 478.350000 199.500000 479.650000 ;
      RECT 157.500000 478.350000 158.500000 479.650000 ;
      RECT 116.500000 478.350000 149.500000 479.650000 ;
      RECT 107.500000 478.350000 108.500000 479.650000 ;
      RECT 66.500000 478.350000 99.500000 479.650000 ;
      RECT 57.500000 478.350000 58.500000 479.650000 ;
      RECT 29.500000 478.350000 49.500000 479.650000 ;
      RECT 15.500000 478.350000 16.500000 479.650000 ;
      RECT 1157.500000 477.650000 1186.000000 478.350000 ;
      RECT 707.500000 477.650000 723.500000 478.350000 ;
      RECT 657.500000 477.650000 699.500000 478.350000 ;
      RECT 607.500000 477.650000 649.500000 478.350000 ;
      RECT 557.500000 477.650000 599.500000 478.350000 ;
      RECT 507.500000 477.650000 549.500000 478.350000 ;
      RECT 457.500000 477.650000 499.500000 478.350000 ;
      RECT 407.500000 477.650000 449.500000 478.350000 ;
      RECT 357.500000 477.650000 399.500000 478.350000 ;
      RECT 307.500000 477.650000 349.500000 478.350000 ;
      RECT 257.500000 477.650000 299.500000 478.350000 ;
      RECT 207.500000 477.650000 249.500000 478.350000 ;
      RECT 157.500000 477.650000 199.500000 478.350000 ;
      RECT 107.500000 477.650000 149.500000 478.350000 ;
      RECT 57.500000 477.650000 99.500000 478.350000 ;
      RECT 15.500000 477.650000 49.500000 478.350000 ;
      RECT 1157.500000 476.350000 1158.500000 477.650000 ;
      RECT 1139.000000 476.350000 1149.500000 479.650000 ;
      RECT 736.500000 476.350000 739.000000 479.650000 ;
      RECT 722.500000 476.350000 723.500000 477.650000 ;
      RECT 707.500000 476.350000 708.500000 477.650000 ;
      RECT 666.500000 476.350000 699.500000 477.650000 ;
      RECT 657.500000 476.350000 658.500000 477.650000 ;
      RECT 616.500000 476.350000 649.500000 477.650000 ;
      RECT 607.500000 476.350000 608.500000 477.650000 ;
      RECT 566.500000 476.350000 599.500000 477.650000 ;
      RECT 557.500000 476.350000 558.500000 477.650000 ;
      RECT 516.500000 476.350000 549.500000 477.650000 ;
      RECT 507.500000 476.350000 508.500000 477.650000 ;
      RECT 466.500000 476.350000 499.500000 477.650000 ;
      RECT 457.500000 476.350000 458.500000 477.650000 ;
      RECT 416.500000 476.350000 449.500000 477.650000 ;
      RECT 407.500000 476.350000 408.500000 477.650000 ;
      RECT 370.000000 476.350000 399.500000 477.650000 ;
      RECT 357.500000 476.350000 362.000000 477.650000 ;
      RECT 316.500000 476.350000 349.500000 477.650000 ;
      RECT 307.500000 476.350000 308.500000 477.650000 ;
      RECT 266.500000 476.350000 299.500000 477.650000 ;
      RECT 257.500000 476.350000 258.500000 477.650000 ;
      RECT 216.500000 476.350000 249.500000 477.650000 ;
      RECT 207.500000 476.350000 208.500000 477.650000 ;
      RECT 166.500000 476.350000 199.500000 477.650000 ;
      RECT 157.500000 476.350000 158.500000 477.650000 ;
      RECT 116.500000 476.350000 149.500000 477.650000 ;
      RECT 107.500000 476.350000 108.500000 477.650000 ;
      RECT 66.500000 476.350000 99.500000 477.650000 ;
      RECT 57.500000 476.350000 58.500000 477.650000 ;
      RECT 29.500000 476.350000 49.500000 477.650000 ;
      RECT 15.500000 476.350000 16.500000 477.650000 ;
      RECT 0.000000 476.350000 2.500000 479.650000 ;
      RECT 1139.000000 475.650000 1158.500000 476.350000 ;
      RECT 722.500000 475.650000 739.000000 476.350000 ;
      RECT 666.500000 475.650000 708.500000 476.350000 ;
      RECT 616.500000 475.650000 658.500000 476.350000 ;
      RECT 566.500000 475.650000 608.500000 476.350000 ;
      RECT 516.500000 475.650000 558.500000 476.350000 ;
      RECT 466.500000 475.650000 508.500000 476.350000 ;
      RECT 416.500000 475.650000 458.500000 476.350000 ;
      RECT 370.000000 475.650000 408.500000 476.350000 ;
      RECT 316.500000 475.650000 362.000000 476.350000 ;
      RECT 266.500000 475.650000 308.500000 476.350000 ;
      RECT 216.500000 475.650000 258.500000 476.350000 ;
      RECT 166.500000 475.650000 208.500000 476.350000 ;
      RECT 116.500000 475.650000 158.500000 476.350000 ;
      RECT 66.500000 475.650000 108.500000 476.350000 ;
      RECT 29.500000 475.650000 58.500000 476.350000 ;
      RECT 0.000000 475.650000 16.500000 476.350000 ;
      RECT 1166.500000 474.350000 1186.000000 477.650000 ;
      RECT 1157.500000 474.350000 1158.500000 475.650000 ;
      RECT 722.500000 474.350000 723.500000 475.650000 ;
      RECT 707.500000 474.350000 708.500000 475.650000 ;
      RECT 666.500000 474.350000 699.500000 475.650000 ;
      RECT 657.500000 474.350000 658.500000 475.650000 ;
      RECT 616.500000 474.350000 649.500000 475.650000 ;
      RECT 607.500000 474.350000 608.500000 475.650000 ;
      RECT 566.500000 474.350000 599.500000 475.650000 ;
      RECT 557.500000 474.350000 558.500000 475.650000 ;
      RECT 516.500000 474.350000 549.500000 475.650000 ;
      RECT 507.500000 474.350000 508.500000 475.650000 ;
      RECT 466.500000 474.350000 499.500000 475.650000 ;
      RECT 457.500000 474.350000 458.500000 475.650000 ;
      RECT 416.500000 474.350000 449.500000 475.650000 ;
      RECT 407.500000 474.350000 408.500000 475.650000 ;
      RECT 370.000000 474.350000 399.500000 475.650000 ;
      RECT 357.500000 474.350000 362.000000 475.650000 ;
      RECT 316.500000 474.350000 349.500000 475.650000 ;
      RECT 307.500000 474.350000 308.500000 475.650000 ;
      RECT 266.500000 474.350000 299.500000 475.650000 ;
      RECT 257.500000 474.350000 258.500000 475.650000 ;
      RECT 216.500000 474.350000 249.500000 475.650000 ;
      RECT 207.500000 474.350000 208.500000 475.650000 ;
      RECT 166.500000 474.350000 199.500000 475.650000 ;
      RECT 157.500000 474.350000 158.500000 475.650000 ;
      RECT 116.500000 474.350000 149.500000 475.650000 ;
      RECT 107.500000 474.350000 108.500000 475.650000 ;
      RECT 66.500000 474.350000 99.500000 475.650000 ;
      RECT 57.500000 474.350000 58.500000 475.650000 ;
      RECT 29.500000 474.350000 49.500000 475.650000 ;
      RECT 15.500000 474.350000 16.500000 475.650000 ;
      RECT 1157.500000 473.650000 1186.000000 474.350000 ;
      RECT 707.500000 473.650000 723.500000 474.350000 ;
      RECT 657.500000 473.650000 699.500000 474.350000 ;
      RECT 607.500000 473.650000 649.500000 474.350000 ;
      RECT 557.500000 473.650000 599.500000 474.350000 ;
      RECT 507.500000 473.650000 549.500000 474.350000 ;
      RECT 457.500000 473.650000 499.500000 474.350000 ;
      RECT 407.500000 473.650000 449.500000 474.350000 ;
      RECT 357.500000 473.650000 399.500000 474.350000 ;
      RECT 307.500000 473.650000 349.500000 474.350000 ;
      RECT 257.500000 473.650000 299.500000 474.350000 ;
      RECT 207.500000 473.650000 249.500000 474.350000 ;
      RECT 157.500000 473.650000 199.500000 474.350000 ;
      RECT 107.500000 473.650000 149.500000 474.350000 ;
      RECT 57.500000 473.650000 99.500000 474.350000 ;
      RECT 15.500000 473.650000 49.500000 474.350000 ;
      RECT 1157.500000 472.350000 1158.500000 473.650000 ;
      RECT 1139.000000 472.350000 1149.500000 475.650000 ;
      RECT 736.500000 472.350000 739.000000 475.650000 ;
      RECT 722.500000 472.350000 723.500000 473.650000 ;
      RECT 707.500000 472.350000 708.500000 473.650000 ;
      RECT 666.500000 472.350000 699.500000 473.650000 ;
      RECT 657.500000 472.350000 658.500000 473.650000 ;
      RECT 616.500000 472.350000 649.500000 473.650000 ;
      RECT 607.500000 472.350000 608.500000 473.650000 ;
      RECT 566.500000 472.350000 599.500000 473.650000 ;
      RECT 557.500000 472.350000 558.500000 473.650000 ;
      RECT 516.500000 472.350000 549.500000 473.650000 ;
      RECT 507.500000 472.350000 508.500000 473.650000 ;
      RECT 466.500000 472.350000 499.500000 473.650000 ;
      RECT 457.500000 472.350000 458.500000 473.650000 ;
      RECT 416.500000 472.350000 449.500000 473.650000 ;
      RECT 407.500000 472.350000 408.500000 473.650000 ;
      RECT 370.000000 472.350000 399.500000 473.650000 ;
      RECT 357.500000 472.350000 358.500000 473.650000 ;
      RECT 316.500000 472.350000 349.500000 473.650000 ;
      RECT 307.500000 472.350000 308.500000 473.650000 ;
      RECT 266.500000 472.350000 299.500000 473.650000 ;
      RECT 257.500000 472.350000 258.500000 473.650000 ;
      RECT 216.500000 472.350000 249.500000 473.650000 ;
      RECT 207.500000 472.350000 208.500000 473.650000 ;
      RECT 166.500000 472.350000 199.500000 473.650000 ;
      RECT 157.500000 472.350000 158.500000 473.650000 ;
      RECT 116.500000 472.350000 149.500000 473.650000 ;
      RECT 107.500000 472.350000 108.500000 473.650000 ;
      RECT 66.500000 472.350000 99.500000 473.650000 ;
      RECT 57.500000 472.350000 58.500000 473.650000 ;
      RECT 29.500000 472.350000 49.500000 473.650000 ;
      RECT 15.500000 472.350000 16.500000 473.650000 ;
      RECT 0.000000 472.350000 2.500000 475.650000 ;
      RECT 1139.000000 471.650000 1158.500000 472.350000 ;
      RECT 722.500000 471.650000 739.000000 472.350000 ;
      RECT 666.500000 471.650000 708.500000 472.350000 ;
      RECT 616.500000 471.650000 658.500000 472.350000 ;
      RECT 566.500000 471.650000 608.500000 472.350000 ;
      RECT 516.500000 471.650000 558.500000 472.350000 ;
      RECT 466.500000 471.650000 508.500000 472.350000 ;
      RECT 416.500000 471.650000 458.500000 472.350000 ;
      RECT 370.000000 471.650000 408.500000 472.350000 ;
      RECT 316.500000 471.650000 358.500000 472.350000 ;
      RECT 266.500000 471.650000 308.500000 472.350000 ;
      RECT 216.500000 471.650000 258.500000 472.350000 ;
      RECT 166.500000 471.650000 208.500000 472.350000 ;
      RECT 116.500000 471.650000 158.500000 472.350000 ;
      RECT 66.500000 471.650000 108.500000 472.350000 ;
      RECT 29.500000 471.650000 58.500000 472.350000 ;
      RECT 0.000000 471.650000 16.500000 472.350000 ;
      RECT 1166.500000 470.350000 1186.000000 473.650000 ;
      RECT 1157.500000 470.350000 1158.500000 471.650000 ;
      RECT 722.500000 470.350000 723.500000 471.650000 ;
      RECT 707.500000 470.350000 708.500000 471.650000 ;
      RECT 666.500000 470.350000 699.500000 471.650000 ;
      RECT 657.500000 470.350000 658.500000 471.650000 ;
      RECT 616.500000 470.350000 649.500000 471.650000 ;
      RECT 607.500000 470.350000 608.500000 471.650000 ;
      RECT 566.500000 470.350000 599.500000 471.650000 ;
      RECT 557.500000 470.350000 558.500000 471.650000 ;
      RECT 516.500000 470.350000 549.500000 471.650000 ;
      RECT 507.500000 470.350000 508.500000 471.650000 ;
      RECT 466.500000 470.350000 499.500000 471.650000 ;
      RECT 457.500000 470.350000 458.500000 471.650000 ;
      RECT 416.500000 470.350000 449.500000 471.650000 ;
      RECT 407.500000 470.350000 408.500000 471.650000 ;
      RECT 370.000000 470.350000 399.500000 471.650000 ;
      RECT 357.500000 470.350000 358.500000 471.650000 ;
      RECT 316.500000 470.350000 349.500000 471.650000 ;
      RECT 307.500000 470.350000 308.500000 471.650000 ;
      RECT 266.500000 470.350000 299.500000 471.650000 ;
      RECT 257.500000 470.350000 258.500000 471.650000 ;
      RECT 216.500000 470.350000 249.500000 471.650000 ;
      RECT 207.500000 470.350000 208.500000 471.650000 ;
      RECT 166.500000 470.350000 199.500000 471.650000 ;
      RECT 157.500000 470.350000 158.500000 471.650000 ;
      RECT 116.500000 470.350000 149.500000 471.650000 ;
      RECT 107.500000 470.350000 108.500000 471.650000 ;
      RECT 66.500000 470.350000 99.500000 471.650000 ;
      RECT 57.500000 470.350000 58.500000 471.650000 ;
      RECT 29.500000 470.350000 49.500000 471.650000 ;
      RECT 15.500000 470.350000 16.500000 471.650000 ;
      RECT 1157.500000 469.650000 1186.000000 470.350000 ;
      RECT 707.500000 469.650000 723.500000 470.350000 ;
      RECT 657.500000 469.650000 699.500000 470.350000 ;
      RECT 607.500000 469.650000 649.500000 470.350000 ;
      RECT 557.500000 469.650000 599.500000 470.350000 ;
      RECT 507.500000 469.650000 549.500000 470.350000 ;
      RECT 457.500000 469.650000 499.500000 470.350000 ;
      RECT 407.500000 469.650000 449.500000 470.350000 ;
      RECT 357.500000 469.650000 399.500000 470.350000 ;
      RECT 307.500000 469.650000 349.500000 470.350000 ;
      RECT 257.500000 469.650000 299.500000 470.350000 ;
      RECT 207.500000 469.650000 249.500000 470.350000 ;
      RECT 157.500000 469.650000 199.500000 470.350000 ;
      RECT 107.500000 469.650000 149.500000 470.350000 ;
      RECT 57.500000 469.650000 99.500000 470.350000 ;
      RECT 15.500000 469.650000 49.500000 470.350000 ;
      RECT 1157.500000 468.350000 1158.500000 469.650000 ;
      RECT 1139.000000 468.350000 1149.500000 471.650000 ;
      RECT 736.500000 468.350000 739.000000 471.650000 ;
      RECT 722.500000 468.350000 723.500000 469.650000 ;
      RECT 707.500000 468.350000 708.500000 469.650000 ;
      RECT 666.500000 468.350000 699.500000 469.650000 ;
      RECT 657.500000 468.350000 658.500000 469.650000 ;
      RECT 616.500000 468.350000 649.500000 469.650000 ;
      RECT 607.500000 468.350000 608.500000 469.650000 ;
      RECT 566.500000 468.350000 599.500000 469.650000 ;
      RECT 557.500000 468.350000 558.500000 469.650000 ;
      RECT 516.500000 468.350000 549.500000 469.650000 ;
      RECT 507.500000 468.350000 508.500000 469.650000 ;
      RECT 466.500000 468.350000 499.500000 469.650000 ;
      RECT 457.500000 468.350000 458.500000 469.650000 ;
      RECT 416.500000 468.350000 449.500000 469.650000 ;
      RECT 407.500000 468.350000 408.500000 469.650000 ;
      RECT 366.500000 468.350000 399.500000 469.650000 ;
      RECT 357.500000 468.350000 358.500000 469.650000 ;
      RECT 316.500000 468.350000 349.500000 469.650000 ;
      RECT 307.500000 468.350000 308.500000 469.650000 ;
      RECT 266.500000 468.350000 299.500000 469.650000 ;
      RECT 257.500000 468.350000 258.500000 469.650000 ;
      RECT 216.500000 468.350000 249.500000 469.650000 ;
      RECT 207.500000 468.350000 208.500000 469.650000 ;
      RECT 166.500000 468.350000 199.500000 469.650000 ;
      RECT 157.500000 468.350000 158.500000 469.650000 ;
      RECT 116.500000 468.350000 149.500000 469.650000 ;
      RECT 107.500000 468.350000 108.500000 469.650000 ;
      RECT 66.500000 468.350000 99.500000 469.650000 ;
      RECT 57.500000 468.350000 58.500000 469.650000 ;
      RECT 29.500000 468.350000 49.500000 469.650000 ;
      RECT 15.500000 468.350000 16.500000 469.650000 ;
      RECT 0.000000 468.350000 2.500000 471.650000 ;
      RECT 1139.000000 467.650000 1158.500000 468.350000 ;
      RECT 722.500000 467.650000 739.000000 468.350000 ;
      RECT 666.500000 467.650000 708.500000 468.350000 ;
      RECT 616.500000 467.650000 658.500000 468.350000 ;
      RECT 566.500000 467.650000 608.500000 468.350000 ;
      RECT 516.500000 467.650000 558.500000 468.350000 ;
      RECT 466.500000 467.650000 508.500000 468.350000 ;
      RECT 416.500000 467.650000 458.500000 468.350000 ;
      RECT 366.500000 467.650000 408.500000 468.350000 ;
      RECT 316.500000 467.650000 358.500000 468.350000 ;
      RECT 266.500000 467.650000 308.500000 468.350000 ;
      RECT 216.500000 467.650000 258.500000 468.350000 ;
      RECT 166.500000 467.650000 208.500000 468.350000 ;
      RECT 116.500000 467.650000 158.500000 468.350000 ;
      RECT 66.500000 467.650000 108.500000 468.350000 ;
      RECT 29.500000 467.650000 58.500000 468.350000 ;
      RECT 0.000000 467.650000 16.500000 468.350000 ;
      RECT 1166.500000 466.350000 1186.000000 469.650000 ;
      RECT 1157.500000 466.350000 1158.500000 467.650000 ;
      RECT 722.500000 466.350000 723.500000 467.650000 ;
      RECT 707.500000 466.350000 708.500000 467.650000 ;
      RECT 666.500000 466.350000 699.500000 467.650000 ;
      RECT 657.500000 466.350000 658.500000 467.650000 ;
      RECT 616.500000 466.350000 649.500000 467.650000 ;
      RECT 607.500000 466.350000 608.500000 467.650000 ;
      RECT 566.500000 466.350000 599.500000 467.650000 ;
      RECT 557.500000 466.350000 558.500000 467.650000 ;
      RECT 516.500000 466.350000 549.500000 467.650000 ;
      RECT 507.500000 466.350000 508.500000 467.650000 ;
      RECT 466.500000 466.350000 499.500000 467.650000 ;
      RECT 457.500000 466.350000 458.500000 467.650000 ;
      RECT 416.500000 466.350000 449.500000 467.650000 ;
      RECT 407.500000 466.350000 408.500000 467.650000 ;
      RECT 366.500000 466.350000 399.500000 467.650000 ;
      RECT 357.500000 466.350000 358.500000 467.650000 ;
      RECT 316.500000 466.350000 349.500000 467.650000 ;
      RECT 307.500000 466.350000 308.500000 467.650000 ;
      RECT 266.500000 466.350000 299.500000 467.650000 ;
      RECT 257.500000 466.350000 258.500000 467.650000 ;
      RECT 216.500000 466.350000 249.500000 467.650000 ;
      RECT 207.500000 466.350000 208.500000 467.650000 ;
      RECT 166.500000 466.350000 199.500000 467.650000 ;
      RECT 157.500000 466.350000 158.500000 467.650000 ;
      RECT 116.500000 466.350000 149.500000 467.650000 ;
      RECT 107.500000 466.350000 108.500000 467.650000 ;
      RECT 66.500000 466.350000 99.500000 467.650000 ;
      RECT 57.500000 466.350000 58.500000 467.650000 ;
      RECT 29.500000 466.350000 49.500000 467.650000 ;
      RECT 15.500000 466.350000 16.500000 467.650000 ;
      RECT 1157.500000 465.650000 1186.000000 466.350000 ;
      RECT 707.500000 465.650000 723.500000 466.350000 ;
      RECT 657.500000 465.650000 699.500000 466.350000 ;
      RECT 607.500000 465.650000 649.500000 466.350000 ;
      RECT 557.500000 465.650000 599.500000 466.350000 ;
      RECT 507.500000 465.650000 549.500000 466.350000 ;
      RECT 457.500000 465.650000 499.500000 466.350000 ;
      RECT 407.500000 465.650000 449.500000 466.350000 ;
      RECT 357.500000 465.650000 399.500000 466.350000 ;
      RECT 307.500000 465.650000 349.500000 466.350000 ;
      RECT 257.500000 465.650000 299.500000 466.350000 ;
      RECT 207.500000 465.650000 249.500000 466.350000 ;
      RECT 157.500000 465.650000 199.500000 466.350000 ;
      RECT 107.500000 465.650000 149.500000 466.350000 ;
      RECT 57.500000 465.650000 99.500000 466.350000 ;
      RECT 15.500000 465.650000 49.500000 466.350000 ;
      RECT 1157.500000 464.350000 1158.500000 465.650000 ;
      RECT 1139.000000 464.350000 1149.500000 467.650000 ;
      RECT 736.500000 464.350000 739.000000 467.650000 ;
      RECT 722.500000 464.350000 723.500000 465.650000 ;
      RECT 707.500000 464.350000 708.500000 465.650000 ;
      RECT 666.500000 464.350000 699.500000 465.650000 ;
      RECT 657.500000 464.350000 658.500000 465.650000 ;
      RECT 616.500000 464.350000 649.500000 465.650000 ;
      RECT 607.500000 464.350000 608.500000 465.650000 ;
      RECT 566.500000 464.350000 599.500000 465.650000 ;
      RECT 557.500000 464.350000 558.500000 465.650000 ;
      RECT 516.500000 464.350000 549.500000 465.650000 ;
      RECT 507.500000 464.350000 508.500000 465.650000 ;
      RECT 466.500000 464.350000 499.500000 465.650000 ;
      RECT 457.500000 464.350000 458.500000 465.650000 ;
      RECT 416.500000 464.350000 449.500000 465.650000 ;
      RECT 407.500000 464.350000 408.500000 465.650000 ;
      RECT 366.500000 464.350000 399.500000 465.650000 ;
      RECT 357.500000 464.350000 358.500000 465.650000 ;
      RECT 316.500000 464.350000 349.500000 465.650000 ;
      RECT 307.500000 464.350000 308.500000 465.650000 ;
      RECT 266.500000 464.350000 299.500000 465.650000 ;
      RECT 257.500000 464.350000 258.500000 465.650000 ;
      RECT 216.500000 464.350000 249.500000 465.650000 ;
      RECT 207.500000 464.350000 208.500000 465.650000 ;
      RECT 166.500000 464.350000 199.500000 465.650000 ;
      RECT 157.500000 464.350000 158.500000 465.650000 ;
      RECT 116.500000 464.350000 149.500000 465.650000 ;
      RECT 107.500000 464.350000 108.500000 465.650000 ;
      RECT 66.500000 464.350000 99.500000 465.650000 ;
      RECT 57.500000 464.350000 58.500000 465.650000 ;
      RECT 29.500000 464.350000 49.500000 465.650000 ;
      RECT 15.500000 464.350000 16.500000 465.650000 ;
      RECT 0.000000 464.350000 2.500000 467.650000 ;
      RECT 1139.000000 463.650000 1158.500000 464.350000 ;
      RECT 722.500000 463.650000 739.000000 464.350000 ;
      RECT 666.500000 463.650000 708.500000 464.350000 ;
      RECT 616.500000 463.650000 658.500000 464.350000 ;
      RECT 566.500000 463.650000 608.500000 464.350000 ;
      RECT 516.500000 463.650000 558.500000 464.350000 ;
      RECT 466.500000 463.650000 508.500000 464.350000 ;
      RECT 416.500000 463.650000 458.500000 464.350000 ;
      RECT 366.500000 463.650000 408.500000 464.350000 ;
      RECT 316.500000 463.650000 358.500000 464.350000 ;
      RECT 266.500000 463.650000 308.500000 464.350000 ;
      RECT 216.500000 463.650000 258.500000 464.350000 ;
      RECT 166.500000 463.650000 208.500000 464.350000 ;
      RECT 116.500000 463.650000 158.500000 464.350000 ;
      RECT 66.500000 463.650000 108.500000 464.350000 ;
      RECT 29.500000 463.650000 58.500000 464.350000 ;
      RECT 0.000000 463.650000 16.500000 464.350000 ;
      RECT 1166.500000 462.350000 1186.000000 465.650000 ;
      RECT 1157.500000 462.350000 1158.500000 463.650000 ;
      RECT 722.500000 462.350000 723.500000 463.650000 ;
      RECT 707.500000 462.350000 708.500000 463.650000 ;
      RECT 666.500000 462.350000 699.500000 463.650000 ;
      RECT 657.500000 462.350000 658.500000 463.650000 ;
      RECT 616.500000 462.350000 649.500000 463.650000 ;
      RECT 607.500000 462.350000 608.500000 463.650000 ;
      RECT 566.500000 462.350000 599.500000 463.650000 ;
      RECT 557.500000 462.350000 558.500000 463.650000 ;
      RECT 516.500000 462.350000 549.500000 463.650000 ;
      RECT 507.500000 462.350000 508.500000 463.650000 ;
      RECT 466.500000 462.350000 499.500000 463.650000 ;
      RECT 457.500000 462.350000 458.500000 463.650000 ;
      RECT 416.500000 462.350000 449.500000 463.650000 ;
      RECT 407.500000 462.350000 408.500000 463.650000 ;
      RECT 366.500000 462.350000 399.500000 463.650000 ;
      RECT 357.500000 462.350000 358.500000 463.650000 ;
      RECT 316.500000 462.350000 349.500000 463.650000 ;
      RECT 307.500000 462.350000 308.500000 463.650000 ;
      RECT 266.500000 462.350000 299.500000 463.650000 ;
      RECT 257.500000 462.350000 258.500000 463.650000 ;
      RECT 216.500000 462.350000 249.500000 463.650000 ;
      RECT 207.500000 462.350000 208.500000 463.650000 ;
      RECT 166.500000 462.350000 199.500000 463.650000 ;
      RECT 157.500000 462.350000 158.500000 463.650000 ;
      RECT 116.500000 462.350000 149.500000 463.650000 ;
      RECT 107.500000 462.350000 108.500000 463.650000 ;
      RECT 66.500000 462.350000 99.500000 463.650000 ;
      RECT 57.500000 462.350000 58.500000 463.650000 ;
      RECT 29.500000 462.350000 49.500000 463.650000 ;
      RECT 15.500000 462.350000 16.500000 463.650000 ;
      RECT 1157.500000 461.650000 1186.000000 462.350000 ;
      RECT 707.500000 461.650000 723.500000 462.350000 ;
      RECT 657.500000 461.650000 699.500000 462.350000 ;
      RECT 607.500000 461.650000 649.500000 462.350000 ;
      RECT 557.500000 461.650000 599.500000 462.350000 ;
      RECT 507.500000 461.650000 549.500000 462.350000 ;
      RECT 457.500000 461.650000 499.500000 462.350000 ;
      RECT 407.500000 461.650000 449.500000 462.350000 ;
      RECT 357.500000 461.650000 399.500000 462.350000 ;
      RECT 307.500000 461.650000 349.500000 462.350000 ;
      RECT 207.500000 461.650000 249.500000 462.350000 ;
      RECT 107.500000 461.650000 149.500000 462.350000 ;
      RECT 57.500000 461.650000 99.500000 462.350000 ;
      RECT 15.500000 461.650000 49.500000 462.350000 ;
      RECT 1157.500000 460.350000 1158.500000 461.650000 ;
      RECT 1139.000000 460.350000 1149.500000 463.650000 ;
      RECT 736.500000 460.350000 739.000000 463.650000 ;
      RECT 722.500000 460.350000 723.500000 461.650000 ;
      RECT 707.500000 460.350000 708.500000 461.650000 ;
      RECT 666.500000 460.350000 699.500000 461.650000 ;
      RECT 657.500000 460.350000 658.500000 461.650000 ;
      RECT 616.500000 460.350000 649.500000 461.650000 ;
      RECT 607.500000 460.350000 608.500000 461.650000 ;
      RECT 566.500000 460.350000 599.500000 461.650000 ;
      RECT 557.500000 460.350000 558.500000 461.650000 ;
      RECT 516.500000 460.350000 549.500000 461.650000 ;
      RECT 507.500000 460.350000 508.500000 461.650000 ;
      RECT 466.500000 460.350000 499.500000 461.650000 ;
      RECT 457.500000 460.350000 458.500000 461.650000 ;
      RECT 416.500000 460.350000 449.500000 461.650000 ;
      RECT 407.500000 460.350000 408.500000 461.650000 ;
      RECT 366.500000 460.350000 399.500000 461.650000 ;
      RECT 357.500000 460.350000 358.500000 461.650000 ;
      RECT 316.500000 460.350000 349.500000 461.650000 ;
      RECT 307.500000 460.350000 308.500000 461.650000 ;
      RECT 257.500000 460.350000 299.500000 462.350000 ;
      RECT 216.500000 460.350000 249.500000 461.650000 ;
      RECT 207.500000 460.350000 208.500000 461.650000 ;
      RECT 157.500000 460.350000 199.500000 462.350000 ;
      RECT 116.500000 460.350000 149.500000 461.650000 ;
      RECT 107.500000 460.350000 108.500000 461.650000 ;
      RECT 66.500000 460.350000 99.500000 461.650000 ;
      RECT 57.500000 460.350000 58.500000 461.650000 ;
      RECT 29.500000 460.350000 49.500000 461.650000 ;
      RECT 15.500000 460.350000 16.500000 461.650000 ;
      RECT 0.000000 460.350000 2.500000 463.650000 ;
      RECT 1139.000000 459.650000 1158.500000 460.350000 ;
      RECT 722.500000 459.650000 739.000000 460.350000 ;
      RECT 666.500000 459.650000 708.500000 460.350000 ;
      RECT 616.500000 459.650000 658.500000 460.350000 ;
      RECT 566.500000 459.650000 608.500000 460.350000 ;
      RECT 516.500000 459.650000 558.500000 460.350000 ;
      RECT 466.500000 459.650000 508.500000 460.350000 ;
      RECT 416.500000 459.650000 458.500000 460.350000 ;
      RECT 366.500000 459.650000 408.500000 460.350000 ;
      RECT 316.500000 459.650000 358.500000 460.350000 ;
      RECT 216.500000 459.650000 308.500000 460.350000 ;
      RECT 116.500000 459.650000 208.500000 460.350000 ;
      RECT 66.500000 459.650000 108.500000 460.350000 ;
      RECT 29.500000 459.650000 58.500000 460.350000 ;
      RECT 0.000000 459.650000 16.500000 460.350000 ;
      RECT 1166.500000 458.350000 1186.000000 461.650000 ;
      RECT 1157.500000 458.350000 1158.500000 459.650000 ;
      RECT 722.500000 458.350000 723.500000 459.650000 ;
      RECT 707.500000 458.350000 708.500000 459.650000 ;
      RECT 666.500000 458.350000 699.500000 459.650000 ;
      RECT 657.500000 458.350000 658.500000 459.650000 ;
      RECT 616.500000 458.350000 649.500000 459.650000 ;
      RECT 607.500000 458.350000 608.500000 459.650000 ;
      RECT 566.500000 458.350000 599.500000 459.650000 ;
      RECT 557.500000 458.350000 558.500000 459.650000 ;
      RECT 516.500000 458.350000 549.500000 459.650000 ;
      RECT 507.500000 458.350000 508.500000 459.650000 ;
      RECT 466.500000 458.350000 499.500000 459.650000 ;
      RECT 457.500000 458.350000 458.500000 459.650000 ;
      RECT 416.500000 458.350000 449.500000 459.650000 ;
      RECT 407.500000 458.350000 408.500000 459.650000 ;
      RECT 366.500000 458.350000 399.500000 459.650000 ;
      RECT 357.500000 458.350000 358.500000 459.650000 ;
      RECT 316.500000 458.350000 349.500000 459.650000 ;
      RECT 307.500000 458.350000 308.500000 459.650000 ;
      RECT 216.500000 458.350000 249.500000 459.650000 ;
      RECT 207.500000 458.350000 208.500000 459.650000 ;
      RECT 116.500000 458.350000 149.500000 459.650000 ;
      RECT 107.500000 458.350000 108.500000 459.650000 ;
      RECT 66.500000 458.350000 99.500000 459.650000 ;
      RECT 57.500000 458.350000 58.500000 459.650000 ;
      RECT 29.500000 458.350000 49.500000 459.650000 ;
      RECT 15.500000 458.350000 16.500000 459.650000 ;
      RECT 1157.500000 457.650000 1186.000000 458.350000 ;
      RECT 707.500000 457.650000 723.500000 458.350000 ;
      RECT 657.500000 457.650000 699.500000 458.350000 ;
      RECT 607.500000 457.650000 649.500000 458.350000 ;
      RECT 557.500000 457.650000 599.500000 458.350000 ;
      RECT 507.500000 457.650000 549.500000 458.350000 ;
      RECT 457.500000 457.650000 499.500000 458.350000 ;
      RECT 407.500000 457.650000 449.500000 458.350000 ;
      RECT 357.500000 457.650000 399.500000 458.350000 ;
      RECT 307.500000 457.650000 349.500000 458.350000 ;
      RECT 207.500000 457.650000 249.500000 458.350000 ;
      RECT 107.500000 457.650000 149.500000 458.350000 ;
      RECT 57.500000 457.650000 99.500000 458.350000 ;
      RECT 15.500000 457.650000 49.500000 458.350000 ;
      RECT 1157.500000 456.350000 1158.500000 457.650000 ;
      RECT 1139.000000 456.350000 1149.500000 459.650000 ;
      RECT 736.500000 456.350000 739.000000 459.650000 ;
      RECT 722.500000 456.350000 723.500000 457.650000 ;
      RECT 707.500000 456.350000 708.500000 457.650000 ;
      RECT 666.500000 456.350000 699.500000 457.650000 ;
      RECT 657.500000 456.350000 658.500000 457.650000 ;
      RECT 616.500000 456.350000 649.500000 457.650000 ;
      RECT 607.500000 456.350000 608.500000 457.650000 ;
      RECT 566.500000 456.350000 599.500000 457.650000 ;
      RECT 557.500000 456.350000 558.500000 457.650000 ;
      RECT 516.500000 456.350000 549.500000 457.650000 ;
      RECT 507.500000 456.350000 508.500000 457.650000 ;
      RECT 466.500000 456.350000 499.500000 457.650000 ;
      RECT 457.500000 456.350000 458.500000 457.650000 ;
      RECT 416.500000 456.350000 449.500000 457.650000 ;
      RECT 407.500000 456.350000 408.500000 457.650000 ;
      RECT 366.500000 456.350000 399.500000 457.650000 ;
      RECT 357.500000 456.350000 358.500000 457.650000 ;
      RECT 316.500000 456.350000 349.500000 457.650000 ;
      RECT 307.500000 456.350000 308.500000 457.650000 ;
      RECT 257.500000 456.350000 299.500000 459.650000 ;
      RECT 216.500000 456.350000 249.500000 457.650000 ;
      RECT 207.500000 456.350000 208.500000 457.650000 ;
      RECT 157.500000 456.350000 199.500000 459.650000 ;
      RECT 116.500000 456.350000 149.500000 457.650000 ;
      RECT 107.500000 456.350000 108.500000 457.650000 ;
      RECT 66.500000 456.350000 99.500000 457.650000 ;
      RECT 57.500000 456.350000 58.500000 457.650000 ;
      RECT 29.500000 456.350000 49.500000 457.650000 ;
      RECT 15.500000 456.350000 16.500000 457.650000 ;
      RECT 0.000000 456.350000 2.500000 459.650000 ;
      RECT 1139.000000 455.650000 1158.500000 456.350000 ;
      RECT 722.500000 455.650000 739.000000 456.350000 ;
      RECT 666.500000 455.650000 708.500000 456.350000 ;
      RECT 616.500000 455.650000 658.500000 456.350000 ;
      RECT 566.500000 455.650000 608.500000 456.350000 ;
      RECT 516.500000 455.650000 558.500000 456.350000 ;
      RECT 466.500000 455.650000 508.500000 456.350000 ;
      RECT 416.500000 455.650000 458.500000 456.350000 ;
      RECT 366.500000 455.650000 408.500000 456.350000 ;
      RECT 316.500000 455.650000 358.500000 456.350000 ;
      RECT 216.500000 455.650000 308.500000 456.350000 ;
      RECT 116.500000 455.650000 208.500000 456.350000 ;
      RECT 66.500000 455.650000 108.500000 456.350000 ;
      RECT 29.500000 455.650000 58.500000 456.350000 ;
      RECT 0.000000 455.650000 16.500000 456.350000 ;
      RECT 1166.500000 454.350000 1186.000000 457.650000 ;
      RECT 1157.500000 454.350000 1158.500000 455.650000 ;
      RECT 722.500000 454.350000 723.500000 455.650000 ;
      RECT 707.500000 454.350000 708.500000 455.650000 ;
      RECT 666.500000 454.350000 699.500000 455.650000 ;
      RECT 657.500000 454.350000 658.500000 455.650000 ;
      RECT 616.500000 454.350000 649.500000 455.650000 ;
      RECT 607.500000 454.350000 608.500000 455.650000 ;
      RECT 566.500000 454.350000 599.500000 455.650000 ;
      RECT 557.500000 454.350000 558.500000 455.650000 ;
      RECT 516.500000 454.350000 549.500000 455.650000 ;
      RECT 507.500000 454.350000 508.500000 455.650000 ;
      RECT 466.500000 454.350000 499.500000 455.650000 ;
      RECT 457.500000 454.350000 458.500000 455.650000 ;
      RECT 416.500000 454.350000 449.500000 455.650000 ;
      RECT 407.500000 454.350000 408.500000 455.650000 ;
      RECT 366.500000 454.350000 399.500000 455.650000 ;
      RECT 357.500000 454.350000 358.500000 455.650000 ;
      RECT 316.500000 454.350000 349.500000 455.650000 ;
      RECT 307.500000 454.350000 308.500000 455.650000 ;
      RECT 216.500000 454.350000 249.500000 455.650000 ;
      RECT 207.500000 454.350000 208.500000 455.650000 ;
      RECT 116.500000 454.350000 149.500000 455.650000 ;
      RECT 107.500000 454.350000 108.500000 455.650000 ;
      RECT 66.500000 454.350000 99.500000 455.650000 ;
      RECT 57.500000 454.350000 58.500000 455.650000 ;
      RECT 29.500000 454.350000 49.500000 455.650000 ;
      RECT 15.500000 454.350000 16.500000 455.650000 ;
      RECT 1157.500000 453.650000 1186.000000 454.350000 ;
      RECT 707.500000 453.650000 723.500000 454.350000 ;
      RECT 657.500000 453.650000 699.500000 454.350000 ;
      RECT 607.500000 453.650000 649.500000 454.350000 ;
      RECT 557.500000 453.650000 599.500000 454.350000 ;
      RECT 507.500000 453.650000 549.500000 454.350000 ;
      RECT 457.500000 453.650000 499.500000 454.350000 ;
      RECT 407.500000 453.650000 449.500000 454.350000 ;
      RECT 357.500000 453.650000 399.500000 454.350000 ;
      RECT 307.500000 453.650000 349.500000 454.350000 ;
      RECT 207.500000 453.650000 249.500000 454.350000 ;
      RECT 107.500000 453.650000 149.500000 454.350000 ;
      RECT 57.500000 453.650000 99.500000 454.350000 ;
      RECT 15.500000 453.650000 49.500000 454.350000 ;
      RECT 1157.500000 452.350000 1158.500000 453.650000 ;
      RECT 1139.000000 452.350000 1149.500000 455.650000 ;
      RECT 736.500000 452.350000 739.000000 455.650000 ;
      RECT 722.500000 452.350000 723.500000 453.650000 ;
      RECT 707.500000 452.350000 708.500000 453.650000 ;
      RECT 666.500000 452.350000 699.500000 453.650000 ;
      RECT 657.500000 452.350000 658.500000 453.650000 ;
      RECT 616.500000 452.350000 649.500000 453.650000 ;
      RECT 607.500000 452.350000 608.500000 453.650000 ;
      RECT 566.500000 452.350000 599.500000 453.650000 ;
      RECT 557.500000 452.350000 558.500000 453.650000 ;
      RECT 516.500000 452.350000 549.500000 453.650000 ;
      RECT 507.500000 452.350000 508.500000 453.650000 ;
      RECT 466.500000 452.350000 499.500000 453.650000 ;
      RECT 457.500000 452.350000 458.500000 453.650000 ;
      RECT 416.500000 452.350000 449.500000 453.650000 ;
      RECT 407.500000 452.350000 408.500000 453.650000 ;
      RECT 366.500000 452.350000 399.500000 453.650000 ;
      RECT 357.500000 452.350000 358.500000 453.650000 ;
      RECT 316.500000 452.350000 349.500000 453.650000 ;
      RECT 307.500000 452.350000 308.500000 453.650000 ;
      RECT 257.500000 452.350000 299.500000 455.650000 ;
      RECT 216.500000 452.350000 249.500000 453.650000 ;
      RECT 207.500000 452.350000 208.500000 453.650000 ;
      RECT 157.500000 452.350000 199.500000 455.650000 ;
      RECT 116.500000 452.350000 149.500000 453.650000 ;
      RECT 107.500000 452.350000 108.500000 453.650000 ;
      RECT 66.500000 452.350000 99.500000 453.650000 ;
      RECT 57.500000 452.350000 58.500000 453.650000 ;
      RECT 29.500000 452.350000 49.500000 453.650000 ;
      RECT 15.500000 452.350000 16.500000 453.650000 ;
      RECT 0.000000 452.350000 2.500000 455.650000 ;
      RECT 1139.000000 451.650000 1158.500000 452.350000 ;
      RECT 722.500000 451.650000 739.000000 452.350000 ;
      RECT 666.500000 451.650000 708.500000 452.350000 ;
      RECT 616.500000 451.650000 658.500000 452.350000 ;
      RECT 566.500000 451.650000 608.500000 452.350000 ;
      RECT 516.500000 451.650000 558.500000 452.350000 ;
      RECT 466.500000 451.650000 508.500000 452.350000 ;
      RECT 416.500000 451.650000 458.500000 452.350000 ;
      RECT 366.500000 451.650000 408.500000 452.350000 ;
      RECT 316.500000 451.650000 358.500000 452.350000 ;
      RECT 216.500000 451.650000 308.500000 452.350000 ;
      RECT 116.500000 451.650000 208.500000 452.350000 ;
      RECT 66.500000 451.650000 108.500000 452.350000 ;
      RECT 29.500000 451.650000 58.500000 452.350000 ;
      RECT 0.000000 451.650000 16.500000 452.350000 ;
      RECT 1166.500000 450.350000 1186.000000 453.650000 ;
      RECT 1157.500000 450.350000 1158.500000 451.650000 ;
      RECT 722.500000 450.350000 723.500000 451.650000 ;
      RECT 707.500000 450.350000 708.500000 451.650000 ;
      RECT 666.500000 450.350000 699.500000 451.650000 ;
      RECT 657.500000 450.350000 658.500000 451.650000 ;
      RECT 616.500000 450.350000 649.500000 451.650000 ;
      RECT 607.500000 450.350000 608.500000 451.650000 ;
      RECT 566.500000 450.350000 599.500000 451.650000 ;
      RECT 557.500000 450.350000 558.500000 451.650000 ;
      RECT 516.500000 450.350000 549.500000 451.650000 ;
      RECT 507.500000 450.350000 508.500000 451.650000 ;
      RECT 466.500000 450.350000 499.500000 451.650000 ;
      RECT 457.500000 450.350000 458.500000 451.650000 ;
      RECT 416.500000 450.350000 449.500000 451.650000 ;
      RECT 407.500000 450.350000 408.500000 451.650000 ;
      RECT 366.500000 450.350000 399.500000 451.650000 ;
      RECT 357.500000 450.350000 358.500000 451.650000 ;
      RECT 316.500000 450.350000 349.500000 451.650000 ;
      RECT 307.500000 450.350000 308.500000 451.650000 ;
      RECT 216.500000 450.350000 299.500000 451.650000 ;
      RECT 207.500000 450.350000 208.500000 451.650000 ;
      RECT 116.500000 450.350000 199.500000 451.650000 ;
      RECT 107.500000 450.350000 108.500000 451.650000 ;
      RECT 66.500000 450.350000 99.500000 451.650000 ;
      RECT 57.500000 450.350000 58.500000 451.650000 ;
      RECT 29.500000 450.350000 49.500000 451.650000 ;
      RECT 15.500000 450.350000 16.500000 451.650000 ;
      RECT 1157.500000 449.650000 1186.000000 450.350000 ;
      RECT 707.500000 449.650000 723.500000 450.350000 ;
      RECT 657.500000 449.650000 699.500000 450.350000 ;
      RECT 607.500000 449.650000 649.500000 450.350000 ;
      RECT 557.500000 449.650000 599.500000 450.350000 ;
      RECT 507.500000 449.650000 549.500000 450.350000 ;
      RECT 457.500000 449.650000 499.500000 450.350000 ;
      RECT 407.500000 449.650000 449.500000 450.350000 ;
      RECT 357.500000 449.650000 399.500000 450.350000 ;
      RECT 307.500000 449.650000 349.500000 450.350000 ;
      RECT 207.500000 449.650000 299.500000 450.350000 ;
      RECT 107.500000 449.650000 199.500000 450.350000 ;
      RECT 57.500000 449.650000 99.500000 450.350000 ;
      RECT 15.500000 449.650000 49.500000 450.350000 ;
      RECT 1157.500000 448.350000 1158.500000 449.650000 ;
      RECT 1139.000000 448.350000 1149.500000 451.650000 ;
      RECT 736.500000 448.350000 739.000000 451.650000 ;
      RECT 722.500000 448.350000 723.500000 449.650000 ;
      RECT 707.500000 448.350000 708.500000 449.650000 ;
      RECT 666.500000 448.350000 699.500000 449.650000 ;
      RECT 657.500000 448.350000 658.500000 449.650000 ;
      RECT 616.500000 448.350000 649.500000 449.650000 ;
      RECT 607.500000 448.350000 608.500000 449.650000 ;
      RECT 566.500000 448.350000 599.500000 449.650000 ;
      RECT 557.500000 448.350000 558.500000 449.650000 ;
      RECT 516.500000 448.350000 549.500000 449.650000 ;
      RECT 507.500000 448.350000 508.500000 449.650000 ;
      RECT 466.500000 448.350000 499.500000 449.650000 ;
      RECT 457.500000 448.350000 458.500000 449.650000 ;
      RECT 416.500000 448.350000 449.500000 449.650000 ;
      RECT 407.500000 448.350000 408.500000 449.650000 ;
      RECT 366.500000 448.350000 399.500000 449.650000 ;
      RECT 357.500000 448.350000 358.500000 449.650000 ;
      RECT 316.500000 448.350000 349.500000 449.650000 ;
      RECT 307.500000 448.350000 308.500000 449.650000 ;
      RECT 216.500000 448.350000 299.500000 449.650000 ;
      RECT 207.500000 448.350000 208.500000 449.650000 ;
      RECT 116.500000 448.350000 199.500000 449.650000 ;
      RECT 107.500000 448.350000 108.500000 449.650000 ;
      RECT 66.500000 448.350000 99.500000 449.650000 ;
      RECT 57.500000 448.350000 58.500000 449.650000 ;
      RECT 29.500000 448.350000 49.500000 449.650000 ;
      RECT 15.500000 448.350000 16.500000 449.650000 ;
      RECT 0.000000 448.350000 2.500000 451.650000 ;
      RECT 1139.000000 447.650000 1158.500000 448.350000 ;
      RECT 722.500000 447.650000 739.000000 448.350000 ;
      RECT 666.500000 447.650000 708.500000 448.350000 ;
      RECT 616.500000 447.650000 658.500000 448.350000 ;
      RECT 566.500000 447.650000 608.500000 448.350000 ;
      RECT 516.500000 447.650000 558.500000 448.350000 ;
      RECT 466.500000 447.650000 508.500000 448.350000 ;
      RECT 416.500000 447.650000 458.500000 448.350000 ;
      RECT 366.500000 447.650000 408.500000 448.350000 ;
      RECT 316.500000 447.650000 358.500000 448.350000 ;
      RECT 216.500000 447.650000 308.500000 448.350000 ;
      RECT 116.500000 447.650000 208.500000 448.350000 ;
      RECT 66.500000 447.650000 108.500000 448.350000 ;
      RECT 29.500000 447.650000 58.500000 448.350000 ;
      RECT 0.000000 447.650000 16.500000 448.350000 ;
      RECT 1166.500000 446.350000 1186.000000 449.650000 ;
      RECT 1157.500000 446.350000 1158.500000 447.650000 ;
      RECT 722.500000 446.350000 723.500000 447.650000 ;
      RECT 707.500000 446.350000 708.500000 447.650000 ;
      RECT 666.500000 446.350000 699.500000 447.650000 ;
      RECT 657.500000 446.350000 658.500000 447.650000 ;
      RECT 616.500000 446.350000 649.500000 447.650000 ;
      RECT 607.500000 446.350000 608.500000 447.650000 ;
      RECT 566.500000 446.350000 599.500000 447.650000 ;
      RECT 557.500000 446.350000 558.500000 447.650000 ;
      RECT 516.500000 446.350000 549.500000 447.650000 ;
      RECT 507.500000 446.350000 508.500000 447.650000 ;
      RECT 466.500000 446.350000 499.500000 447.650000 ;
      RECT 457.500000 446.350000 458.500000 447.650000 ;
      RECT 416.500000 446.350000 449.500000 447.650000 ;
      RECT 407.500000 446.350000 408.500000 447.650000 ;
      RECT 366.500000 446.350000 399.500000 447.650000 ;
      RECT 357.500000 446.350000 358.500000 447.650000 ;
      RECT 316.500000 446.350000 349.500000 447.650000 ;
      RECT 307.500000 446.350000 308.500000 447.650000 ;
      RECT 216.500000 446.350000 299.500000 447.650000 ;
      RECT 207.500000 446.350000 208.500000 447.650000 ;
      RECT 116.500000 446.350000 199.500000 447.650000 ;
      RECT 107.500000 446.350000 108.500000 447.650000 ;
      RECT 66.500000 446.350000 99.500000 447.650000 ;
      RECT 57.500000 446.350000 58.500000 447.650000 ;
      RECT 29.500000 446.350000 49.500000 447.650000 ;
      RECT 15.500000 446.350000 16.500000 447.650000 ;
      RECT 1139.000000 446.000000 1149.500000 447.650000 ;
      RECT 736.500000 446.000000 739.000000 447.650000 ;
      RECT 1157.500000 445.650000 1186.000000 446.350000 ;
      RECT 736.500000 445.650000 1149.500000 446.000000 ;
      RECT 707.500000 445.650000 723.500000 446.350000 ;
      RECT 657.500000 445.650000 699.500000 446.350000 ;
      RECT 607.500000 445.650000 649.500000 446.350000 ;
      RECT 557.500000 445.650000 599.500000 446.350000 ;
      RECT 507.500000 445.650000 549.500000 446.350000 ;
      RECT 457.500000 445.650000 499.500000 446.350000 ;
      RECT 407.500000 445.650000 449.500000 446.350000 ;
      RECT 357.500000 445.650000 399.500000 446.350000 ;
      RECT 307.500000 445.650000 349.500000 446.350000 ;
      RECT 207.500000 445.650000 299.500000 446.350000 ;
      RECT 107.500000 445.650000 199.500000 446.350000 ;
      RECT 57.500000 445.650000 99.500000 446.350000 ;
      RECT 15.500000 445.650000 49.500000 446.350000 ;
      RECT 1157.500000 444.350000 1158.500000 445.650000 ;
      RECT 1116.500000 444.350000 1149.500000 445.650000 ;
      RECT 736.500000 444.350000 758.500000 445.650000 ;
      RECT 722.500000 444.350000 723.500000 445.650000 ;
      RECT 707.500000 444.350000 708.500000 445.650000 ;
      RECT 666.500000 444.350000 699.500000 445.650000 ;
      RECT 657.500000 444.350000 658.500000 445.650000 ;
      RECT 616.500000 444.350000 649.500000 445.650000 ;
      RECT 607.500000 444.350000 608.500000 445.650000 ;
      RECT 566.500000 444.350000 599.500000 445.650000 ;
      RECT 557.500000 444.350000 558.500000 445.650000 ;
      RECT 516.500000 444.350000 549.500000 445.650000 ;
      RECT 507.500000 444.350000 508.500000 445.650000 ;
      RECT 466.500000 444.350000 499.500000 445.650000 ;
      RECT 457.500000 444.350000 458.500000 445.650000 ;
      RECT 416.500000 444.350000 449.500000 445.650000 ;
      RECT 407.500000 444.350000 408.500000 445.650000 ;
      RECT 366.500000 444.350000 399.500000 445.650000 ;
      RECT 357.500000 444.350000 358.500000 445.650000 ;
      RECT 316.500000 444.350000 349.500000 445.650000 ;
      RECT 307.500000 444.350000 308.500000 445.650000 ;
      RECT 216.500000 444.350000 299.500000 445.650000 ;
      RECT 207.500000 444.350000 208.500000 445.650000 ;
      RECT 116.500000 444.350000 199.500000 445.650000 ;
      RECT 107.500000 444.350000 108.500000 445.650000 ;
      RECT 66.500000 444.350000 99.500000 445.650000 ;
      RECT 57.500000 444.350000 58.500000 445.650000 ;
      RECT 29.500000 444.350000 49.500000 445.650000 ;
      RECT 15.500000 444.350000 16.500000 445.650000 ;
      RECT 0.000000 444.350000 2.500000 447.650000 ;
      RECT 1166.500000 443.650000 1186.000000 445.650000 ;
      RECT 1116.500000 443.650000 1158.500000 444.350000 ;
      RECT 1066.500000 443.650000 1108.500000 445.650000 ;
      RECT 1016.500000 443.650000 1058.500000 445.650000 ;
      RECT 966.500000 443.650000 1008.500000 445.650000 ;
      RECT 916.500000 443.650000 958.500000 445.650000 ;
      RECT 866.500000 443.650000 908.500000 445.650000 ;
      RECT 816.500000 443.650000 858.500000 445.650000 ;
      RECT 766.500000 443.650000 808.500000 445.650000 ;
      RECT 722.500000 443.650000 758.500000 444.350000 ;
      RECT 666.500000 443.650000 708.500000 444.350000 ;
      RECT 616.500000 443.650000 658.500000 444.350000 ;
      RECT 566.500000 443.650000 608.500000 444.350000 ;
      RECT 516.500000 443.650000 558.500000 444.350000 ;
      RECT 466.500000 443.650000 508.500000 444.350000 ;
      RECT 416.500000 443.650000 458.500000 444.350000 ;
      RECT 366.500000 443.650000 408.500000 444.350000 ;
      RECT 316.500000 443.650000 358.500000 444.350000 ;
      RECT 216.500000 443.650000 308.500000 444.350000 ;
      RECT 116.500000 443.650000 208.500000 444.350000 ;
      RECT 66.500000 443.650000 108.500000 444.350000 ;
      RECT 29.500000 443.650000 58.500000 444.350000 ;
      RECT 0.000000 443.650000 16.500000 444.350000 ;
      RECT 1166.500000 442.350000 1170.500000 443.650000 ;
      RECT 1157.500000 442.350000 1158.500000 443.650000 ;
      RECT 1116.500000 442.350000 1149.500000 443.650000 ;
      RECT 1107.500000 442.350000 1108.500000 443.650000 ;
      RECT 1066.500000 442.350000 1099.500000 443.650000 ;
      RECT 1057.500000 442.350000 1058.500000 443.650000 ;
      RECT 1016.500000 442.350000 1049.500000 443.650000 ;
      RECT 1007.500000 442.350000 1008.500000 443.650000 ;
      RECT 966.500000 442.350000 999.500000 443.650000 ;
      RECT 957.500000 442.350000 958.500000 443.650000 ;
      RECT 916.500000 442.350000 949.500000 443.650000 ;
      RECT 907.500000 442.350000 908.500000 443.650000 ;
      RECT 866.500000 442.350000 899.500000 443.650000 ;
      RECT 857.500000 442.350000 858.500000 443.650000 ;
      RECT 816.500000 442.350000 849.500000 443.650000 ;
      RECT 807.500000 442.350000 808.500000 443.650000 ;
      RECT 766.500000 442.350000 799.500000 443.650000 ;
      RECT 757.500000 442.350000 758.500000 443.650000 ;
      RECT 722.500000 442.350000 723.500000 443.650000 ;
      RECT 707.500000 442.350000 708.500000 443.650000 ;
      RECT 666.500000 442.350000 699.500000 443.650000 ;
      RECT 657.500000 442.350000 658.500000 443.650000 ;
      RECT 616.500000 442.350000 649.500000 443.650000 ;
      RECT 607.500000 442.350000 608.500000 443.650000 ;
      RECT 566.500000 442.350000 599.500000 443.650000 ;
      RECT 557.500000 442.350000 558.500000 443.650000 ;
      RECT 516.500000 442.350000 549.500000 443.650000 ;
      RECT 507.500000 442.350000 508.500000 443.650000 ;
      RECT 466.500000 442.350000 499.500000 443.650000 ;
      RECT 457.500000 442.350000 458.500000 443.650000 ;
      RECT 416.500000 442.350000 449.500000 443.650000 ;
      RECT 407.500000 442.350000 408.500000 443.650000 ;
      RECT 366.500000 442.350000 399.500000 443.650000 ;
      RECT 357.500000 442.350000 358.500000 443.650000 ;
      RECT 316.500000 442.350000 349.500000 443.650000 ;
      RECT 307.500000 442.350000 308.500000 443.650000 ;
      RECT 216.500000 442.350000 299.500000 443.650000 ;
      RECT 207.500000 442.350000 208.500000 443.650000 ;
      RECT 116.500000 442.350000 199.500000 443.650000 ;
      RECT 107.500000 442.350000 108.500000 443.650000 ;
      RECT 66.500000 442.350000 99.500000 443.650000 ;
      RECT 57.500000 442.350000 58.500000 443.650000 ;
      RECT 29.500000 442.350000 49.500000 443.650000 ;
      RECT 15.500000 442.350000 16.500000 443.650000 ;
      RECT 1157.500000 441.650000 1170.500000 442.350000 ;
      RECT 1107.500000 441.650000 1149.500000 442.350000 ;
      RECT 1057.500000 441.650000 1099.500000 442.350000 ;
      RECT 1007.500000 441.650000 1049.500000 442.350000 ;
      RECT 957.500000 441.650000 999.500000 442.350000 ;
      RECT 907.500000 441.650000 949.500000 442.350000 ;
      RECT 857.500000 441.650000 899.500000 442.350000 ;
      RECT 807.500000 441.650000 849.500000 442.350000 ;
      RECT 757.500000 441.650000 799.500000 442.350000 ;
      RECT 707.500000 441.650000 723.500000 442.350000 ;
      RECT 657.500000 441.650000 699.500000 442.350000 ;
      RECT 607.500000 441.650000 649.500000 442.350000 ;
      RECT 557.500000 441.650000 599.500000 442.350000 ;
      RECT 507.500000 441.650000 549.500000 442.350000 ;
      RECT 457.500000 441.650000 499.500000 442.350000 ;
      RECT 407.500000 441.650000 449.500000 442.350000 ;
      RECT 357.500000 441.650000 399.500000 442.350000 ;
      RECT 307.500000 441.650000 349.500000 442.350000 ;
      RECT 207.500000 441.650000 299.500000 442.350000 ;
      RECT 107.500000 441.650000 199.500000 442.350000 ;
      RECT 57.500000 441.650000 99.500000 442.350000 ;
      RECT 15.500000 441.650000 49.500000 442.350000 ;
      RECT 1183.500000 440.350000 1186.000000 443.650000 ;
      RECT 1166.500000 440.350000 1170.500000 441.650000 ;
      RECT 1157.500000 440.350000 1158.500000 441.650000 ;
      RECT 1116.500000 440.350000 1149.500000 441.650000 ;
      RECT 1107.500000 440.350000 1108.500000 441.650000 ;
      RECT 1066.500000 440.350000 1099.500000 441.650000 ;
      RECT 1057.500000 440.350000 1058.500000 441.650000 ;
      RECT 1016.500000 440.350000 1049.500000 441.650000 ;
      RECT 1007.500000 440.350000 1008.500000 441.650000 ;
      RECT 966.500000 440.350000 999.500000 441.650000 ;
      RECT 957.500000 440.350000 958.500000 441.650000 ;
      RECT 916.500000 440.350000 949.500000 441.650000 ;
      RECT 907.500000 440.350000 908.500000 441.650000 ;
      RECT 866.500000 440.350000 899.500000 441.650000 ;
      RECT 857.500000 440.350000 858.500000 441.650000 ;
      RECT 816.500000 440.350000 849.500000 441.650000 ;
      RECT 807.500000 440.350000 808.500000 441.650000 ;
      RECT 766.500000 440.350000 799.500000 441.650000 ;
      RECT 757.500000 440.350000 758.500000 441.650000 ;
      RECT 736.500000 440.350000 749.500000 443.650000 ;
      RECT 722.500000 440.350000 723.500000 441.650000 ;
      RECT 707.500000 440.350000 708.500000 441.650000 ;
      RECT 666.500000 440.350000 699.500000 441.650000 ;
      RECT 657.500000 440.350000 658.500000 441.650000 ;
      RECT 616.500000 440.350000 649.500000 441.650000 ;
      RECT 607.500000 440.350000 608.500000 441.650000 ;
      RECT 566.500000 440.350000 599.500000 441.650000 ;
      RECT 557.500000 440.350000 558.500000 441.650000 ;
      RECT 516.500000 440.350000 549.500000 441.650000 ;
      RECT 507.500000 440.350000 508.500000 441.650000 ;
      RECT 466.500000 440.350000 499.500000 441.650000 ;
      RECT 457.500000 440.350000 458.500000 441.650000 ;
      RECT 416.500000 440.350000 449.500000 441.650000 ;
      RECT 407.500000 440.350000 408.500000 441.650000 ;
      RECT 366.500000 440.350000 399.500000 441.650000 ;
      RECT 357.500000 440.350000 358.500000 441.650000 ;
      RECT 316.500000 440.350000 349.500000 441.650000 ;
      RECT 307.500000 440.350000 308.500000 441.650000 ;
      RECT 216.500000 440.350000 299.500000 441.650000 ;
      RECT 207.500000 440.350000 208.500000 441.650000 ;
      RECT 116.500000 440.350000 199.500000 441.650000 ;
      RECT 107.500000 440.350000 108.500000 441.650000 ;
      RECT 66.500000 440.350000 99.500000 441.650000 ;
      RECT 57.500000 440.350000 58.500000 441.650000 ;
      RECT 29.500000 440.350000 49.500000 441.650000 ;
      RECT 15.500000 440.350000 16.500000 441.650000 ;
      RECT 0.000000 440.350000 2.500000 443.650000 ;
      RECT 1166.500000 439.650000 1186.000000 440.350000 ;
      RECT 1116.500000 439.650000 1158.500000 440.350000 ;
      RECT 1066.500000 439.650000 1108.500000 440.350000 ;
      RECT 1016.500000 439.650000 1058.500000 440.350000 ;
      RECT 966.500000 439.650000 1008.500000 440.350000 ;
      RECT 916.500000 439.650000 958.500000 440.350000 ;
      RECT 866.500000 439.650000 908.500000 440.350000 ;
      RECT 816.500000 439.650000 858.500000 440.350000 ;
      RECT 766.500000 439.650000 808.500000 440.350000 ;
      RECT 722.500000 439.650000 758.500000 440.350000 ;
      RECT 666.500000 439.650000 708.500000 440.350000 ;
      RECT 616.500000 439.650000 658.500000 440.350000 ;
      RECT 566.500000 439.650000 608.500000 440.350000 ;
      RECT 516.500000 439.650000 558.500000 440.350000 ;
      RECT 466.500000 439.650000 508.500000 440.350000 ;
      RECT 416.500000 439.650000 458.500000 440.350000 ;
      RECT 366.500000 439.650000 408.500000 440.350000 ;
      RECT 316.500000 439.650000 358.500000 440.350000 ;
      RECT 216.500000 439.650000 308.500000 440.350000 ;
      RECT 116.500000 439.650000 208.500000 440.350000 ;
      RECT 66.500000 439.650000 108.500000 440.350000 ;
      RECT 29.500000 439.650000 58.500000 440.350000 ;
      RECT 0.000000 439.650000 16.500000 440.350000 ;
      RECT 1166.500000 438.350000 1170.500000 439.650000 ;
      RECT 1157.500000 438.350000 1158.500000 439.650000 ;
      RECT 1116.500000 438.350000 1149.500000 439.650000 ;
      RECT 1107.500000 438.350000 1108.500000 439.650000 ;
      RECT 1066.500000 438.350000 1099.500000 439.650000 ;
      RECT 1057.500000 438.350000 1058.500000 439.650000 ;
      RECT 1016.500000 438.350000 1049.500000 439.650000 ;
      RECT 1007.500000 438.350000 1008.500000 439.650000 ;
      RECT 966.500000 438.350000 999.500000 439.650000 ;
      RECT 957.500000 438.350000 958.500000 439.650000 ;
      RECT 916.500000 438.350000 949.500000 439.650000 ;
      RECT 907.500000 438.350000 908.500000 439.650000 ;
      RECT 866.500000 438.350000 899.500000 439.650000 ;
      RECT 857.500000 438.350000 858.500000 439.650000 ;
      RECT 816.500000 438.350000 849.500000 439.650000 ;
      RECT 807.500000 438.350000 808.500000 439.650000 ;
      RECT 766.500000 438.350000 799.500000 439.650000 ;
      RECT 757.500000 438.350000 758.500000 439.650000 ;
      RECT 722.500000 438.350000 723.500000 439.650000 ;
      RECT 707.500000 438.350000 708.500000 439.650000 ;
      RECT 666.500000 438.350000 699.500000 439.650000 ;
      RECT 657.500000 438.350000 658.500000 439.650000 ;
      RECT 616.500000 438.350000 649.500000 439.650000 ;
      RECT 607.500000 438.350000 608.500000 439.650000 ;
      RECT 566.500000 438.350000 599.500000 439.650000 ;
      RECT 557.500000 438.350000 558.500000 439.650000 ;
      RECT 516.500000 438.350000 549.500000 439.650000 ;
      RECT 507.500000 438.350000 508.500000 439.650000 ;
      RECT 466.500000 438.350000 499.500000 439.650000 ;
      RECT 457.500000 438.350000 458.500000 439.650000 ;
      RECT 416.500000 438.350000 449.500000 439.650000 ;
      RECT 407.500000 438.350000 408.500000 439.650000 ;
      RECT 366.500000 438.350000 399.500000 439.650000 ;
      RECT 357.500000 438.350000 358.500000 439.650000 ;
      RECT 316.500000 438.350000 349.500000 439.650000 ;
      RECT 307.500000 438.350000 308.500000 439.650000 ;
      RECT 216.500000 438.350000 299.500000 439.650000 ;
      RECT 207.500000 438.350000 208.500000 439.650000 ;
      RECT 116.500000 438.350000 199.500000 439.650000 ;
      RECT 107.500000 438.350000 108.500000 439.650000 ;
      RECT 66.500000 438.350000 99.500000 439.650000 ;
      RECT 57.500000 438.350000 58.500000 439.650000 ;
      RECT 29.500000 438.350000 49.500000 439.650000 ;
      RECT 15.500000 438.350000 16.500000 439.650000 ;
      RECT 1157.500000 437.650000 1170.500000 438.350000 ;
      RECT 1107.500000 437.650000 1149.500000 438.350000 ;
      RECT 1057.500000 437.650000 1099.500000 438.350000 ;
      RECT 1007.500000 437.650000 1049.500000 438.350000 ;
      RECT 957.500000 437.650000 999.500000 438.350000 ;
      RECT 907.500000 437.650000 949.500000 438.350000 ;
      RECT 857.500000 437.650000 899.500000 438.350000 ;
      RECT 807.500000 437.650000 849.500000 438.350000 ;
      RECT 757.500000 437.650000 799.500000 438.350000 ;
      RECT 707.500000 437.650000 723.500000 438.350000 ;
      RECT 657.500000 437.650000 699.500000 438.350000 ;
      RECT 607.500000 437.650000 649.500000 438.350000 ;
      RECT 557.500000 437.650000 599.500000 438.350000 ;
      RECT 507.500000 437.650000 549.500000 438.350000 ;
      RECT 457.500000 437.650000 499.500000 438.350000 ;
      RECT 407.500000 437.650000 449.500000 438.350000 ;
      RECT 357.500000 437.650000 399.500000 438.350000 ;
      RECT 307.500000 437.650000 349.500000 438.350000 ;
      RECT 207.500000 437.650000 299.500000 438.350000 ;
      RECT 107.500000 437.650000 199.500000 438.350000 ;
      RECT 57.500000 437.650000 99.500000 438.350000 ;
      RECT 15.500000 437.650000 49.500000 438.350000 ;
      RECT 1183.500000 436.350000 1186.000000 439.650000 ;
      RECT 1166.500000 436.350000 1170.500000 437.650000 ;
      RECT 1157.500000 436.350000 1158.500000 437.650000 ;
      RECT 1116.500000 436.350000 1149.500000 437.650000 ;
      RECT 1107.500000 436.350000 1108.500000 437.650000 ;
      RECT 1066.500000 436.350000 1099.500000 437.650000 ;
      RECT 1057.500000 436.350000 1058.500000 437.650000 ;
      RECT 1016.500000 436.350000 1049.500000 437.650000 ;
      RECT 1007.500000 436.350000 1008.500000 437.650000 ;
      RECT 966.500000 436.350000 999.500000 437.650000 ;
      RECT 957.500000 436.350000 958.500000 437.650000 ;
      RECT 916.500000 436.350000 949.500000 437.650000 ;
      RECT 907.500000 436.350000 908.500000 437.650000 ;
      RECT 866.500000 436.350000 899.500000 437.650000 ;
      RECT 857.500000 436.350000 858.500000 437.650000 ;
      RECT 816.500000 436.350000 849.500000 437.650000 ;
      RECT 807.500000 436.350000 808.500000 437.650000 ;
      RECT 766.500000 436.350000 799.500000 437.650000 ;
      RECT 757.500000 436.350000 758.500000 437.650000 ;
      RECT 736.500000 436.350000 749.500000 439.650000 ;
      RECT 722.500000 436.350000 723.500000 437.650000 ;
      RECT 707.500000 436.350000 708.500000 437.650000 ;
      RECT 666.500000 436.350000 699.500000 437.650000 ;
      RECT 657.500000 436.350000 658.500000 437.650000 ;
      RECT 616.500000 436.350000 649.500000 437.650000 ;
      RECT 607.500000 436.350000 608.500000 437.650000 ;
      RECT 566.500000 436.350000 599.500000 437.650000 ;
      RECT 557.500000 436.350000 558.500000 437.650000 ;
      RECT 516.500000 436.350000 549.500000 437.650000 ;
      RECT 507.500000 436.350000 508.500000 437.650000 ;
      RECT 466.500000 436.350000 499.500000 437.650000 ;
      RECT 457.500000 436.350000 458.500000 437.650000 ;
      RECT 416.500000 436.350000 449.500000 437.650000 ;
      RECT 407.500000 436.350000 408.500000 437.650000 ;
      RECT 366.500000 436.350000 399.500000 437.650000 ;
      RECT 357.500000 436.350000 358.500000 437.650000 ;
      RECT 316.500000 436.350000 349.500000 437.650000 ;
      RECT 307.500000 436.350000 308.500000 437.650000 ;
      RECT 216.500000 436.350000 299.500000 437.650000 ;
      RECT 207.500000 436.350000 208.500000 437.650000 ;
      RECT 116.500000 436.350000 199.500000 437.650000 ;
      RECT 107.500000 436.350000 108.500000 437.650000 ;
      RECT 66.500000 436.350000 99.500000 437.650000 ;
      RECT 57.500000 436.350000 58.500000 437.650000 ;
      RECT 29.500000 436.350000 49.500000 437.650000 ;
      RECT 15.500000 436.350000 16.500000 437.650000 ;
      RECT 0.000000 436.350000 2.500000 439.650000 ;
      RECT 1166.500000 435.650000 1186.000000 436.350000 ;
      RECT 1116.500000 435.650000 1158.500000 436.350000 ;
      RECT 1066.500000 435.650000 1108.500000 436.350000 ;
      RECT 1016.500000 435.650000 1058.500000 436.350000 ;
      RECT 966.500000 435.650000 1008.500000 436.350000 ;
      RECT 916.500000 435.650000 958.500000 436.350000 ;
      RECT 866.500000 435.650000 908.500000 436.350000 ;
      RECT 816.500000 435.650000 858.500000 436.350000 ;
      RECT 766.500000 435.650000 808.500000 436.350000 ;
      RECT 722.500000 435.650000 758.500000 436.350000 ;
      RECT 666.500000 435.650000 708.500000 436.350000 ;
      RECT 616.500000 435.650000 658.500000 436.350000 ;
      RECT 566.500000 435.650000 608.500000 436.350000 ;
      RECT 516.500000 435.650000 558.500000 436.350000 ;
      RECT 466.500000 435.650000 508.500000 436.350000 ;
      RECT 416.500000 435.650000 458.500000 436.350000 ;
      RECT 366.500000 435.650000 408.500000 436.350000 ;
      RECT 316.500000 435.650000 358.500000 436.350000 ;
      RECT 216.500000 435.650000 308.500000 436.350000 ;
      RECT 116.500000 435.650000 208.500000 436.350000 ;
      RECT 66.500000 435.650000 108.500000 436.350000 ;
      RECT 29.500000 435.650000 58.500000 436.350000 ;
      RECT 0.000000 435.650000 16.500000 436.350000 ;
      RECT 1166.500000 434.350000 1170.500000 435.650000 ;
      RECT 1157.500000 434.350000 1158.500000 435.650000 ;
      RECT 1116.500000 434.350000 1149.500000 435.650000 ;
      RECT 1107.500000 434.350000 1108.500000 435.650000 ;
      RECT 1066.500000 434.350000 1099.500000 435.650000 ;
      RECT 1057.500000 434.350000 1058.500000 435.650000 ;
      RECT 1016.500000 434.350000 1049.500000 435.650000 ;
      RECT 1007.500000 434.350000 1008.500000 435.650000 ;
      RECT 966.500000 434.350000 999.500000 435.650000 ;
      RECT 957.500000 434.350000 958.500000 435.650000 ;
      RECT 916.500000 434.350000 949.500000 435.650000 ;
      RECT 907.500000 434.350000 908.500000 435.650000 ;
      RECT 866.500000 434.350000 899.500000 435.650000 ;
      RECT 857.500000 434.350000 858.500000 435.650000 ;
      RECT 816.500000 434.350000 849.500000 435.650000 ;
      RECT 807.500000 434.350000 808.500000 435.650000 ;
      RECT 766.500000 434.350000 799.500000 435.650000 ;
      RECT 757.500000 434.350000 758.500000 435.650000 ;
      RECT 722.500000 434.350000 723.500000 435.650000 ;
      RECT 707.500000 434.350000 708.500000 435.650000 ;
      RECT 666.500000 434.350000 699.500000 435.650000 ;
      RECT 657.500000 434.350000 658.500000 435.650000 ;
      RECT 616.500000 434.350000 649.500000 435.650000 ;
      RECT 607.500000 434.350000 608.500000 435.650000 ;
      RECT 566.500000 434.350000 599.500000 435.650000 ;
      RECT 557.500000 434.350000 558.500000 435.650000 ;
      RECT 516.500000 434.350000 549.500000 435.650000 ;
      RECT 507.500000 434.350000 508.500000 435.650000 ;
      RECT 466.500000 434.350000 499.500000 435.650000 ;
      RECT 457.500000 434.350000 458.500000 435.650000 ;
      RECT 416.500000 434.350000 449.500000 435.650000 ;
      RECT 407.500000 434.350000 408.500000 435.650000 ;
      RECT 366.500000 434.350000 399.500000 435.650000 ;
      RECT 357.500000 434.350000 358.500000 435.650000 ;
      RECT 316.500000 434.350000 349.500000 435.650000 ;
      RECT 307.500000 434.350000 308.500000 435.650000 ;
      RECT 216.500000 434.350000 299.500000 435.650000 ;
      RECT 207.500000 434.350000 208.500000 435.650000 ;
      RECT 116.500000 434.350000 199.500000 435.650000 ;
      RECT 107.500000 434.350000 108.500000 435.650000 ;
      RECT 66.500000 434.350000 99.500000 435.650000 ;
      RECT 57.500000 434.350000 58.500000 435.650000 ;
      RECT 29.500000 434.350000 49.500000 435.650000 ;
      RECT 15.500000 434.350000 16.500000 435.650000 ;
      RECT 1157.500000 433.650000 1170.500000 434.350000 ;
      RECT 1107.500000 433.650000 1149.500000 434.350000 ;
      RECT 1057.500000 433.650000 1099.500000 434.350000 ;
      RECT 1007.500000 433.650000 1049.500000 434.350000 ;
      RECT 957.500000 433.650000 999.500000 434.350000 ;
      RECT 907.500000 433.650000 949.500000 434.350000 ;
      RECT 857.500000 433.650000 899.500000 434.350000 ;
      RECT 807.500000 433.650000 849.500000 434.350000 ;
      RECT 757.500000 433.650000 799.500000 434.350000 ;
      RECT 707.500000 433.650000 723.500000 434.350000 ;
      RECT 657.500000 433.650000 699.500000 434.350000 ;
      RECT 607.500000 433.650000 649.500000 434.350000 ;
      RECT 557.500000 433.650000 599.500000 434.350000 ;
      RECT 507.500000 433.650000 549.500000 434.350000 ;
      RECT 457.500000 433.650000 499.500000 434.350000 ;
      RECT 407.500000 433.650000 449.500000 434.350000 ;
      RECT 357.500000 433.650000 399.500000 434.350000 ;
      RECT 307.500000 433.650000 349.500000 434.350000 ;
      RECT 207.500000 433.650000 299.500000 434.350000 ;
      RECT 107.500000 433.650000 199.500000 434.350000 ;
      RECT 57.500000 433.650000 99.500000 434.350000 ;
      RECT 15.500000 433.650000 49.500000 434.350000 ;
      RECT 1183.500000 432.350000 1186.000000 435.650000 ;
      RECT 1166.500000 432.350000 1170.500000 433.650000 ;
      RECT 1157.500000 432.350000 1158.500000 433.650000 ;
      RECT 1116.500000 432.350000 1149.500000 433.650000 ;
      RECT 1107.500000 432.350000 1108.500000 433.650000 ;
      RECT 1066.500000 432.350000 1099.500000 433.650000 ;
      RECT 1057.500000 432.350000 1058.500000 433.650000 ;
      RECT 1016.500000 432.350000 1049.500000 433.650000 ;
      RECT 1007.500000 432.350000 1008.500000 433.650000 ;
      RECT 966.500000 432.350000 999.500000 433.650000 ;
      RECT 957.500000 432.350000 958.500000 433.650000 ;
      RECT 916.500000 432.350000 949.500000 433.650000 ;
      RECT 907.500000 432.350000 908.500000 433.650000 ;
      RECT 866.500000 432.350000 899.500000 433.650000 ;
      RECT 857.500000 432.350000 858.500000 433.650000 ;
      RECT 816.500000 432.350000 849.500000 433.650000 ;
      RECT 807.500000 432.350000 808.500000 433.650000 ;
      RECT 766.500000 432.350000 799.500000 433.650000 ;
      RECT 757.500000 432.350000 758.500000 433.650000 ;
      RECT 736.500000 432.350000 749.500000 435.650000 ;
      RECT 722.500000 432.350000 723.500000 433.650000 ;
      RECT 707.500000 432.350000 708.500000 433.650000 ;
      RECT 666.500000 432.350000 699.500000 433.650000 ;
      RECT 657.500000 432.350000 658.500000 433.650000 ;
      RECT 616.500000 432.350000 649.500000 433.650000 ;
      RECT 607.500000 432.350000 608.500000 433.650000 ;
      RECT 566.500000 432.350000 599.500000 433.650000 ;
      RECT 557.500000 432.350000 558.500000 433.650000 ;
      RECT 516.500000 432.350000 549.500000 433.650000 ;
      RECT 507.500000 432.350000 508.500000 433.650000 ;
      RECT 466.500000 432.350000 499.500000 433.650000 ;
      RECT 457.500000 432.350000 458.500000 433.650000 ;
      RECT 416.500000 432.350000 449.500000 433.650000 ;
      RECT 407.500000 432.350000 408.500000 433.650000 ;
      RECT 366.500000 432.350000 399.500000 433.650000 ;
      RECT 357.500000 432.350000 358.500000 433.650000 ;
      RECT 316.500000 432.350000 349.500000 433.650000 ;
      RECT 307.500000 432.350000 308.500000 433.650000 ;
      RECT 216.500000 432.350000 299.500000 433.650000 ;
      RECT 207.500000 432.350000 208.500000 433.650000 ;
      RECT 116.500000 432.350000 199.500000 433.650000 ;
      RECT 107.500000 432.350000 108.500000 433.650000 ;
      RECT 66.500000 432.350000 99.500000 433.650000 ;
      RECT 57.500000 432.350000 58.500000 433.650000 ;
      RECT 29.500000 432.350000 49.500000 433.650000 ;
      RECT 15.500000 432.350000 16.500000 433.650000 ;
      RECT 0.000000 432.350000 2.500000 435.650000 ;
      RECT 1166.500000 431.650000 1186.000000 432.350000 ;
      RECT 1116.500000 431.650000 1158.500000 432.350000 ;
      RECT 1066.500000 431.650000 1108.500000 432.350000 ;
      RECT 1016.500000 431.650000 1058.500000 432.350000 ;
      RECT 966.500000 431.650000 1008.500000 432.350000 ;
      RECT 916.500000 431.650000 958.500000 432.350000 ;
      RECT 866.500000 431.650000 908.500000 432.350000 ;
      RECT 816.500000 431.650000 858.500000 432.350000 ;
      RECT 766.500000 431.650000 808.500000 432.350000 ;
      RECT 722.500000 431.650000 758.500000 432.350000 ;
      RECT 666.500000 431.650000 708.500000 432.350000 ;
      RECT 616.500000 431.650000 658.500000 432.350000 ;
      RECT 566.500000 431.650000 608.500000 432.350000 ;
      RECT 516.500000 431.650000 558.500000 432.350000 ;
      RECT 466.500000 431.650000 508.500000 432.350000 ;
      RECT 416.500000 431.650000 458.500000 432.350000 ;
      RECT 366.500000 431.650000 408.500000 432.350000 ;
      RECT 316.500000 431.650000 358.500000 432.350000 ;
      RECT 216.500000 431.650000 308.500000 432.350000 ;
      RECT 116.500000 431.650000 208.500000 432.350000 ;
      RECT 66.500000 431.650000 108.500000 432.350000 ;
      RECT 29.500000 431.650000 58.500000 432.350000 ;
      RECT 0.000000 431.650000 16.500000 432.350000 ;
      RECT 1166.500000 430.350000 1170.500000 431.650000 ;
      RECT 1157.500000 430.350000 1158.500000 431.650000 ;
      RECT 1116.500000 430.350000 1149.500000 431.650000 ;
      RECT 1107.500000 430.350000 1108.500000 431.650000 ;
      RECT 1066.500000 430.350000 1099.500000 431.650000 ;
      RECT 1057.500000 430.350000 1058.500000 431.650000 ;
      RECT 1016.500000 430.350000 1049.500000 431.650000 ;
      RECT 1007.500000 430.350000 1008.500000 431.650000 ;
      RECT 966.500000 430.350000 999.500000 431.650000 ;
      RECT 957.500000 430.350000 958.500000 431.650000 ;
      RECT 916.500000 430.350000 949.500000 431.650000 ;
      RECT 907.500000 430.350000 908.500000 431.650000 ;
      RECT 866.500000 430.350000 899.500000 431.650000 ;
      RECT 857.500000 430.350000 858.500000 431.650000 ;
      RECT 816.500000 430.350000 849.500000 431.650000 ;
      RECT 807.500000 430.350000 808.500000 431.650000 ;
      RECT 766.500000 430.350000 799.500000 431.650000 ;
      RECT 757.500000 430.350000 758.500000 431.650000 ;
      RECT 722.500000 430.350000 749.500000 431.650000 ;
      RECT 707.500000 430.350000 708.500000 431.650000 ;
      RECT 666.500000 430.350000 699.500000 431.650000 ;
      RECT 657.500000 430.350000 658.500000 431.650000 ;
      RECT 616.500000 430.350000 649.500000 431.650000 ;
      RECT 607.500000 430.350000 608.500000 431.650000 ;
      RECT 566.500000 430.350000 599.500000 431.650000 ;
      RECT 557.500000 430.350000 558.500000 431.650000 ;
      RECT 516.500000 430.350000 549.500000 431.650000 ;
      RECT 507.500000 430.350000 508.500000 431.650000 ;
      RECT 466.500000 430.350000 499.500000 431.650000 ;
      RECT 457.500000 430.350000 458.500000 431.650000 ;
      RECT 416.500000 430.350000 449.500000 431.650000 ;
      RECT 407.500000 430.350000 408.500000 431.650000 ;
      RECT 366.500000 430.350000 399.500000 431.650000 ;
      RECT 357.500000 430.350000 358.500000 431.650000 ;
      RECT 316.500000 430.350000 349.500000 431.650000 ;
      RECT 307.500000 430.350000 308.500000 431.650000 ;
      RECT 216.500000 430.350000 299.500000 431.650000 ;
      RECT 207.500000 430.350000 208.500000 431.650000 ;
      RECT 116.500000 430.350000 199.500000 431.650000 ;
      RECT 107.500000 430.350000 108.500000 431.650000 ;
      RECT 66.500000 430.350000 99.500000 431.650000 ;
      RECT 57.500000 430.350000 58.500000 431.650000 ;
      RECT 29.500000 430.350000 49.500000 431.650000 ;
      RECT 15.500000 430.350000 16.500000 431.650000 ;
      RECT 1157.500000 429.650000 1170.500000 430.350000 ;
      RECT 1107.500000 429.650000 1149.500000 430.350000 ;
      RECT 1057.500000 429.650000 1099.500000 430.350000 ;
      RECT 1007.500000 429.650000 1049.500000 430.350000 ;
      RECT 957.500000 429.650000 999.500000 430.350000 ;
      RECT 907.500000 429.650000 949.500000 430.350000 ;
      RECT 857.500000 429.650000 899.500000 430.350000 ;
      RECT 807.500000 429.650000 849.500000 430.350000 ;
      RECT 757.500000 429.650000 799.500000 430.350000 ;
      RECT 707.500000 429.650000 749.500000 430.350000 ;
      RECT 657.500000 429.650000 699.500000 430.350000 ;
      RECT 607.500000 429.650000 649.500000 430.350000 ;
      RECT 557.500000 429.650000 599.500000 430.350000 ;
      RECT 507.500000 429.650000 549.500000 430.350000 ;
      RECT 457.500000 429.650000 499.500000 430.350000 ;
      RECT 407.500000 429.650000 449.500000 430.350000 ;
      RECT 357.500000 429.650000 399.500000 430.350000 ;
      RECT 307.500000 429.650000 349.500000 430.350000 ;
      RECT 207.500000 429.650000 299.500000 430.350000 ;
      RECT 107.500000 429.650000 199.500000 430.350000 ;
      RECT 57.500000 429.650000 99.500000 430.350000 ;
      RECT 15.500000 429.650000 49.500000 430.350000 ;
      RECT 1183.500000 428.350000 1186.000000 431.650000 ;
      RECT 1169.500000 428.350000 1170.500000 429.650000 ;
      RECT 1116.500000 428.350000 1149.500000 429.650000 ;
      RECT 1107.500000 428.350000 1108.500000 429.650000 ;
      RECT 1066.500000 428.350000 1099.500000 429.650000 ;
      RECT 1057.500000 428.350000 1058.500000 429.650000 ;
      RECT 1016.500000 428.350000 1049.500000 429.650000 ;
      RECT 1007.500000 428.350000 1008.500000 429.650000 ;
      RECT 966.500000 428.350000 999.500000 429.650000 ;
      RECT 957.500000 428.350000 958.500000 429.650000 ;
      RECT 916.500000 428.350000 949.500000 429.650000 ;
      RECT 907.500000 428.350000 908.500000 429.650000 ;
      RECT 866.500000 428.350000 899.500000 429.650000 ;
      RECT 857.500000 428.350000 858.500000 429.650000 ;
      RECT 816.500000 428.350000 849.500000 429.650000 ;
      RECT 807.500000 428.350000 808.500000 429.650000 ;
      RECT 766.500000 428.350000 799.500000 429.650000 ;
      RECT 757.500000 428.350000 758.500000 429.650000 ;
      RECT 722.500000 428.350000 749.500000 429.650000 ;
      RECT 707.500000 428.350000 709.500000 429.650000 ;
      RECT 666.500000 428.350000 699.500000 429.650000 ;
      RECT 657.500000 428.350000 658.500000 429.650000 ;
      RECT 616.500000 428.350000 649.500000 429.650000 ;
      RECT 607.500000 428.350000 608.500000 429.650000 ;
      RECT 566.500000 428.350000 599.500000 429.650000 ;
      RECT 557.500000 428.350000 558.500000 429.650000 ;
      RECT 516.500000 428.350000 549.500000 429.650000 ;
      RECT 507.500000 428.350000 508.500000 429.650000 ;
      RECT 466.500000 428.350000 499.500000 429.650000 ;
      RECT 457.500000 428.350000 458.500000 429.650000 ;
      RECT 416.500000 428.350000 449.500000 429.650000 ;
      RECT 407.500000 428.350000 408.500000 429.650000 ;
      RECT 366.500000 428.350000 399.500000 429.650000 ;
      RECT 357.500000 428.350000 358.500000 429.650000 ;
      RECT 316.500000 428.350000 349.500000 429.650000 ;
      RECT 307.500000 428.350000 308.500000 429.650000 ;
      RECT 216.500000 428.350000 299.500000 429.650000 ;
      RECT 207.500000 428.350000 208.500000 429.650000 ;
      RECT 116.500000 428.350000 199.500000 429.650000 ;
      RECT 107.500000 428.350000 108.500000 429.650000 ;
      RECT 66.500000 428.350000 99.500000 429.650000 ;
      RECT 57.500000 428.350000 58.500000 429.650000 ;
      RECT 29.500000 428.350000 49.500000 429.650000 ;
      RECT 15.500000 428.350000 16.500000 429.650000 ;
      RECT 0.000000 428.350000 2.500000 431.650000 ;
      RECT 1169.500000 427.650000 1186.000000 428.350000 ;
      RECT 1116.500000 427.650000 1156.500000 428.350000 ;
      RECT 1066.500000 427.650000 1108.500000 428.350000 ;
      RECT 1016.500000 427.650000 1058.500000 428.350000 ;
      RECT 966.500000 427.650000 1008.500000 428.350000 ;
      RECT 916.500000 427.650000 958.500000 428.350000 ;
      RECT 866.500000 427.650000 908.500000 428.350000 ;
      RECT 816.500000 427.650000 858.500000 428.350000 ;
      RECT 766.500000 427.650000 808.500000 428.350000 ;
      RECT 722.500000 427.650000 758.500000 428.350000 ;
      RECT 666.500000 427.650000 709.500000 428.350000 ;
      RECT 616.500000 427.650000 658.500000 428.350000 ;
      RECT 566.500000 427.650000 608.500000 428.350000 ;
      RECT 516.500000 427.650000 558.500000 428.350000 ;
      RECT 466.500000 427.650000 508.500000 428.350000 ;
      RECT 416.500000 427.650000 458.500000 428.350000 ;
      RECT 366.500000 427.650000 408.500000 428.350000 ;
      RECT 316.500000 427.650000 358.500000 428.350000 ;
      RECT 216.500000 427.650000 308.500000 428.350000 ;
      RECT 116.500000 427.650000 208.500000 428.350000 ;
      RECT 66.500000 427.650000 108.500000 428.350000 ;
      RECT 29.500000 427.650000 58.500000 428.350000 ;
      RECT 0.000000 427.650000 16.500000 428.350000 ;
      RECT 1169.500000 426.350000 1170.500000 427.650000 ;
      RECT 1116.500000 426.350000 1149.500000 427.650000 ;
      RECT 1107.500000 426.350000 1108.500000 427.650000 ;
      RECT 1066.500000 426.350000 1099.500000 427.650000 ;
      RECT 1057.500000 426.350000 1058.500000 427.650000 ;
      RECT 1016.500000 426.350000 1049.500000 427.650000 ;
      RECT 1007.500000 426.350000 1008.500000 427.650000 ;
      RECT 966.500000 426.350000 999.500000 427.650000 ;
      RECT 957.500000 426.350000 958.500000 427.650000 ;
      RECT 916.500000 426.350000 949.500000 427.650000 ;
      RECT 907.500000 426.350000 908.500000 427.650000 ;
      RECT 866.500000 426.350000 899.500000 427.650000 ;
      RECT 857.500000 426.350000 858.500000 427.650000 ;
      RECT 816.500000 426.350000 849.500000 427.650000 ;
      RECT 807.500000 426.350000 808.500000 427.650000 ;
      RECT 766.500000 426.350000 799.500000 427.650000 ;
      RECT 757.500000 426.350000 758.500000 427.650000 ;
      RECT 722.500000 426.350000 749.500000 427.650000 ;
      RECT 707.500000 426.350000 709.500000 427.650000 ;
      RECT 666.500000 426.350000 699.500000 427.650000 ;
      RECT 657.500000 426.350000 658.500000 427.650000 ;
      RECT 616.500000 426.350000 649.500000 427.650000 ;
      RECT 607.500000 426.350000 608.500000 427.650000 ;
      RECT 566.500000 426.350000 599.500000 427.650000 ;
      RECT 557.500000 426.350000 558.500000 427.650000 ;
      RECT 516.500000 426.350000 549.500000 427.650000 ;
      RECT 507.500000 426.350000 508.500000 427.650000 ;
      RECT 466.500000 426.350000 499.500000 427.650000 ;
      RECT 457.500000 426.350000 458.500000 427.650000 ;
      RECT 416.500000 426.350000 449.500000 427.650000 ;
      RECT 407.500000 426.350000 408.500000 427.650000 ;
      RECT 366.500000 426.350000 399.500000 427.650000 ;
      RECT 357.500000 426.350000 358.500000 427.650000 ;
      RECT 316.500000 426.350000 349.500000 427.650000 ;
      RECT 307.500000 426.350000 308.500000 427.650000 ;
      RECT 216.500000 426.350000 299.500000 427.650000 ;
      RECT 207.500000 426.350000 208.500000 427.650000 ;
      RECT 116.500000 426.350000 199.500000 427.650000 ;
      RECT 107.500000 426.350000 108.500000 427.650000 ;
      RECT 66.500000 426.350000 99.500000 427.650000 ;
      RECT 57.500000 426.350000 58.500000 427.650000 ;
      RECT 29.500000 426.350000 49.500000 427.650000 ;
      RECT 15.500000 426.350000 16.500000 427.650000 ;
      RECT 1157.500000 425.650000 1170.500000 426.350000 ;
      RECT 1107.500000 425.650000 1149.500000 426.350000 ;
      RECT 1057.500000 425.650000 1099.500000 426.350000 ;
      RECT 1007.500000 425.650000 1049.500000 426.350000 ;
      RECT 957.500000 425.650000 999.500000 426.350000 ;
      RECT 907.500000 425.650000 949.500000 426.350000 ;
      RECT 857.500000 425.650000 899.500000 426.350000 ;
      RECT 807.500000 425.650000 849.500000 426.350000 ;
      RECT 757.500000 425.650000 799.500000 426.350000 ;
      RECT 707.500000 425.650000 749.500000 426.350000 ;
      RECT 657.500000 425.650000 699.500000 426.350000 ;
      RECT 607.500000 425.650000 649.500000 426.350000 ;
      RECT 557.500000 425.650000 599.500000 426.350000 ;
      RECT 507.500000 425.650000 549.500000 426.350000 ;
      RECT 457.500000 425.650000 499.500000 426.350000 ;
      RECT 407.500000 425.650000 449.500000 426.350000 ;
      RECT 357.500000 425.650000 399.500000 426.350000 ;
      RECT 307.500000 425.650000 349.500000 426.350000 ;
      RECT 207.500000 425.650000 299.500000 426.350000 ;
      RECT 107.500000 425.650000 199.500000 426.350000 ;
      RECT 57.500000 425.650000 99.500000 426.350000 ;
      RECT 15.500000 425.650000 49.500000 426.350000 ;
      RECT 1183.500000 424.350000 1186.000000 427.650000 ;
      RECT 1169.500000 424.350000 1170.500000 425.650000 ;
      RECT 1116.500000 424.350000 1149.500000 425.650000 ;
      RECT 1107.500000 424.350000 1108.500000 425.650000 ;
      RECT 1066.500000 424.350000 1099.500000 425.650000 ;
      RECT 1057.500000 424.350000 1058.500000 425.650000 ;
      RECT 1016.500000 424.350000 1049.500000 425.650000 ;
      RECT 1007.500000 424.350000 1008.500000 425.650000 ;
      RECT 966.500000 424.350000 999.500000 425.650000 ;
      RECT 957.500000 424.350000 958.500000 425.650000 ;
      RECT 916.500000 424.350000 949.500000 425.650000 ;
      RECT 907.500000 424.350000 908.500000 425.650000 ;
      RECT 866.500000 424.350000 899.500000 425.650000 ;
      RECT 857.500000 424.350000 858.500000 425.650000 ;
      RECT 816.500000 424.350000 849.500000 425.650000 ;
      RECT 807.500000 424.350000 808.500000 425.650000 ;
      RECT 766.500000 424.350000 799.500000 425.650000 ;
      RECT 757.500000 424.350000 758.500000 425.650000 ;
      RECT 722.500000 424.350000 749.500000 425.650000 ;
      RECT 707.500000 424.350000 709.500000 425.650000 ;
      RECT 666.500000 424.350000 699.500000 425.650000 ;
      RECT 657.500000 424.350000 658.500000 425.650000 ;
      RECT 616.500000 424.350000 649.500000 425.650000 ;
      RECT 607.500000 424.350000 608.500000 425.650000 ;
      RECT 566.500000 424.350000 599.500000 425.650000 ;
      RECT 557.500000 424.350000 558.500000 425.650000 ;
      RECT 516.500000 424.350000 549.500000 425.650000 ;
      RECT 507.500000 424.350000 508.500000 425.650000 ;
      RECT 466.500000 424.350000 499.500000 425.650000 ;
      RECT 457.500000 424.350000 458.500000 425.650000 ;
      RECT 416.500000 424.350000 449.500000 425.650000 ;
      RECT 407.500000 424.350000 408.500000 425.650000 ;
      RECT 366.500000 424.350000 399.500000 425.650000 ;
      RECT 357.500000 424.350000 358.500000 425.650000 ;
      RECT 316.500000 424.350000 349.500000 425.650000 ;
      RECT 307.500000 424.350000 308.500000 425.650000 ;
      RECT 216.500000 424.350000 299.500000 425.650000 ;
      RECT 207.500000 424.350000 208.500000 425.650000 ;
      RECT 116.500000 424.350000 199.500000 425.650000 ;
      RECT 107.500000 424.350000 108.500000 425.650000 ;
      RECT 66.500000 424.350000 99.500000 425.650000 ;
      RECT 57.500000 424.350000 58.500000 425.650000 ;
      RECT 29.500000 424.350000 49.500000 425.650000 ;
      RECT 15.500000 424.350000 16.500000 425.650000 ;
      RECT 0.000000 424.350000 2.500000 427.650000 ;
      RECT 1169.500000 423.650000 1186.000000 424.350000 ;
      RECT 1116.500000 423.650000 1156.500000 424.350000 ;
      RECT 1066.500000 423.650000 1108.500000 424.350000 ;
      RECT 1016.500000 423.650000 1058.500000 424.350000 ;
      RECT 966.500000 423.650000 1008.500000 424.350000 ;
      RECT 916.500000 423.650000 958.500000 424.350000 ;
      RECT 866.500000 423.650000 908.500000 424.350000 ;
      RECT 816.500000 423.650000 858.500000 424.350000 ;
      RECT 766.500000 423.650000 808.500000 424.350000 ;
      RECT 722.500000 423.650000 758.500000 424.350000 ;
      RECT 666.500000 423.650000 709.500000 424.350000 ;
      RECT 616.500000 423.650000 658.500000 424.350000 ;
      RECT 566.500000 423.650000 608.500000 424.350000 ;
      RECT 516.500000 423.650000 558.500000 424.350000 ;
      RECT 466.500000 423.650000 508.500000 424.350000 ;
      RECT 416.500000 423.650000 458.500000 424.350000 ;
      RECT 366.500000 423.650000 408.500000 424.350000 ;
      RECT 316.500000 423.650000 358.500000 424.350000 ;
      RECT 216.500000 423.650000 308.500000 424.350000 ;
      RECT 116.500000 423.650000 208.500000 424.350000 ;
      RECT 66.500000 423.650000 108.500000 424.350000 ;
      RECT 29.500000 423.650000 58.500000 424.350000 ;
      RECT 0.000000 423.650000 16.500000 424.350000 ;
      RECT 1169.500000 422.350000 1170.500000 423.650000 ;
      RECT 1116.500000 422.350000 1149.500000 423.650000 ;
      RECT 1107.500000 422.350000 1108.500000 423.650000 ;
      RECT 1066.500000 422.350000 1099.500000 423.650000 ;
      RECT 1057.500000 422.350000 1058.500000 423.650000 ;
      RECT 1016.500000 422.350000 1049.500000 423.650000 ;
      RECT 1007.500000 422.350000 1008.500000 423.650000 ;
      RECT 966.500000 422.350000 999.500000 423.650000 ;
      RECT 957.500000 422.350000 958.500000 423.650000 ;
      RECT 916.500000 422.350000 949.500000 423.650000 ;
      RECT 907.500000 422.350000 908.500000 423.650000 ;
      RECT 866.500000 422.350000 899.500000 423.650000 ;
      RECT 857.500000 422.350000 858.500000 423.650000 ;
      RECT 816.500000 422.350000 849.500000 423.650000 ;
      RECT 807.500000 422.350000 808.500000 423.650000 ;
      RECT 766.500000 422.350000 799.500000 423.650000 ;
      RECT 757.500000 422.350000 758.500000 423.650000 ;
      RECT 722.500000 422.350000 749.500000 423.650000 ;
      RECT 707.500000 422.350000 709.500000 423.650000 ;
      RECT 666.500000 422.350000 699.500000 423.650000 ;
      RECT 657.500000 422.350000 658.500000 423.650000 ;
      RECT 616.500000 422.350000 649.500000 423.650000 ;
      RECT 607.500000 422.350000 608.500000 423.650000 ;
      RECT 566.500000 422.350000 599.500000 423.650000 ;
      RECT 557.500000 422.350000 558.500000 423.650000 ;
      RECT 516.500000 422.350000 549.500000 423.650000 ;
      RECT 507.500000 422.350000 508.500000 423.650000 ;
      RECT 466.500000 422.350000 499.500000 423.650000 ;
      RECT 457.500000 422.350000 458.500000 423.650000 ;
      RECT 416.500000 422.350000 449.500000 423.650000 ;
      RECT 407.500000 422.350000 408.500000 423.650000 ;
      RECT 366.500000 422.350000 399.500000 423.650000 ;
      RECT 357.500000 422.350000 358.500000 423.650000 ;
      RECT 316.500000 422.350000 349.500000 423.650000 ;
      RECT 307.500000 422.350000 308.500000 423.650000 ;
      RECT 216.500000 422.350000 299.500000 423.650000 ;
      RECT 207.500000 422.350000 208.500000 423.650000 ;
      RECT 116.500000 422.350000 199.500000 423.650000 ;
      RECT 107.500000 422.350000 108.500000 423.650000 ;
      RECT 66.500000 422.350000 99.500000 423.650000 ;
      RECT 57.500000 422.350000 58.500000 423.650000 ;
      RECT 29.500000 422.350000 49.500000 423.650000 ;
      RECT 15.500000 422.350000 16.500000 423.650000 ;
      RECT 1157.500000 421.650000 1170.500000 422.350000 ;
      RECT 1107.500000 421.650000 1149.500000 422.350000 ;
      RECT 1057.500000 421.650000 1099.500000 422.350000 ;
      RECT 1007.500000 421.650000 1049.500000 422.350000 ;
      RECT 957.500000 421.650000 999.500000 422.350000 ;
      RECT 907.500000 421.650000 949.500000 422.350000 ;
      RECT 857.500000 421.650000 899.500000 422.350000 ;
      RECT 807.500000 421.650000 849.500000 422.350000 ;
      RECT 757.500000 421.650000 799.500000 422.350000 ;
      RECT 707.500000 421.650000 749.500000 422.350000 ;
      RECT 657.500000 421.650000 699.500000 422.350000 ;
      RECT 607.500000 421.650000 649.500000 422.350000 ;
      RECT 557.500000 421.650000 599.500000 422.350000 ;
      RECT 507.500000 421.650000 549.500000 422.350000 ;
      RECT 457.500000 421.650000 499.500000 422.350000 ;
      RECT 407.500000 421.650000 449.500000 422.350000 ;
      RECT 357.500000 421.650000 399.500000 422.350000 ;
      RECT 307.500000 421.650000 349.500000 422.350000 ;
      RECT 207.500000 421.650000 299.500000 422.350000 ;
      RECT 107.500000 421.650000 199.500000 422.350000 ;
      RECT 57.500000 421.650000 99.500000 422.350000 ;
      RECT 15.500000 421.650000 49.500000 422.350000 ;
      RECT 1183.500000 420.350000 1186.000000 423.650000 ;
      RECT 1169.500000 420.350000 1170.500000 421.650000 ;
      RECT 1116.500000 420.350000 1149.500000 421.650000 ;
      RECT 1107.500000 420.350000 1108.500000 421.650000 ;
      RECT 1066.500000 420.350000 1099.500000 421.650000 ;
      RECT 1057.500000 420.350000 1058.500000 421.650000 ;
      RECT 1016.500000 420.350000 1049.500000 421.650000 ;
      RECT 1007.500000 420.350000 1008.500000 421.650000 ;
      RECT 966.500000 420.350000 999.500000 421.650000 ;
      RECT 957.500000 420.350000 958.500000 421.650000 ;
      RECT 916.500000 420.350000 949.500000 421.650000 ;
      RECT 907.500000 420.350000 908.500000 421.650000 ;
      RECT 866.500000 420.350000 899.500000 421.650000 ;
      RECT 857.500000 420.350000 858.500000 421.650000 ;
      RECT 816.500000 420.350000 849.500000 421.650000 ;
      RECT 807.500000 420.350000 808.500000 421.650000 ;
      RECT 766.500000 420.350000 799.500000 421.650000 ;
      RECT 757.500000 420.350000 758.500000 421.650000 ;
      RECT 722.500000 420.350000 749.500000 421.650000 ;
      RECT 707.500000 420.350000 709.500000 421.650000 ;
      RECT 666.500000 420.350000 699.500000 421.650000 ;
      RECT 657.500000 420.350000 658.500000 421.650000 ;
      RECT 616.500000 420.350000 649.500000 421.650000 ;
      RECT 607.500000 420.350000 608.500000 421.650000 ;
      RECT 566.500000 420.350000 599.500000 421.650000 ;
      RECT 557.500000 420.350000 558.500000 421.650000 ;
      RECT 516.500000 420.350000 549.500000 421.650000 ;
      RECT 507.500000 420.350000 508.500000 421.650000 ;
      RECT 466.500000 420.350000 499.500000 421.650000 ;
      RECT 457.500000 420.350000 458.500000 421.650000 ;
      RECT 416.500000 420.350000 449.500000 421.650000 ;
      RECT 407.500000 420.350000 408.500000 421.650000 ;
      RECT 366.500000 420.350000 399.500000 421.650000 ;
      RECT 357.500000 420.350000 358.500000 421.650000 ;
      RECT 316.500000 420.350000 349.500000 421.650000 ;
      RECT 307.500000 420.350000 308.500000 421.650000 ;
      RECT 216.500000 420.350000 299.500000 421.650000 ;
      RECT 207.500000 420.350000 208.500000 421.650000 ;
      RECT 116.500000 420.350000 199.500000 421.650000 ;
      RECT 107.500000 420.350000 108.500000 421.650000 ;
      RECT 66.500000 420.350000 99.500000 421.650000 ;
      RECT 57.500000 420.350000 58.500000 421.650000 ;
      RECT 29.500000 420.350000 49.500000 421.650000 ;
      RECT 15.500000 420.350000 16.500000 421.650000 ;
      RECT 0.000000 420.350000 2.500000 423.650000 ;
      RECT 1169.500000 419.650000 1186.000000 420.350000 ;
      RECT 1116.500000 419.650000 1156.500000 420.350000 ;
      RECT 1066.500000 419.650000 1108.500000 420.350000 ;
      RECT 1016.500000 419.650000 1058.500000 420.350000 ;
      RECT 966.500000 419.650000 1008.500000 420.350000 ;
      RECT 916.500000 419.650000 958.500000 420.350000 ;
      RECT 866.500000 419.650000 908.500000 420.350000 ;
      RECT 816.500000 419.650000 858.500000 420.350000 ;
      RECT 766.500000 419.650000 808.500000 420.350000 ;
      RECT 722.500000 419.650000 758.500000 420.350000 ;
      RECT 666.500000 419.650000 709.500000 420.350000 ;
      RECT 616.500000 419.650000 658.500000 420.350000 ;
      RECT 566.500000 419.650000 608.500000 420.350000 ;
      RECT 516.500000 419.650000 558.500000 420.350000 ;
      RECT 466.500000 419.650000 508.500000 420.350000 ;
      RECT 366.500000 419.650000 408.500000 420.350000 ;
      RECT 316.500000 419.650000 358.500000 420.350000 ;
      RECT 216.500000 419.650000 308.500000 420.350000 ;
      RECT 116.500000 419.650000 208.500000 420.350000 ;
      RECT 66.500000 419.650000 108.500000 420.350000 ;
      RECT 29.500000 419.650000 58.500000 420.350000 ;
      RECT 0.000000 419.650000 16.500000 420.350000 ;
      RECT 416.500000 418.605000 458.500000 420.350000 ;
      RECT 1169.500000 418.350000 1170.500000 419.650000 ;
      RECT 1116.500000 418.350000 1149.500000 419.650000 ;
      RECT 1107.500000 418.350000 1108.500000 419.650000 ;
      RECT 1066.500000 418.350000 1099.500000 419.650000 ;
      RECT 1057.500000 418.350000 1058.500000 419.650000 ;
      RECT 1016.500000 418.350000 1049.500000 419.650000 ;
      RECT 1007.500000 418.350000 1008.500000 419.650000 ;
      RECT 966.500000 418.350000 999.500000 419.650000 ;
      RECT 957.500000 418.350000 958.500000 419.650000 ;
      RECT 916.500000 418.350000 949.500000 419.650000 ;
      RECT 907.500000 418.350000 908.500000 419.650000 ;
      RECT 866.500000 418.350000 899.500000 419.650000 ;
      RECT 857.500000 418.350000 858.500000 419.650000 ;
      RECT 816.500000 418.350000 849.500000 419.650000 ;
      RECT 807.500000 418.350000 808.500000 419.650000 ;
      RECT 766.500000 418.350000 799.500000 419.650000 ;
      RECT 757.500000 418.350000 758.500000 419.650000 ;
      RECT 722.500000 418.350000 749.500000 419.650000 ;
      RECT 707.500000 418.350000 709.500000 419.650000 ;
      RECT 666.500000 418.350000 699.500000 419.650000 ;
      RECT 657.500000 418.350000 658.500000 419.650000 ;
      RECT 616.500000 418.350000 649.500000 419.650000 ;
      RECT 607.500000 418.350000 608.500000 419.650000 ;
      RECT 566.500000 418.350000 599.500000 419.650000 ;
      RECT 557.500000 418.350000 558.500000 419.650000 ;
      RECT 516.500000 418.350000 549.500000 419.650000 ;
      RECT 507.500000 418.350000 508.500000 419.650000 ;
      RECT 466.500000 418.350000 499.500000 419.650000 ;
      RECT 457.500000 418.350000 458.500000 418.605000 ;
      RECT 416.500000 418.350000 449.500000 418.605000 ;
      RECT 407.500000 418.350000 408.500000 419.650000 ;
      RECT 366.500000 418.350000 399.500000 419.650000 ;
      RECT 357.500000 418.350000 358.500000 419.650000 ;
      RECT 316.500000 418.350000 349.500000 419.650000 ;
      RECT 307.500000 418.350000 308.500000 419.650000 ;
      RECT 216.500000 418.350000 299.500000 419.650000 ;
      RECT 207.500000 418.350000 208.500000 419.650000 ;
      RECT 116.500000 418.350000 199.500000 419.650000 ;
      RECT 107.500000 418.350000 108.500000 419.650000 ;
      RECT 66.500000 418.350000 99.500000 419.650000 ;
      RECT 57.500000 418.350000 58.500000 419.650000 ;
      RECT 29.500000 418.350000 49.500000 419.650000 ;
      RECT 15.500000 418.350000 16.500000 419.650000 ;
      RECT 1157.500000 417.650000 1170.500000 418.350000 ;
      RECT 1107.500000 417.650000 1149.500000 418.350000 ;
      RECT 1057.500000 417.650000 1099.500000 418.350000 ;
      RECT 1007.500000 417.650000 1049.500000 418.350000 ;
      RECT 957.500000 417.650000 999.500000 418.350000 ;
      RECT 907.500000 417.650000 949.500000 418.350000 ;
      RECT 857.500000 417.650000 899.500000 418.350000 ;
      RECT 807.500000 417.650000 849.500000 418.350000 ;
      RECT 757.500000 417.650000 799.500000 418.350000 ;
      RECT 707.500000 417.650000 749.500000 418.350000 ;
      RECT 657.500000 417.650000 699.500000 418.350000 ;
      RECT 607.500000 417.650000 649.500000 418.350000 ;
      RECT 557.500000 417.650000 599.500000 418.350000 ;
      RECT 507.500000 417.650000 549.500000 418.350000 ;
      RECT 407.500000 417.650000 449.500000 418.350000 ;
      RECT 357.500000 417.650000 399.500000 418.350000 ;
      RECT 307.500000 417.650000 349.500000 418.350000 ;
      RECT 207.500000 417.650000 299.500000 418.350000 ;
      RECT 107.500000 417.650000 199.500000 418.350000 ;
      RECT 57.500000 417.650000 99.500000 418.350000 ;
      RECT 15.500000 417.650000 49.500000 418.350000 ;
      RECT 1183.500000 416.350000 1186.000000 419.650000 ;
      RECT 1169.500000 416.350000 1170.500000 417.650000 ;
      RECT 1116.500000 416.350000 1149.500000 417.650000 ;
      RECT 1107.500000 416.350000 1108.500000 417.650000 ;
      RECT 1066.500000 416.350000 1099.500000 417.650000 ;
      RECT 1057.500000 416.350000 1058.500000 417.650000 ;
      RECT 1016.500000 416.350000 1049.500000 417.650000 ;
      RECT 1007.500000 416.350000 1008.500000 417.650000 ;
      RECT 966.500000 416.350000 999.500000 417.650000 ;
      RECT 957.500000 416.350000 958.500000 417.650000 ;
      RECT 916.500000 416.350000 949.500000 417.650000 ;
      RECT 907.500000 416.350000 908.500000 417.650000 ;
      RECT 866.500000 416.350000 899.500000 417.650000 ;
      RECT 857.500000 416.350000 858.500000 417.650000 ;
      RECT 816.500000 416.350000 849.500000 417.650000 ;
      RECT 807.500000 416.350000 808.500000 417.650000 ;
      RECT 766.500000 416.350000 799.500000 417.650000 ;
      RECT 757.500000 416.350000 758.500000 417.650000 ;
      RECT 720.000000 416.350000 749.500000 417.650000 ;
      RECT 707.500000 416.350000 712.000000 417.650000 ;
      RECT 666.500000 416.350000 699.500000 417.650000 ;
      RECT 657.500000 416.350000 658.500000 417.650000 ;
      RECT 616.500000 416.350000 649.500000 417.650000 ;
      RECT 607.500000 416.350000 608.500000 417.650000 ;
      RECT 566.500000 416.350000 599.500000 417.650000 ;
      RECT 557.500000 416.350000 558.500000 417.650000 ;
      RECT 516.500000 416.350000 549.500000 417.650000 ;
      RECT 507.500000 416.350000 508.500000 417.650000 ;
      RECT 457.500000 416.350000 499.500000 418.350000 ;
      RECT 407.500000 416.350000 408.500000 417.650000 ;
      RECT 366.500000 416.350000 399.500000 417.650000 ;
      RECT 357.500000 416.350000 358.500000 417.650000 ;
      RECT 316.500000 416.350000 349.500000 417.650000 ;
      RECT 307.500000 416.350000 308.500000 417.650000 ;
      RECT 216.500000 416.350000 299.500000 417.650000 ;
      RECT 207.500000 416.350000 208.500000 417.650000 ;
      RECT 116.500000 416.350000 199.500000 417.650000 ;
      RECT 107.500000 416.350000 108.500000 417.650000 ;
      RECT 66.500000 416.350000 99.500000 417.650000 ;
      RECT 57.500000 416.350000 58.500000 417.650000 ;
      RECT 29.500000 416.350000 49.500000 417.650000 ;
      RECT 15.500000 416.350000 16.500000 417.650000 ;
      RECT 0.000000 416.350000 2.500000 419.650000 ;
      RECT 1169.500000 415.650000 1186.000000 416.350000 ;
      RECT 1116.500000 415.650000 1156.500000 416.350000 ;
      RECT 1066.500000 415.650000 1108.500000 416.350000 ;
      RECT 1016.500000 415.650000 1058.500000 416.350000 ;
      RECT 966.500000 415.650000 1008.500000 416.350000 ;
      RECT 916.500000 415.650000 958.500000 416.350000 ;
      RECT 866.500000 415.650000 908.500000 416.350000 ;
      RECT 816.500000 415.650000 858.500000 416.350000 ;
      RECT 766.500000 415.650000 808.500000 416.350000 ;
      RECT 720.000000 415.650000 758.500000 416.350000 ;
      RECT 666.500000 415.650000 712.000000 416.350000 ;
      RECT 616.500000 415.650000 658.500000 416.350000 ;
      RECT 566.500000 415.650000 608.500000 416.350000 ;
      RECT 516.500000 415.650000 558.500000 416.350000 ;
      RECT 457.500000 415.650000 508.500000 416.350000 ;
      RECT 366.500000 415.650000 408.500000 416.350000 ;
      RECT 316.500000 415.650000 358.500000 416.350000 ;
      RECT 216.500000 415.650000 308.500000 416.350000 ;
      RECT 116.500000 415.650000 208.500000 416.350000 ;
      RECT 66.500000 415.650000 108.500000 416.350000 ;
      RECT 29.500000 415.650000 58.500000 416.350000 ;
      RECT 0.000000 415.650000 16.500000 416.350000 ;
      RECT 457.500000 414.605000 499.500000 415.650000 ;
      RECT 416.500000 414.605000 449.500000 417.650000 ;
      RECT 1169.500000 414.350000 1170.500000 415.650000 ;
      RECT 1116.500000 414.350000 1149.500000 415.650000 ;
      RECT 1107.500000 414.350000 1108.500000 415.650000 ;
      RECT 1066.500000 414.350000 1099.500000 415.650000 ;
      RECT 1057.500000 414.350000 1058.500000 415.650000 ;
      RECT 1016.500000 414.350000 1049.500000 415.650000 ;
      RECT 1007.500000 414.350000 1008.500000 415.650000 ;
      RECT 966.500000 414.350000 999.500000 415.650000 ;
      RECT 957.500000 414.350000 958.500000 415.650000 ;
      RECT 916.500000 414.350000 949.500000 415.650000 ;
      RECT 907.500000 414.350000 908.500000 415.650000 ;
      RECT 866.500000 414.350000 899.500000 415.650000 ;
      RECT 857.500000 414.350000 858.500000 415.650000 ;
      RECT 816.500000 414.350000 849.500000 415.650000 ;
      RECT 807.500000 414.350000 808.500000 415.650000 ;
      RECT 766.500000 414.350000 799.500000 415.650000 ;
      RECT 757.500000 414.350000 758.500000 415.650000 ;
      RECT 720.000000 414.350000 749.500000 415.650000 ;
      RECT 707.500000 414.350000 712.000000 415.650000 ;
      RECT 666.500000 414.350000 699.500000 415.650000 ;
      RECT 657.500000 414.350000 658.500000 415.650000 ;
      RECT 616.500000 414.350000 649.500000 415.650000 ;
      RECT 607.500000 414.350000 608.500000 415.650000 ;
      RECT 566.500000 414.350000 599.500000 415.650000 ;
      RECT 557.500000 414.350000 558.500000 415.650000 ;
      RECT 516.500000 414.350000 549.500000 415.650000 ;
      RECT 507.500000 414.350000 508.500000 415.650000 ;
      RECT 416.500000 414.350000 499.500000 414.605000 ;
      RECT 407.500000 414.350000 408.500000 415.650000 ;
      RECT 366.500000 414.350000 399.500000 415.650000 ;
      RECT 357.500000 414.350000 358.500000 415.650000 ;
      RECT 316.500000 414.350000 349.500000 415.650000 ;
      RECT 307.500000 414.350000 308.500000 415.650000 ;
      RECT 216.500000 414.350000 299.500000 415.650000 ;
      RECT 207.500000 414.350000 208.500000 415.650000 ;
      RECT 116.500000 414.350000 199.500000 415.650000 ;
      RECT 107.500000 414.350000 108.500000 415.650000 ;
      RECT 66.500000 414.350000 99.500000 415.650000 ;
      RECT 57.500000 414.350000 58.500000 415.650000 ;
      RECT 29.500000 414.350000 49.500000 415.650000 ;
      RECT 15.500000 414.350000 16.500000 415.650000 ;
      RECT 1157.500000 413.650000 1170.500000 414.350000 ;
      RECT 1107.500000 413.650000 1149.500000 414.350000 ;
      RECT 1057.500000 413.650000 1099.500000 414.350000 ;
      RECT 1007.500000 413.650000 1049.500000 414.350000 ;
      RECT 957.500000 413.650000 999.500000 414.350000 ;
      RECT 907.500000 413.650000 949.500000 414.350000 ;
      RECT 857.500000 413.650000 899.500000 414.350000 ;
      RECT 807.500000 413.650000 849.500000 414.350000 ;
      RECT 757.500000 413.650000 799.500000 414.350000 ;
      RECT 707.500000 413.650000 749.500000 414.350000 ;
      RECT 657.500000 413.650000 699.500000 414.350000 ;
      RECT 607.500000 413.650000 649.500000 414.350000 ;
      RECT 557.500000 413.650000 599.500000 414.350000 ;
      RECT 507.500000 413.650000 549.500000 414.350000 ;
      RECT 407.500000 413.650000 499.500000 414.350000 ;
      RECT 357.500000 413.650000 399.500000 414.350000 ;
      RECT 307.500000 413.650000 349.500000 414.350000 ;
      RECT 207.500000 413.650000 299.500000 414.350000 ;
      RECT 107.500000 413.650000 199.500000 414.350000 ;
      RECT 57.500000 413.650000 99.500000 414.350000 ;
      RECT 15.500000 413.650000 49.500000 414.350000 ;
      RECT 1183.500000 412.350000 1186.000000 415.650000 ;
      RECT 1169.500000 412.350000 1170.500000 413.650000 ;
      RECT 1116.500000 412.350000 1149.500000 413.650000 ;
      RECT 1107.500000 412.350000 1108.500000 413.650000 ;
      RECT 1066.500000 412.350000 1099.500000 413.650000 ;
      RECT 1057.500000 412.350000 1058.500000 413.650000 ;
      RECT 1016.500000 412.350000 1049.500000 413.650000 ;
      RECT 1007.500000 412.350000 1008.500000 413.650000 ;
      RECT 966.500000 412.350000 999.500000 413.650000 ;
      RECT 957.500000 412.350000 958.500000 413.650000 ;
      RECT 916.500000 412.350000 949.500000 413.650000 ;
      RECT 907.500000 412.350000 908.500000 413.650000 ;
      RECT 866.500000 412.350000 899.500000 413.650000 ;
      RECT 857.500000 412.350000 858.500000 413.650000 ;
      RECT 816.500000 412.350000 849.500000 413.650000 ;
      RECT 807.500000 412.350000 808.500000 413.650000 ;
      RECT 766.500000 412.350000 799.500000 413.650000 ;
      RECT 757.500000 412.350000 758.500000 413.650000 ;
      RECT 720.000000 412.350000 749.500000 413.650000 ;
      RECT 707.500000 412.350000 708.500000 413.650000 ;
      RECT 666.500000 412.350000 699.500000 413.650000 ;
      RECT 657.500000 412.350000 658.500000 413.650000 ;
      RECT 616.500000 412.350000 649.500000 413.650000 ;
      RECT 607.500000 412.350000 608.500000 413.650000 ;
      RECT 566.500000 412.350000 599.500000 413.650000 ;
      RECT 557.500000 412.350000 558.500000 413.650000 ;
      RECT 516.500000 412.350000 549.500000 413.650000 ;
      RECT 507.500000 412.350000 508.500000 413.650000 ;
      RECT 416.500000 412.350000 499.500000 413.650000 ;
      RECT 407.500000 412.350000 408.500000 413.650000 ;
      RECT 366.500000 412.350000 399.500000 413.650000 ;
      RECT 357.500000 412.350000 358.500000 413.650000 ;
      RECT 316.500000 412.350000 349.500000 413.650000 ;
      RECT 307.500000 412.350000 308.500000 413.650000 ;
      RECT 216.500000 412.350000 299.500000 413.650000 ;
      RECT 207.500000 412.350000 208.500000 413.650000 ;
      RECT 116.500000 412.350000 199.500000 413.650000 ;
      RECT 107.500000 412.350000 108.500000 413.650000 ;
      RECT 66.500000 412.350000 99.500000 413.650000 ;
      RECT 57.500000 412.350000 58.500000 413.650000 ;
      RECT 29.500000 412.350000 49.500000 413.650000 ;
      RECT 15.500000 412.350000 16.500000 413.650000 ;
      RECT 0.000000 412.350000 2.500000 415.650000 ;
      RECT 1169.500000 411.650000 1186.000000 412.350000 ;
      RECT 1116.500000 411.650000 1156.500000 412.350000 ;
      RECT 1066.500000 411.650000 1108.500000 412.350000 ;
      RECT 1016.500000 411.650000 1058.500000 412.350000 ;
      RECT 966.500000 411.650000 1008.500000 412.350000 ;
      RECT 916.500000 411.650000 958.500000 412.350000 ;
      RECT 866.500000 411.650000 908.500000 412.350000 ;
      RECT 816.500000 411.650000 858.500000 412.350000 ;
      RECT 766.500000 411.650000 808.500000 412.350000 ;
      RECT 720.000000 411.650000 758.500000 412.350000 ;
      RECT 666.500000 411.650000 708.500000 412.350000 ;
      RECT 616.500000 411.650000 658.500000 412.350000 ;
      RECT 566.500000 411.650000 608.500000 412.350000 ;
      RECT 516.500000 411.650000 558.500000 412.350000 ;
      RECT 416.500000 411.650000 508.500000 412.350000 ;
      RECT 366.500000 411.650000 408.500000 412.350000 ;
      RECT 316.500000 411.650000 358.500000 412.350000 ;
      RECT 216.500000 411.650000 308.500000 412.350000 ;
      RECT 116.500000 411.650000 208.500000 412.350000 ;
      RECT 66.500000 411.650000 108.500000 412.350000 ;
      RECT 29.500000 411.650000 58.500000 412.350000 ;
      RECT 0.000000 411.650000 16.500000 412.350000 ;
      RECT 1169.500000 410.350000 1170.500000 411.650000 ;
      RECT 1116.500000 410.350000 1149.500000 411.650000 ;
      RECT 1107.500000 410.350000 1108.500000 411.650000 ;
      RECT 1066.500000 410.350000 1099.500000 411.650000 ;
      RECT 1057.500000 410.350000 1058.500000 411.650000 ;
      RECT 1016.500000 410.350000 1049.500000 411.650000 ;
      RECT 1007.500000 410.350000 1008.500000 411.650000 ;
      RECT 966.500000 410.350000 999.500000 411.650000 ;
      RECT 957.500000 410.350000 958.500000 411.650000 ;
      RECT 916.500000 410.350000 949.500000 411.650000 ;
      RECT 907.500000 410.350000 908.500000 411.650000 ;
      RECT 866.500000 410.350000 899.500000 411.650000 ;
      RECT 857.500000 410.350000 858.500000 411.650000 ;
      RECT 816.500000 410.350000 849.500000 411.650000 ;
      RECT 807.500000 410.350000 808.500000 411.650000 ;
      RECT 766.500000 410.350000 799.500000 411.650000 ;
      RECT 757.500000 410.350000 758.500000 411.650000 ;
      RECT 720.000000 410.350000 749.500000 411.650000 ;
      RECT 707.500000 410.350000 708.500000 411.650000 ;
      RECT 666.500000 410.350000 699.500000 411.650000 ;
      RECT 657.500000 410.350000 658.500000 411.650000 ;
      RECT 616.500000 410.350000 649.500000 411.650000 ;
      RECT 607.500000 410.350000 608.500000 411.650000 ;
      RECT 566.500000 410.350000 599.500000 411.650000 ;
      RECT 557.500000 410.350000 558.500000 411.650000 ;
      RECT 516.500000 410.350000 549.500000 411.650000 ;
      RECT 507.500000 410.350000 508.500000 411.650000 ;
      RECT 416.500000 410.350000 499.500000 411.650000 ;
      RECT 407.500000 410.350000 408.500000 411.650000 ;
      RECT 366.500000 410.350000 399.500000 411.650000 ;
      RECT 357.500000 410.350000 358.500000 411.650000 ;
      RECT 316.500000 410.350000 349.500000 411.650000 ;
      RECT 307.500000 410.350000 308.500000 411.650000 ;
      RECT 216.500000 410.350000 299.500000 411.650000 ;
      RECT 207.500000 410.350000 208.500000 411.650000 ;
      RECT 116.500000 410.350000 199.500000 411.650000 ;
      RECT 107.500000 410.350000 108.500000 411.650000 ;
      RECT 66.500000 410.350000 99.500000 411.650000 ;
      RECT 57.500000 410.350000 58.500000 411.650000 ;
      RECT 29.500000 410.350000 49.500000 411.650000 ;
      RECT 15.500000 410.350000 16.500000 411.650000 ;
      RECT 1157.500000 409.650000 1170.500000 410.350000 ;
      RECT 1107.500000 409.650000 1149.500000 410.350000 ;
      RECT 1057.500000 409.650000 1099.500000 410.350000 ;
      RECT 1007.500000 409.650000 1049.500000 410.350000 ;
      RECT 957.500000 409.650000 999.500000 410.350000 ;
      RECT 907.500000 409.650000 949.500000 410.350000 ;
      RECT 857.500000 409.650000 899.500000 410.350000 ;
      RECT 807.500000 409.650000 849.500000 410.350000 ;
      RECT 757.500000 409.650000 799.500000 410.350000 ;
      RECT 707.500000 409.650000 749.500000 410.350000 ;
      RECT 657.500000 409.650000 699.500000 410.350000 ;
      RECT 607.500000 409.650000 649.500000 410.350000 ;
      RECT 557.500000 409.650000 599.500000 410.350000 ;
      RECT 507.500000 409.650000 549.500000 410.350000 ;
      RECT 407.500000 409.650000 499.500000 410.350000 ;
      RECT 357.500000 409.650000 399.500000 410.350000 ;
      RECT 307.500000 409.650000 349.500000 410.350000 ;
      RECT 207.500000 409.650000 299.500000 410.350000 ;
      RECT 107.500000 409.650000 199.500000 410.350000 ;
      RECT 57.500000 409.650000 99.500000 410.350000 ;
      RECT 15.500000 409.650000 49.500000 410.350000 ;
      RECT 1183.500000 408.350000 1186.000000 411.650000 ;
      RECT 1169.500000 408.350000 1170.500000 409.650000 ;
      RECT 1116.500000 408.350000 1149.500000 409.650000 ;
      RECT 1107.500000 408.350000 1108.500000 409.650000 ;
      RECT 1066.500000 408.350000 1099.500000 409.650000 ;
      RECT 1057.500000 408.350000 1058.500000 409.650000 ;
      RECT 1016.500000 408.350000 1049.500000 409.650000 ;
      RECT 1007.500000 408.350000 1008.500000 409.650000 ;
      RECT 966.500000 408.350000 999.500000 409.650000 ;
      RECT 957.500000 408.350000 958.500000 409.650000 ;
      RECT 916.500000 408.350000 949.500000 409.650000 ;
      RECT 907.500000 408.350000 908.500000 409.650000 ;
      RECT 866.500000 408.350000 899.500000 409.650000 ;
      RECT 857.500000 408.350000 858.500000 409.650000 ;
      RECT 816.500000 408.350000 849.500000 409.650000 ;
      RECT 807.500000 408.350000 808.500000 409.650000 ;
      RECT 766.500000 408.350000 799.500000 409.650000 ;
      RECT 757.500000 408.350000 758.500000 409.650000 ;
      RECT 716.500000 408.350000 749.500000 409.650000 ;
      RECT 707.500000 408.350000 708.500000 409.650000 ;
      RECT 666.500000 408.350000 699.500000 409.650000 ;
      RECT 657.500000 408.350000 658.500000 409.650000 ;
      RECT 616.500000 408.350000 649.500000 409.650000 ;
      RECT 607.500000 408.350000 608.500000 409.650000 ;
      RECT 566.500000 408.350000 599.500000 409.650000 ;
      RECT 557.500000 408.350000 558.500000 409.650000 ;
      RECT 516.500000 408.350000 549.500000 409.650000 ;
      RECT 507.500000 408.350000 508.500000 409.650000 ;
      RECT 416.500000 408.350000 499.500000 409.650000 ;
      RECT 407.500000 408.350000 408.500000 409.650000 ;
      RECT 366.500000 408.350000 399.500000 409.650000 ;
      RECT 357.500000 408.350000 358.500000 409.650000 ;
      RECT 316.500000 408.350000 349.500000 409.650000 ;
      RECT 307.500000 408.350000 308.500000 409.650000 ;
      RECT 216.500000 408.350000 299.500000 409.650000 ;
      RECT 207.500000 408.350000 208.500000 409.650000 ;
      RECT 116.500000 408.350000 199.500000 409.650000 ;
      RECT 107.500000 408.350000 108.500000 409.650000 ;
      RECT 66.500000 408.350000 99.500000 409.650000 ;
      RECT 57.500000 408.350000 58.500000 409.650000 ;
      RECT 29.500000 408.350000 49.500000 409.650000 ;
      RECT 15.500000 408.350000 16.500000 409.650000 ;
      RECT 0.000000 408.350000 2.500000 411.650000 ;
      RECT 1169.500000 407.650000 1186.000000 408.350000 ;
      RECT 1116.500000 407.650000 1156.500000 408.350000 ;
      RECT 1066.500000 407.650000 1108.500000 408.350000 ;
      RECT 1016.500000 407.650000 1058.500000 408.350000 ;
      RECT 966.500000 407.650000 1008.500000 408.350000 ;
      RECT 916.500000 407.650000 958.500000 408.350000 ;
      RECT 866.500000 407.650000 908.500000 408.350000 ;
      RECT 816.500000 407.650000 858.500000 408.350000 ;
      RECT 766.500000 407.650000 808.500000 408.350000 ;
      RECT 716.500000 407.650000 758.500000 408.350000 ;
      RECT 666.500000 407.650000 708.500000 408.350000 ;
      RECT 616.500000 407.650000 658.500000 408.350000 ;
      RECT 566.500000 407.650000 608.500000 408.350000 ;
      RECT 516.500000 407.650000 558.500000 408.350000 ;
      RECT 416.500000 407.650000 508.500000 408.350000 ;
      RECT 366.500000 407.650000 408.500000 408.350000 ;
      RECT 316.500000 407.650000 358.500000 408.350000 ;
      RECT 216.500000 407.650000 308.500000 408.350000 ;
      RECT 116.500000 407.650000 208.500000 408.350000 ;
      RECT 66.500000 407.650000 108.500000 408.350000 ;
      RECT 29.500000 407.650000 58.500000 408.350000 ;
      RECT 0.000000 407.650000 16.500000 408.350000 ;
      RECT 1169.500000 406.350000 1170.500000 407.650000 ;
      RECT 1116.500000 406.350000 1149.500000 407.650000 ;
      RECT 1107.500000 406.350000 1108.500000 407.650000 ;
      RECT 1066.500000 406.350000 1099.500000 407.650000 ;
      RECT 1057.500000 406.350000 1058.500000 407.650000 ;
      RECT 1016.500000 406.350000 1049.500000 407.650000 ;
      RECT 1007.500000 406.350000 1008.500000 407.650000 ;
      RECT 966.500000 406.350000 999.500000 407.650000 ;
      RECT 957.500000 406.350000 958.500000 407.650000 ;
      RECT 916.500000 406.350000 949.500000 407.650000 ;
      RECT 907.500000 406.350000 908.500000 407.650000 ;
      RECT 866.500000 406.350000 899.500000 407.650000 ;
      RECT 857.500000 406.350000 858.500000 407.650000 ;
      RECT 816.500000 406.350000 849.500000 407.650000 ;
      RECT 807.500000 406.350000 808.500000 407.650000 ;
      RECT 766.500000 406.350000 799.500000 407.650000 ;
      RECT 757.500000 406.350000 758.500000 407.650000 ;
      RECT 716.500000 406.350000 749.500000 407.650000 ;
      RECT 707.500000 406.350000 708.500000 407.650000 ;
      RECT 666.500000 406.350000 699.500000 407.650000 ;
      RECT 657.500000 406.350000 658.500000 407.650000 ;
      RECT 616.500000 406.350000 649.500000 407.650000 ;
      RECT 607.500000 406.350000 608.500000 407.650000 ;
      RECT 566.500000 406.350000 599.500000 407.650000 ;
      RECT 557.500000 406.350000 558.500000 407.650000 ;
      RECT 516.500000 406.350000 549.500000 407.650000 ;
      RECT 507.500000 406.350000 508.500000 407.650000 ;
      RECT 416.500000 406.350000 499.500000 407.650000 ;
      RECT 407.500000 406.350000 408.500000 407.650000 ;
      RECT 366.500000 406.350000 399.500000 407.650000 ;
      RECT 357.500000 406.350000 358.500000 407.650000 ;
      RECT 316.500000 406.350000 349.500000 407.650000 ;
      RECT 307.500000 406.350000 308.500000 407.650000 ;
      RECT 216.500000 406.350000 299.500000 407.650000 ;
      RECT 207.500000 406.350000 208.500000 407.650000 ;
      RECT 116.500000 406.350000 199.500000 407.650000 ;
      RECT 107.500000 406.350000 108.500000 407.650000 ;
      RECT 66.500000 406.350000 99.500000 407.650000 ;
      RECT 57.500000 406.350000 58.500000 407.650000 ;
      RECT 29.500000 406.350000 49.500000 407.650000 ;
      RECT 15.500000 406.350000 16.500000 407.650000 ;
      RECT 1157.500000 405.650000 1170.500000 406.350000 ;
      RECT 1107.500000 405.650000 1149.500000 406.350000 ;
      RECT 1057.500000 405.650000 1099.500000 406.350000 ;
      RECT 1007.500000 405.650000 1049.500000 406.350000 ;
      RECT 957.500000 405.650000 999.500000 406.350000 ;
      RECT 907.500000 405.650000 949.500000 406.350000 ;
      RECT 857.500000 405.650000 899.500000 406.350000 ;
      RECT 807.500000 405.650000 849.500000 406.350000 ;
      RECT 757.500000 405.650000 799.500000 406.350000 ;
      RECT 707.500000 405.650000 749.500000 406.350000 ;
      RECT 657.500000 405.650000 699.500000 406.350000 ;
      RECT 607.500000 405.650000 649.500000 406.350000 ;
      RECT 557.500000 405.650000 599.500000 406.350000 ;
      RECT 507.500000 405.650000 549.500000 406.350000 ;
      RECT 407.500000 405.650000 499.500000 406.350000 ;
      RECT 357.500000 405.650000 399.500000 406.350000 ;
      RECT 307.500000 405.650000 349.500000 406.350000 ;
      RECT 207.500000 405.650000 299.500000 406.350000 ;
      RECT 107.500000 405.650000 199.500000 406.350000 ;
      RECT 57.500000 405.650000 99.500000 406.350000 ;
      RECT 15.500000 405.650000 49.500000 406.350000 ;
      RECT 1183.500000 404.350000 1186.000000 407.650000 ;
      RECT 1169.500000 404.350000 1170.500000 405.650000 ;
      RECT 1116.500000 404.350000 1149.500000 405.650000 ;
      RECT 1107.500000 404.350000 1108.500000 405.650000 ;
      RECT 1066.500000 404.350000 1099.500000 405.650000 ;
      RECT 1057.500000 404.350000 1058.500000 405.650000 ;
      RECT 1016.500000 404.350000 1049.500000 405.650000 ;
      RECT 1007.500000 404.350000 1008.500000 405.650000 ;
      RECT 966.500000 404.350000 999.500000 405.650000 ;
      RECT 957.500000 404.350000 958.500000 405.650000 ;
      RECT 916.500000 404.350000 949.500000 405.650000 ;
      RECT 907.500000 404.350000 908.500000 405.650000 ;
      RECT 866.500000 404.350000 899.500000 405.650000 ;
      RECT 857.500000 404.350000 858.500000 405.650000 ;
      RECT 816.500000 404.350000 849.500000 405.650000 ;
      RECT 807.500000 404.350000 808.500000 405.650000 ;
      RECT 766.500000 404.350000 799.500000 405.650000 ;
      RECT 757.500000 404.350000 758.500000 405.650000 ;
      RECT 716.500000 404.350000 749.500000 405.650000 ;
      RECT 707.500000 404.350000 708.500000 405.650000 ;
      RECT 666.500000 404.350000 699.500000 405.650000 ;
      RECT 657.500000 404.350000 658.500000 405.650000 ;
      RECT 616.500000 404.350000 649.500000 405.650000 ;
      RECT 607.500000 404.350000 608.500000 405.650000 ;
      RECT 566.500000 404.350000 599.500000 405.650000 ;
      RECT 557.500000 404.350000 558.500000 405.650000 ;
      RECT 516.500000 404.350000 549.500000 405.650000 ;
      RECT 507.500000 404.350000 508.500000 405.650000 ;
      RECT 416.500000 404.350000 499.500000 405.650000 ;
      RECT 407.500000 404.350000 408.500000 405.650000 ;
      RECT 366.500000 404.350000 399.500000 405.650000 ;
      RECT 357.500000 404.350000 358.500000 405.650000 ;
      RECT 316.500000 404.350000 349.500000 405.650000 ;
      RECT 307.500000 404.350000 308.500000 405.650000 ;
      RECT 216.500000 404.350000 299.500000 405.650000 ;
      RECT 207.500000 404.350000 208.500000 405.650000 ;
      RECT 116.500000 404.350000 199.500000 405.650000 ;
      RECT 107.500000 404.350000 108.500000 405.650000 ;
      RECT 66.500000 404.350000 99.500000 405.650000 ;
      RECT 57.500000 404.350000 58.500000 405.650000 ;
      RECT 29.500000 404.350000 49.500000 405.650000 ;
      RECT 15.500000 404.350000 16.500000 405.650000 ;
      RECT 0.000000 404.350000 2.500000 407.650000 ;
      RECT 416.500000 403.730000 508.500000 404.350000 ;
      RECT 1169.500000 403.650000 1186.000000 404.350000 ;
      RECT 1116.500000 403.650000 1156.500000 404.350000 ;
      RECT 1066.500000 403.650000 1108.500000 404.350000 ;
      RECT 1016.500000 403.650000 1058.500000 404.350000 ;
      RECT 966.500000 403.650000 1008.500000 404.350000 ;
      RECT 916.500000 403.650000 958.500000 404.350000 ;
      RECT 866.500000 403.650000 908.500000 404.350000 ;
      RECT 816.500000 403.650000 858.500000 404.350000 ;
      RECT 766.500000 403.650000 808.500000 404.350000 ;
      RECT 716.500000 403.650000 758.500000 404.350000 ;
      RECT 666.500000 403.650000 708.500000 404.350000 ;
      RECT 616.500000 403.650000 658.500000 404.350000 ;
      RECT 566.500000 403.650000 608.500000 404.350000 ;
      RECT 516.500000 403.650000 558.500000 404.350000 ;
      RECT 466.500000 403.650000 508.500000 403.730000 ;
      RECT 366.500000 403.650000 408.500000 404.350000 ;
      RECT 316.500000 403.650000 358.500000 404.350000 ;
      RECT 216.500000 403.650000 308.500000 404.350000 ;
      RECT 116.500000 403.650000 208.500000 404.350000 ;
      RECT 66.500000 403.650000 108.500000 404.350000 ;
      RECT 29.500000 403.650000 58.500000 404.350000 ;
      RECT 0.000000 403.650000 16.500000 404.350000 ;
      RECT 1169.500000 402.350000 1170.500000 403.650000 ;
      RECT 1116.500000 402.350000 1149.500000 403.650000 ;
      RECT 1107.500000 402.350000 1108.500000 403.650000 ;
      RECT 1066.500000 402.350000 1099.500000 403.650000 ;
      RECT 1057.500000 402.350000 1058.500000 403.650000 ;
      RECT 1016.500000 402.350000 1049.500000 403.650000 ;
      RECT 1007.500000 402.350000 1008.500000 403.650000 ;
      RECT 966.500000 402.350000 999.500000 403.650000 ;
      RECT 957.500000 402.350000 958.500000 403.650000 ;
      RECT 916.500000 402.350000 949.500000 403.650000 ;
      RECT 907.500000 402.350000 908.500000 403.650000 ;
      RECT 866.500000 402.350000 899.500000 403.650000 ;
      RECT 857.500000 402.350000 858.500000 403.650000 ;
      RECT 816.500000 402.350000 849.500000 403.650000 ;
      RECT 807.500000 402.350000 808.500000 403.650000 ;
      RECT 766.500000 402.350000 799.500000 403.650000 ;
      RECT 757.500000 402.350000 758.500000 403.650000 ;
      RECT 716.500000 402.350000 749.500000 403.650000 ;
      RECT 707.500000 402.350000 708.500000 403.650000 ;
      RECT 666.500000 402.350000 699.500000 403.650000 ;
      RECT 657.500000 402.350000 658.500000 403.650000 ;
      RECT 616.500000 402.350000 649.500000 403.650000 ;
      RECT 607.500000 402.350000 608.500000 403.650000 ;
      RECT 566.500000 402.350000 599.500000 403.650000 ;
      RECT 557.500000 402.350000 558.500000 403.650000 ;
      RECT 516.500000 402.350000 549.500000 403.650000 ;
      RECT 507.500000 402.350000 508.500000 403.650000 ;
      RECT 416.500000 402.350000 458.500000 403.730000 ;
      RECT 407.500000 402.350000 408.500000 403.650000 ;
      RECT 366.500000 402.350000 399.500000 403.650000 ;
      RECT 357.500000 402.350000 358.500000 403.650000 ;
      RECT 316.500000 402.350000 349.500000 403.650000 ;
      RECT 307.500000 402.350000 308.500000 403.650000 ;
      RECT 216.500000 402.350000 249.500000 403.650000 ;
      RECT 207.500000 402.350000 208.500000 403.650000 ;
      RECT 116.500000 402.350000 149.500000 403.650000 ;
      RECT 107.500000 402.350000 108.500000 403.650000 ;
      RECT 66.500000 402.350000 99.500000 403.650000 ;
      RECT 57.500000 402.350000 58.500000 403.650000 ;
      RECT 29.500000 402.350000 49.500000 403.650000 ;
      RECT 15.500000 402.350000 16.500000 403.650000 ;
      RECT 1157.500000 401.650000 1170.500000 402.350000 ;
      RECT 1107.500000 401.650000 1149.500000 402.350000 ;
      RECT 1057.500000 401.650000 1099.500000 402.350000 ;
      RECT 1007.500000 401.650000 1049.500000 402.350000 ;
      RECT 957.500000 401.650000 999.500000 402.350000 ;
      RECT 907.500000 401.650000 949.500000 402.350000 ;
      RECT 857.500000 401.650000 899.500000 402.350000 ;
      RECT 807.500000 401.650000 849.500000 402.350000 ;
      RECT 757.500000 401.650000 799.500000 402.350000 ;
      RECT 707.500000 401.650000 749.500000 402.350000 ;
      RECT 657.500000 401.650000 699.500000 402.350000 ;
      RECT 607.500000 401.650000 649.500000 402.350000 ;
      RECT 557.500000 401.650000 599.500000 402.350000 ;
      RECT 507.500000 401.650000 549.500000 402.350000 ;
      RECT 407.500000 401.650000 458.500000 402.350000 ;
      RECT 357.500000 401.650000 399.500000 402.350000 ;
      RECT 307.500000 401.650000 349.500000 402.350000 ;
      RECT 257.500000 401.650000 299.500000 403.650000 ;
      RECT 207.500000 401.650000 249.500000 402.350000 ;
      RECT 157.500000 401.650000 199.500000 403.650000 ;
      RECT 107.500000 401.650000 149.500000 402.350000 ;
      RECT 57.500000 401.650000 99.500000 402.350000 ;
      RECT 15.500000 401.650000 49.500000 402.350000 ;
      RECT 1183.500000 400.350000 1186.000000 403.650000 ;
      RECT 1169.500000 400.350000 1170.500000 401.650000 ;
      RECT 1116.500000 400.350000 1149.500000 401.650000 ;
      RECT 1107.500000 400.350000 1108.500000 401.650000 ;
      RECT 1066.500000 400.350000 1099.500000 401.650000 ;
      RECT 1057.500000 400.350000 1058.500000 401.650000 ;
      RECT 1016.500000 400.350000 1049.500000 401.650000 ;
      RECT 1007.500000 400.350000 1008.500000 401.650000 ;
      RECT 966.500000 400.350000 999.500000 401.650000 ;
      RECT 957.500000 400.350000 958.500000 401.650000 ;
      RECT 916.500000 400.350000 949.500000 401.650000 ;
      RECT 907.500000 400.350000 908.500000 401.650000 ;
      RECT 866.500000 400.350000 899.500000 401.650000 ;
      RECT 857.500000 400.350000 858.500000 401.650000 ;
      RECT 816.500000 400.350000 849.500000 401.650000 ;
      RECT 807.500000 400.350000 808.500000 401.650000 ;
      RECT 766.500000 400.350000 799.500000 401.650000 ;
      RECT 757.500000 400.350000 758.500000 401.650000 ;
      RECT 716.500000 400.350000 749.500000 401.650000 ;
      RECT 707.500000 400.350000 708.500000 401.650000 ;
      RECT 666.500000 400.350000 699.500000 401.650000 ;
      RECT 657.500000 400.350000 658.500000 401.650000 ;
      RECT 616.500000 400.350000 649.500000 401.650000 ;
      RECT 607.500000 400.350000 608.500000 401.650000 ;
      RECT 566.500000 400.350000 599.500000 401.650000 ;
      RECT 557.500000 400.350000 558.500000 401.650000 ;
      RECT 516.500000 400.350000 549.500000 401.650000 ;
      RECT 507.500000 400.350000 508.500000 401.650000 ;
      RECT 466.500000 400.350000 499.500000 403.650000 ;
      RECT 407.500000 400.350000 408.500000 401.650000 ;
      RECT 366.500000 400.350000 399.500000 401.650000 ;
      RECT 357.500000 400.350000 358.500000 401.650000 ;
      RECT 316.500000 400.350000 349.500000 401.650000 ;
      RECT 307.500000 400.350000 308.500000 401.650000 ;
      RECT 266.500000 400.350000 299.500000 401.650000 ;
      RECT 257.500000 400.350000 258.500000 401.650000 ;
      RECT 216.500000 400.350000 249.500000 401.650000 ;
      RECT 207.500000 400.350000 208.500000 401.650000 ;
      RECT 166.500000 400.350000 199.500000 401.650000 ;
      RECT 157.500000 400.350000 158.500000 401.650000 ;
      RECT 116.500000 400.350000 149.500000 401.650000 ;
      RECT 107.500000 400.350000 108.500000 401.650000 ;
      RECT 66.500000 400.350000 99.500000 401.650000 ;
      RECT 57.500000 400.350000 58.500000 401.650000 ;
      RECT 29.500000 400.350000 49.500000 401.650000 ;
      RECT 15.500000 400.350000 16.500000 401.650000 ;
      RECT 0.000000 400.350000 2.500000 403.650000 ;
      RECT 466.500000 399.730000 508.500000 400.350000 ;
      RECT 416.500000 399.730000 458.500000 401.650000 ;
      RECT 1169.500000 399.650000 1186.000000 400.350000 ;
      RECT 1116.500000 399.650000 1156.500000 400.350000 ;
      RECT 1066.500000 399.650000 1108.500000 400.350000 ;
      RECT 1016.500000 399.650000 1058.500000 400.350000 ;
      RECT 966.500000 399.650000 1008.500000 400.350000 ;
      RECT 916.500000 399.650000 958.500000 400.350000 ;
      RECT 866.500000 399.650000 908.500000 400.350000 ;
      RECT 816.500000 399.650000 858.500000 400.350000 ;
      RECT 766.500000 399.650000 808.500000 400.350000 ;
      RECT 716.500000 399.650000 758.500000 400.350000 ;
      RECT 666.500000 399.650000 708.500000 400.350000 ;
      RECT 616.500000 399.650000 658.500000 400.350000 ;
      RECT 566.500000 399.650000 608.500000 400.350000 ;
      RECT 516.500000 399.650000 558.500000 400.350000 ;
      RECT 416.500000 399.650000 508.500000 399.730000 ;
      RECT 366.500000 399.650000 408.500000 400.350000 ;
      RECT 316.500000 399.650000 358.500000 400.350000 ;
      RECT 266.500000 399.650000 308.500000 400.350000 ;
      RECT 216.500000 399.650000 258.500000 400.350000 ;
      RECT 166.500000 399.650000 208.500000 400.350000 ;
      RECT 116.500000 399.650000 158.500000 400.350000 ;
      RECT 66.500000 399.650000 108.500000 400.350000 ;
      RECT 29.500000 399.650000 58.500000 400.350000 ;
      RECT 0.000000 399.650000 16.500000 400.350000 ;
      RECT 1169.500000 398.350000 1170.500000 399.650000 ;
      RECT 1116.500000 398.350000 1149.500000 399.650000 ;
      RECT 1107.500000 398.350000 1108.500000 399.650000 ;
      RECT 1066.500000 398.350000 1099.500000 399.650000 ;
      RECT 1057.500000 398.350000 1058.500000 399.650000 ;
      RECT 1016.500000 398.350000 1049.500000 399.650000 ;
      RECT 1007.500000 398.350000 1008.500000 399.650000 ;
      RECT 966.500000 398.350000 999.500000 399.650000 ;
      RECT 957.500000 398.350000 958.500000 399.650000 ;
      RECT 916.500000 398.350000 949.500000 399.650000 ;
      RECT 907.500000 398.350000 908.500000 399.650000 ;
      RECT 866.500000 398.350000 899.500000 399.650000 ;
      RECT 857.500000 398.350000 858.500000 399.650000 ;
      RECT 816.500000 398.350000 849.500000 399.650000 ;
      RECT 807.500000 398.350000 808.500000 399.650000 ;
      RECT 766.500000 398.350000 799.500000 399.650000 ;
      RECT 757.500000 398.350000 758.500000 399.650000 ;
      RECT 716.500000 398.350000 749.500000 399.650000 ;
      RECT 707.500000 398.350000 708.500000 399.650000 ;
      RECT 666.500000 398.350000 699.500000 399.650000 ;
      RECT 657.500000 398.350000 658.500000 399.650000 ;
      RECT 616.500000 398.350000 649.500000 399.650000 ;
      RECT 607.500000 398.350000 608.500000 399.650000 ;
      RECT 566.500000 398.350000 599.500000 399.650000 ;
      RECT 557.500000 398.350000 558.500000 399.650000 ;
      RECT 516.500000 398.350000 549.500000 399.650000 ;
      RECT 507.500000 398.350000 508.500000 399.650000 ;
      RECT 416.500000 398.350000 449.500000 399.650000 ;
      RECT 407.500000 398.350000 408.500000 399.650000 ;
      RECT 366.500000 398.350000 399.500000 399.650000 ;
      RECT 357.500000 398.350000 358.500000 399.650000 ;
      RECT 316.500000 398.350000 349.500000 399.650000 ;
      RECT 307.500000 398.350000 308.500000 399.650000 ;
      RECT 266.500000 398.350000 299.500000 399.650000 ;
      RECT 257.500000 398.350000 258.500000 399.650000 ;
      RECT 216.500000 398.350000 249.500000 399.650000 ;
      RECT 207.500000 398.350000 208.500000 399.650000 ;
      RECT 166.500000 398.350000 199.500000 399.650000 ;
      RECT 157.500000 398.350000 158.500000 399.650000 ;
      RECT 116.500000 398.350000 149.500000 399.650000 ;
      RECT 107.500000 398.350000 108.500000 399.650000 ;
      RECT 66.500000 398.350000 99.500000 399.650000 ;
      RECT 57.500000 398.350000 58.500000 399.650000 ;
      RECT 29.500000 398.350000 49.500000 399.650000 ;
      RECT 15.500000 398.350000 16.500000 399.650000 ;
      RECT 1157.500000 397.650000 1170.500000 398.350000 ;
      RECT 1107.500000 397.650000 1149.500000 398.350000 ;
      RECT 1057.500000 397.650000 1099.500000 398.350000 ;
      RECT 1007.500000 397.650000 1049.500000 398.350000 ;
      RECT 957.500000 397.650000 999.500000 398.350000 ;
      RECT 907.500000 397.650000 949.500000 398.350000 ;
      RECT 857.500000 397.650000 899.500000 398.350000 ;
      RECT 807.500000 397.650000 849.500000 398.350000 ;
      RECT 757.500000 397.650000 799.500000 398.350000 ;
      RECT 707.500000 397.650000 749.500000 398.350000 ;
      RECT 657.500000 397.650000 699.500000 398.350000 ;
      RECT 607.500000 397.650000 649.500000 398.350000 ;
      RECT 557.500000 397.650000 599.500000 398.350000 ;
      RECT 507.500000 397.650000 549.500000 398.350000 ;
      RECT 457.500000 397.650000 499.500000 399.650000 ;
      RECT 407.500000 397.650000 449.500000 398.350000 ;
      RECT 357.500000 397.650000 399.500000 398.350000 ;
      RECT 307.500000 397.650000 349.500000 398.350000 ;
      RECT 257.500000 397.650000 299.500000 398.350000 ;
      RECT 207.500000 397.650000 249.500000 398.350000 ;
      RECT 157.500000 397.650000 199.500000 398.350000 ;
      RECT 107.500000 397.650000 149.500000 398.350000 ;
      RECT 57.500000 397.650000 99.500000 398.350000 ;
      RECT 15.500000 397.650000 49.500000 398.350000 ;
      RECT 1183.500000 396.350000 1186.000000 399.650000 ;
      RECT 1169.500000 396.350000 1170.500000 397.650000 ;
      RECT 1116.500000 396.350000 1149.500000 397.650000 ;
      RECT 1107.500000 396.350000 1108.500000 397.650000 ;
      RECT 1066.500000 396.350000 1099.500000 397.650000 ;
      RECT 1057.500000 396.350000 1058.500000 397.650000 ;
      RECT 1016.500000 396.350000 1049.500000 397.650000 ;
      RECT 1007.500000 396.350000 1008.500000 397.650000 ;
      RECT 966.500000 396.350000 999.500000 397.650000 ;
      RECT 957.500000 396.350000 958.500000 397.650000 ;
      RECT 916.500000 396.350000 949.500000 397.650000 ;
      RECT 907.500000 396.350000 908.500000 397.650000 ;
      RECT 866.500000 396.350000 899.500000 397.650000 ;
      RECT 857.500000 396.350000 858.500000 397.650000 ;
      RECT 816.500000 396.350000 849.500000 397.650000 ;
      RECT 807.500000 396.350000 808.500000 397.650000 ;
      RECT 766.500000 396.350000 799.500000 397.650000 ;
      RECT 757.500000 396.350000 758.500000 397.650000 ;
      RECT 716.500000 396.350000 749.500000 397.650000 ;
      RECT 707.500000 396.350000 708.500000 397.650000 ;
      RECT 666.500000 396.350000 699.500000 397.650000 ;
      RECT 657.500000 396.350000 658.500000 397.650000 ;
      RECT 616.500000 396.350000 649.500000 397.650000 ;
      RECT 607.500000 396.350000 608.500000 397.650000 ;
      RECT 566.500000 396.350000 599.500000 397.650000 ;
      RECT 557.500000 396.350000 558.500000 397.650000 ;
      RECT 516.500000 396.350000 549.500000 397.650000 ;
      RECT 507.500000 396.350000 508.500000 397.650000 ;
      RECT 466.500000 396.350000 499.500000 397.650000 ;
      RECT 457.500000 396.350000 458.500000 397.650000 ;
      RECT 416.500000 396.350000 449.500000 397.650000 ;
      RECT 407.500000 396.350000 408.500000 397.650000 ;
      RECT 366.500000 396.350000 399.500000 397.650000 ;
      RECT 357.500000 396.350000 358.500000 397.650000 ;
      RECT 316.500000 396.350000 349.500000 397.650000 ;
      RECT 307.500000 396.350000 308.500000 397.650000 ;
      RECT 266.500000 396.350000 299.500000 397.650000 ;
      RECT 257.500000 396.350000 258.500000 397.650000 ;
      RECT 216.500000 396.350000 249.500000 397.650000 ;
      RECT 207.500000 396.350000 208.500000 397.650000 ;
      RECT 166.500000 396.350000 199.500000 397.650000 ;
      RECT 157.500000 396.350000 158.500000 397.650000 ;
      RECT 116.500000 396.350000 149.500000 397.650000 ;
      RECT 107.500000 396.350000 108.500000 397.650000 ;
      RECT 66.500000 396.350000 99.500000 397.650000 ;
      RECT 57.500000 396.350000 58.500000 397.650000 ;
      RECT 29.500000 396.350000 49.500000 397.650000 ;
      RECT 15.500000 396.350000 16.500000 397.650000 ;
      RECT 0.000000 396.350000 2.500000 399.650000 ;
      RECT 1169.500000 395.650000 1186.000000 396.350000 ;
      RECT 1116.500000 395.650000 1156.500000 396.350000 ;
      RECT 1066.500000 395.650000 1108.500000 396.350000 ;
      RECT 1016.500000 395.650000 1058.500000 396.350000 ;
      RECT 966.500000 395.650000 1008.500000 396.350000 ;
      RECT 916.500000 395.650000 958.500000 396.350000 ;
      RECT 866.500000 395.650000 908.500000 396.350000 ;
      RECT 816.500000 395.650000 858.500000 396.350000 ;
      RECT 766.500000 395.650000 808.500000 396.350000 ;
      RECT 716.500000 395.650000 758.500000 396.350000 ;
      RECT 666.500000 395.650000 708.500000 396.350000 ;
      RECT 616.500000 395.650000 658.500000 396.350000 ;
      RECT 566.500000 395.650000 608.500000 396.350000 ;
      RECT 516.500000 395.650000 558.500000 396.350000 ;
      RECT 466.500000 395.650000 508.500000 396.350000 ;
      RECT 416.500000 395.650000 458.500000 396.350000 ;
      RECT 366.500000 395.650000 408.500000 396.350000 ;
      RECT 316.500000 395.650000 358.500000 396.350000 ;
      RECT 266.500000 395.650000 308.500000 396.350000 ;
      RECT 216.500000 395.650000 258.500000 396.350000 ;
      RECT 166.500000 395.650000 208.500000 396.350000 ;
      RECT 116.500000 395.650000 158.500000 396.350000 ;
      RECT 66.500000 395.650000 108.500000 396.350000 ;
      RECT 29.500000 395.650000 58.500000 396.350000 ;
      RECT 0.000000 395.650000 16.500000 396.350000 ;
      RECT 1169.500000 394.350000 1170.500000 395.650000 ;
      RECT 1116.500000 394.350000 1149.500000 395.650000 ;
      RECT 1107.500000 394.350000 1108.500000 395.650000 ;
      RECT 1066.500000 394.350000 1099.500000 395.650000 ;
      RECT 1057.500000 394.350000 1058.500000 395.650000 ;
      RECT 1016.500000 394.350000 1049.500000 395.650000 ;
      RECT 1007.500000 394.350000 1008.500000 395.650000 ;
      RECT 966.500000 394.350000 999.500000 395.650000 ;
      RECT 957.500000 394.350000 958.500000 395.650000 ;
      RECT 916.500000 394.350000 949.500000 395.650000 ;
      RECT 907.500000 394.350000 908.500000 395.650000 ;
      RECT 866.500000 394.350000 899.500000 395.650000 ;
      RECT 857.500000 394.350000 858.500000 395.650000 ;
      RECT 816.500000 394.350000 849.500000 395.650000 ;
      RECT 807.500000 394.350000 808.500000 395.650000 ;
      RECT 766.500000 394.350000 799.500000 395.650000 ;
      RECT 757.500000 394.350000 758.500000 395.650000 ;
      RECT 716.500000 394.350000 749.500000 395.650000 ;
      RECT 707.500000 394.350000 708.500000 395.650000 ;
      RECT 666.500000 394.350000 699.500000 395.650000 ;
      RECT 657.500000 394.350000 658.500000 395.650000 ;
      RECT 616.500000 394.350000 649.500000 395.650000 ;
      RECT 607.500000 394.350000 608.500000 395.650000 ;
      RECT 566.500000 394.350000 599.500000 395.650000 ;
      RECT 557.500000 394.350000 558.500000 395.650000 ;
      RECT 516.500000 394.350000 549.500000 395.650000 ;
      RECT 507.500000 394.350000 508.500000 395.650000 ;
      RECT 466.500000 394.350000 499.500000 395.650000 ;
      RECT 457.500000 394.350000 458.500000 395.650000 ;
      RECT 416.500000 394.350000 449.500000 395.650000 ;
      RECT 407.500000 394.350000 408.500000 395.650000 ;
      RECT 366.500000 394.350000 399.500000 395.650000 ;
      RECT 357.500000 394.350000 358.500000 395.650000 ;
      RECT 316.500000 394.350000 349.500000 395.650000 ;
      RECT 307.500000 394.350000 308.500000 395.650000 ;
      RECT 266.500000 394.350000 299.500000 395.650000 ;
      RECT 257.500000 394.350000 258.500000 395.650000 ;
      RECT 216.500000 394.350000 249.500000 395.650000 ;
      RECT 207.500000 394.350000 208.500000 395.650000 ;
      RECT 166.500000 394.350000 199.500000 395.650000 ;
      RECT 157.500000 394.350000 158.500000 395.650000 ;
      RECT 116.500000 394.350000 149.500000 395.650000 ;
      RECT 107.500000 394.350000 108.500000 395.650000 ;
      RECT 66.500000 394.350000 99.500000 395.650000 ;
      RECT 57.500000 394.350000 58.500000 395.650000 ;
      RECT 29.500000 394.350000 49.500000 395.650000 ;
      RECT 15.500000 394.350000 16.500000 395.650000 ;
      RECT 1157.500000 393.650000 1170.500000 394.350000 ;
      RECT 1107.500000 393.650000 1149.500000 394.350000 ;
      RECT 1057.500000 393.650000 1099.500000 394.350000 ;
      RECT 1007.500000 393.650000 1049.500000 394.350000 ;
      RECT 957.500000 393.650000 999.500000 394.350000 ;
      RECT 907.500000 393.650000 949.500000 394.350000 ;
      RECT 857.500000 393.650000 899.500000 394.350000 ;
      RECT 807.500000 393.650000 849.500000 394.350000 ;
      RECT 757.500000 393.650000 799.500000 394.350000 ;
      RECT 707.500000 393.650000 749.500000 394.350000 ;
      RECT 657.500000 393.650000 699.500000 394.350000 ;
      RECT 607.500000 393.650000 649.500000 394.350000 ;
      RECT 557.500000 393.650000 599.500000 394.350000 ;
      RECT 507.500000 393.650000 549.500000 394.350000 ;
      RECT 457.500000 393.650000 499.500000 394.350000 ;
      RECT 407.500000 393.650000 449.500000 394.350000 ;
      RECT 357.500000 393.650000 399.500000 394.350000 ;
      RECT 307.500000 393.650000 349.500000 394.350000 ;
      RECT 257.500000 393.650000 299.500000 394.350000 ;
      RECT 207.500000 393.650000 249.500000 394.350000 ;
      RECT 157.500000 393.650000 199.500000 394.350000 ;
      RECT 107.500000 393.650000 149.500000 394.350000 ;
      RECT 57.500000 393.650000 99.500000 394.350000 ;
      RECT 15.500000 393.650000 49.500000 394.350000 ;
      RECT 1183.500000 392.350000 1186.000000 395.650000 ;
      RECT 1169.500000 392.350000 1170.500000 393.650000 ;
      RECT 1116.500000 392.350000 1149.500000 393.650000 ;
      RECT 1107.500000 392.350000 1108.500000 393.650000 ;
      RECT 1066.500000 392.350000 1099.500000 393.650000 ;
      RECT 1057.500000 392.350000 1058.500000 393.650000 ;
      RECT 1016.500000 392.350000 1049.500000 393.650000 ;
      RECT 1007.500000 392.350000 1008.500000 393.650000 ;
      RECT 966.500000 392.350000 999.500000 393.650000 ;
      RECT 957.500000 392.350000 958.500000 393.650000 ;
      RECT 916.500000 392.350000 949.500000 393.650000 ;
      RECT 907.500000 392.350000 908.500000 393.650000 ;
      RECT 866.500000 392.350000 899.500000 393.650000 ;
      RECT 857.500000 392.350000 858.500000 393.650000 ;
      RECT 816.500000 392.350000 849.500000 393.650000 ;
      RECT 807.500000 392.350000 808.500000 393.650000 ;
      RECT 766.500000 392.350000 799.500000 393.650000 ;
      RECT 757.500000 392.350000 758.500000 393.650000 ;
      RECT 716.500000 392.350000 749.500000 393.650000 ;
      RECT 707.500000 392.350000 708.500000 393.650000 ;
      RECT 666.500000 392.350000 699.500000 393.650000 ;
      RECT 657.500000 392.350000 658.500000 393.650000 ;
      RECT 616.500000 392.350000 649.500000 393.650000 ;
      RECT 607.500000 392.350000 608.500000 393.650000 ;
      RECT 566.500000 392.350000 599.500000 393.650000 ;
      RECT 557.500000 392.350000 558.500000 393.650000 ;
      RECT 516.500000 392.350000 549.500000 393.650000 ;
      RECT 507.500000 392.350000 508.500000 393.650000 ;
      RECT 466.500000 392.350000 499.500000 393.650000 ;
      RECT 457.500000 392.350000 458.500000 393.650000 ;
      RECT 416.500000 392.350000 449.500000 393.650000 ;
      RECT 407.500000 392.350000 408.500000 393.650000 ;
      RECT 366.500000 392.350000 399.500000 393.650000 ;
      RECT 357.500000 392.350000 358.500000 393.650000 ;
      RECT 316.500000 392.350000 349.500000 393.650000 ;
      RECT 307.500000 392.350000 308.500000 393.650000 ;
      RECT 266.500000 392.350000 299.500000 393.650000 ;
      RECT 257.500000 392.350000 258.500000 393.650000 ;
      RECT 216.500000 392.350000 249.500000 393.650000 ;
      RECT 207.500000 392.350000 208.500000 393.650000 ;
      RECT 166.500000 392.350000 199.500000 393.650000 ;
      RECT 157.500000 392.350000 158.500000 393.650000 ;
      RECT 116.500000 392.350000 149.500000 393.650000 ;
      RECT 107.500000 392.350000 108.500000 393.650000 ;
      RECT 66.500000 392.350000 99.500000 393.650000 ;
      RECT 57.500000 392.350000 58.500000 393.650000 ;
      RECT 29.500000 392.350000 49.500000 393.650000 ;
      RECT 15.500000 392.350000 16.500000 393.650000 ;
      RECT 0.000000 392.350000 2.500000 395.650000 ;
      RECT 1169.500000 391.650000 1186.000000 392.350000 ;
      RECT 1116.500000 391.650000 1156.500000 392.350000 ;
      RECT 1066.500000 391.650000 1108.500000 392.350000 ;
      RECT 1016.500000 391.650000 1058.500000 392.350000 ;
      RECT 966.500000 391.650000 1008.500000 392.350000 ;
      RECT 916.500000 391.650000 958.500000 392.350000 ;
      RECT 866.500000 391.650000 908.500000 392.350000 ;
      RECT 816.500000 391.650000 858.500000 392.350000 ;
      RECT 766.500000 391.650000 808.500000 392.350000 ;
      RECT 716.500000 391.650000 758.500000 392.350000 ;
      RECT 666.500000 391.650000 708.500000 392.350000 ;
      RECT 616.500000 391.650000 658.500000 392.350000 ;
      RECT 566.500000 391.650000 608.500000 392.350000 ;
      RECT 516.500000 391.650000 558.500000 392.350000 ;
      RECT 466.500000 391.650000 508.500000 392.350000 ;
      RECT 416.500000 391.650000 458.500000 392.350000 ;
      RECT 366.500000 391.650000 408.500000 392.350000 ;
      RECT 316.500000 391.650000 358.500000 392.350000 ;
      RECT 266.500000 391.650000 308.500000 392.350000 ;
      RECT 216.500000 391.650000 258.500000 392.350000 ;
      RECT 166.500000 391.650000 208.500000 392.350000 ;
      RECT 116.500000 391.650000 158.500000 392.350000 ;
      RECT 66.500000 391.650000 108.500000 392.350000 ;
      RECT 29.500000 391.650000 58.500000 392.350000 ;
      RECT 0.000000 391.650000 16.500000 392.350000 ;
      RECT 1169.500000 390.350000 1170.500000 391.650000 ;
      RECT 1116.500000 390.350000 1149.500000 391.650000 ;
      RECT 1107.500000 390.350000 1108.500000 391.650000 ;
      RECT 1066.500000 390.350000 1099.500000 391.650000 ;
      RECT 1057.500000 390.350000 1058.500000 391.650000 ;
      RECT 1016.500000 390.350000 1049.500000 391.650000 ;
      RECT 1007.500000 390.350000 1008.500000 391.650000 ;
      RECT 966.500000 390.350000 999.500000 391.650000 ;
      RECT 957.500000 390.350000 958.500000 391.650000 ;
      RECT 916.500000 390.350000 949.500000 391.650000 ;
      RECT 907.500000 390.350000 908.500000 391.650000 ;
      RECT 866.500000 390.350000 899.500000 391.650000 ;
      RECT 857.500000 390.350000 858.500000 391.650000 ;
      RECT 816.500000 390.350000 849.500000 391.650000 ;
      RECT 807.500000 390.350000 808.500000 391.650000 ;
      RECT 766.500000 390.350000 799.500000 391.650000 ;
      RECT 757.500000 390.350000 758.500000 391.650000 ;
      RECT 716.500000 390.350000 749.500000 391.650000 ;
      RECT 707.500000 390.350000 708.500000 391.650000 ;
      RECT 666.500000 390.350000 699.500000 391.650000 ;
      RECT 657.500000 390.350000 658.500000 391.650000 ;
      RECT 616.500000 390.350000 649.500000 391.650000 ;
      RECT 607.500000 390.350000 608.500000 391.650000 ;
      RECT 566.500000 390.350000 599.500000 391.650000 ;
      RECT 557.500000 390.350000 558.500000 391.650000 ;
      RECT 516.500000 390.350000 549.500000 391.650000 ;
      RECT 507.500000 390.350000 508.500000 391.650000 ;
      RECT 466.500000 390.350000 499.500000 391.650000 ;
      RECT 457.500000 390.350000 458.500000 391.650000 ;
      RECT 416.500000 390.350000 449.500000 391.650000 ;
      RECT 407.500000 390.350000 408.500000 391.650000 ;
      RECT 366.500000 390.350000 399.500000 391.650000 ;
      RECT 357.500000 390.350000 358.500000 391.650000 ;
      RECT 316.500000 390.350000 349.500000 391.650000 ;
      RECT 307.500000 390.350000 308.500000 391.650000 ;
      RECT 266.500000 390.350000 299.500000 391.650000 ;
      RECT 257.500000 390.350000 258.500000 391.650000 ;
      RECT 216.500000 390.350000 249.500000 391.650000 ;
      RECT 207.500000 390.350000 208.500000 391.650000 ;
      RECT 166.500000 390.350000 199.500000 391.650000 ;
      RECT 157.500000 390.350000 158.500000 391.650000 ;
      RECT 116.500000 390.350000 149.500000 391.650000 ;
      RECT 107.500000 390.350000 108.500000 391.650000 ;
      RECT 66.500000 390.350000 99.500000 391.650000 ;
      RECT 57.500000 390.350000 58.500000 391.650000 ;
      RECT 29.500000 390.350000 49.500000 391.650000 ;
      RECT 15.500000 390.350000 16.500000 391.650000 ;
      RECT 1157.500000 389.650000 1170.500000 390.350000 ;
      RECT 1107.500000 389.650000 1149.500000 390.350000 ;
      RECT 1057.500000 389.650000 1099.500000 390.350000 ;
      RECT 1007.500000 389.650000 1049.500000 390.350000 ;
      RECT 957.500000 389.650000 999.500000 390.350000 ;
      RECT 907.500000 389.650000 949.500000 390.350000 ;
      RECT 857.500000 389.650000 899.500000 390.350000 ;
      RECT 807.500000 389.650000 849.500000 390.350000 ;
      RECT 757.500000 389.650000 799.500000 390.350000 ;
      RECT 707.500000 389.650000 749.500000 390.350000 ;
      RECT 657.500000 389.650000 699.500000 390.350000 ;
      RECT 607.500000 389.650000 649.500000 390.350000 ;
      RECT 557.500000 389.650000 599.500000 390.350000 ;
      RECT 507.500000 389.650000 549.500000 390.350000 ;
      RECT 457.500000 389.650000 499.500000 390.350000 ;
      RECT 407.500000 389.650000 449.500000 390.350000 ;
      RECT 357.500000 389.650000 399.500000 390.350000 ;
      RECT 307.500000 389.650000 349.500000 390.350000 ;
      RECT 257.500000 389.650000 299.500000 390.350000 ;
      RECT 207.500000 389.650000 249.500000 390.350000 ;
      RECT 157.500000 389.650000 199.500000 390.350000 ;
      RECT 107.500000 389.650000 149.500000 390.350000 ;
      RECT 57.500000 389.650000 99.500000 390.350000 ;
      RECT 15.500000 389.650000 49.500000 390.350000 ;
      RECT 1183.500000 388.350000 1186.000000 391.650000 ;
      RECT 1169.500000 388.350000 1170.500000 389.650000 ;
      RECT 1116.500000 388.350000 1149.500000 389.650000 ;
      RECT 1107.500000 388.350000 1108.500000 389.650000 ;
      RECT 1066.500000 388.350000 1099.500000 389.650000 ;
      RECT 1057.500000 388.350000 1058.500000 389.650000 ;
      RECT 1016.500000 388.350000 1049.500000 389.650000 ;
      RECT 1007.500000 388.350000 1008.500000 389.650000 ;
      RECT 966.500000 388.350000 999.500000 389.650000 ;
      RECT 957.500000 388.350000 958.500000 389.650000 ;
      RECT 916.500000 388.350000 949.500000 389.650000 ;
      RECT 907.500000 388.350000 908.500000 389.650000 ;
      RECT 866.500000 388.350000 899.500000 389.650000 ;
      RECT 857.500000 388.350000 858.500000 389.650000 ;
      RECT 816.500000 388.350000 849.500000 389.650000 ;
      RECT 807.500000 388.350000 808.500000 389.650000 ;
      RECT 766.500000 388.350000 799.500000 389.650000 ;
      RECT 757.500000 388.350000 758.500000 389.650000 ;
      RECT 716.500000 388.350000 749.500000 389.650000 ;
      RECT 707.500000 388.350000 708.500000 389.650000 ;
      RECT 666.500000 388.350000 699.500000 389.650000 ;
      RECT 657.500000 388.350000 658.500000 389.650000 ;
      RECT 616.500000 388.350000 649.500000 389.650000 ;
      RECT 607.500000 388.350000 608.500000 389.650000 ;
      RECT 566.500000 388.350000 599.500000 389.650000 ;
      RECT 557.500000 388.350000 558.500000 389.650000 ;
      RECT 516.500000 388.350000 549.500000 389.650000 ;
      RECT 507.500000 388.350000 508.500000 389.650000 ;
      RECT 466.500000 388.350000 499.500000 389.650000 ;
      RECT 457.500000 388.350000 458.500000 389.650000 ;
      RECT 416.500000 388.350000 449.500000 389.650000 ;
      RECT 407.500000 388.350000 408.500000 389.650000 ;
      RECT 366.500000 388.350000 399.500000 389.650000 ;
      RECT 357.500000 388.350000 358.500000 389.650000 ;
      RECT 316.500000 388.350000 349.500000 389.650000 ;
      RECT 307.500000 388.350000 308.500000 389.650000 ;
      RECT 266.500000 388.350000 299.500000 389.650000 ;
      RECT 257.500000 388.350000 258.500000 389.650000 ;
      RECT 216.500000 388.350000 249.500000 389.650000 ;
      RECT 207.500000 388.350000 208.500000 389.650000 ;
      RECT 166.500000 388.350000 199.500000 389.650000 ;
      RECT 157.500000 388.350000 158.500000 389.650000 ;
      RECT 116.500000 388.350000 149.500000 389.650000 ;
      RECT 107.500000 388.350000 108.500000 389.650000 ;
      RECT 66.500000 388.350000 99.500000 389.650000 ;
      RECT 57.500000 388.350000 58.500000 389.650000 ;
      RECT 29.500000 388.350000 49.500000 389.650000 ;
      RECT 15.500000 388.350000 16.500000 389.650000 ;
      RECT 0.000000 388.350000 2.500000 391.650000 ;
      RECT 1169.500000 387.650000 1186.000000 388.350000 ;
      RECT 1116.500000 387.650000 1156.500000 388.350000 ;
      RECT 1066.500000 387.650000 1108.500000 388.350000 ;
      RECT 1016.500000 387.650000 1058.500000 388.350000 ;
      RECT 966.500000 387.650000 1008.500000 388.350000 ;
      RECT 916.500000 387.650000 958.500000 388.350000 ;
      RECT 866.500000 387.650000 908.500000 388.350000 ;
      RECT 816.500000 387.650000 858.500000 388.350000 ;
      RECT 766.500000 387.650000 808.500000 388.350000 ;
      RECT 716.500000 387.650000 758.500000 388.350000 ;
      RECT 666.500000 387.650000 708.500000 388.350000 ;
      RECT 616.500000 387.650000 658.500000 388.350000 ;
      RECT 566.500000 387.650000 608.500000 388.350000 ;
      RECT 516.500000 387.650000 558.500000 388.350000 ;
      RECT 466.500000 387.650000 508.500000 388.350000 ;
      RECT 416.500000 387.650000 458.500000 388.350000 ;
      RECT 366.500000 387.650000 408.500000 388.350000 ;
      RECT 316.500000 387.650000 358.500000 388.350000 ;
      RECT 266.500000 387.650000 308.500000 388.350000 ;
      RECT 216.500000 387.650000 258.500000 388.350000 ;
      RECT 166.500000 387.650000 208.500000 388.350000 ;
      RECT 116.500000 387.650000 158.500000 388.350000 ;
      RECT 66.500000 387.650000 108.500000 388.350000 ;
      RECT 29.500000 387.650000 58.500000 388.350000 ;
      RECT 0.000000 387.650000 16.500000 388.350000 ;
      RECT 1169.500000 386.350000 1170.500000 387.650000 ;
      RECT 1116.500000 386.350000 1149.500000 387.650000 ;
      RECT 1107.500000 386.350000 1108.500000 387.650000 ;
      RECT 1066.500000 386.350000 1099.500000 387.650000 ;
      RECT 1057.500000 386.350000 1058.500000 387.650000 ;
      RECT 1016.500000 386.350000 1049.500000 387.650000 ;
      RECT 1007.500000 386.350000 1008.500000 387.650000 ;
      RECT 966.500000 386.350000 999.500000 387.650000 ;
      RECT 957.500000 386.350000 958.500000 387.650000 ;
      RECT 916.500000 386.350000 949.500000 387.650000 ;
      RECT 907.500000 386.350000 908.500000 387.650000 ;
      RECT 866.500000 386.350000 899.500000 387.650000 ;
      RECT 857.500000 386.350000 858.500000 387.650000 ;
      RECT 816.500000 386.350000 849.500000 387.650000 ;
      RECT 807.500000 386.350000 808.500000 387.650000 ;
      RECT 766.500000 386.350000 799.500000 387.650000 ;
      RECT 757.500000 386.350000 758.500000 387.650000 ;
      RECT 716.500000 386.350000 749.500000 387.650000 ;
      RECT 707.500000 386.350000 708.500000 387.650000 ;
      RECT 666.500000 386.350000 699.500000 387.650000 ;
      RECT 657.500000 386.350000 658.500000 387.650000 ;
      RECT 616.500000 386.350000 649.500000 387.650000 ;
      RECT 607.500000 386.350000 608.500000 387.650000 ;
      RECT 566.500000 386.350000 599.500000 387.650000 ;
      RECT 557.500000 386.350000 558.500000 387.650000 ;
      RECT 516.500000 386.350000 549.500000 387.650000 ;
      RECT 507.500000 386.350000 508.500000 387.650000 ;
      RECT 466.500000 386.350000 499.500000 387.650000 ;
      RECT 457.500000 386.350000 458.500000 387.650000 ;
      RECT 416.500000 386.350000 449.500000 387.650000 ;
      RECT 407.500000 386.350000 408.500000 387.650000 ;
      RECT 366.500000 386.350000 399.500000 387.650000 ;
      RECT 357.500000 386.350000 358.500000 387.650000 ;
      RECT 316.500000 386.350000 349.500000 387.650000 ;
      RECT 307.500000 386.350000 308.500000 387.650000 ;
      RECT 266.500000 386.350000 299.500000 387.650000 ;
      RECT 257.500000 386.350000 258.500000 387.650000 ;
      RECT 216.500000 386.350000 249.500000 387.650000 ;
      RECT 207.500000 386.350000 208.500000 387.650000 ;
      RECT 166.500000 386.350000 199.500000 387.650000 ;
      RECT 157.500000 386.350000 158.500000 387.650000 ;
      RECT 116.500000 386.350000 149.500000 387.650000 ;
      RECT 107.500000 386.350000 108.500000 387.650000 ;
      RECT 66.500000 386.350000 99.500000 387.650000 ;
      RECT 57.500000 386.350000 58.500000 387.650000 ;
      RECT 29.500000 386.350000 49.500000 387.650000 ;
      RECT 15.500000 386.350000 16.500000 387.650000 ;
      RECT 1157.500000 385.650000 1170.500000 386.350000 ;
      RECT 1107.500000 385.650000 1149.500000 386.350000 ;
      RECT 1057.500000 385.650000 1099.500000 386.350000 ;
      RECT 1007.500000 385.650000 1049.500000 386.350000 ;
      RECT 957.500000 385.650000 999.500000 386.350000 ;
      RECT 907.500000 385.650000 949.500000 386.350000 ;
      RECT 857.500000 385.650000 899.500000 386.350000 ;
      RECT 807.500000 385.650000 849.500000 386.350000 ;
      RECT 757.500000 385.650000 799.500000 386.350000 ;
      RECT 707.500000 385.650000 749.500000 386.350000 ;
      RECT 657.500000 385.650000 699.500000 386.350000 ;
      RECT 607.500000 385.650000 649.500000 386.350000 ;
      RECT 557.500000 385.650000 599.500000 386.350000 ;
      RECT 507.500000 385.650000 549.500000 386.350000 ;
      RECT 457.500000 385.650000 499.500000 386.350000 ;
      RECT 407.500000 385.650000 449.500000 386.350000 ;
      RECT 357.500000 385.650000 399.500000 386.350000 ;
      RECT 307.500000 385.650000 349.500000 386.350000 ;
      RECT 257.500000 385.650000 299.500000 386.350000 ;
      RECT 207.500000 385.650000 249.500000 386.350000 ;
      RECT 157.500000 385.650000 199.500000 386.350000 ;
      RECT 107.500000 385.650000 149.500000 386.350000 ;
      RECT 57.500000 385.650000 99.500000 386.350000 ;
      RECT 15.500000 385.650000 49.500000 386.350000 ;
      RECT 1183.500000 384.350000 1186.000000 387.650000 ;
      RECT 1169.500000 384.350000 1170.500000 385.650000 ;
      RECT 1116.500000 384.350000 1149.500000 385.650000 ;
      RECT 1107.500000 384.350000 1108.500000 385.650000 ;
      RECT 1066.500000 384.350000 1099.500000 385.650000 ;
      RECT 1057.500000 384.350000 1058.500000 385.650000 ;
      RECT 1016.500000 384.350000 1049.500000 385.650000 ;
      RECT 1007.500000 384.350000 1008.500000 385.650000 ;
      RECT 966.500000 384.350000 999.500000 385.650000 ;
      RECT 957.500000 384.350000 958.500000 385.650000 ;
      RECT 916.500000 384.350000 949.500000 385.650000 ;
      RECT 907.500000 384.350000 908.500000 385.650000 ;
      RECT 866.500000 384.350000 899.500000 385.650000 ;
      RECT 857.500000 384.350000 858.500000 385.650000 ;
      RECT 816.500000 384.350000 849.500000 385.650000 ;
      RECT 807.500000 384.350000 808.500000 385.650000 ;
      RECT 766.500000 384.350000 799.500000 385.650000 ;
      RECT 757.500000 384.350000 758.500000 385.650000 ;
      RECT 716.500000 384.350000 749.500000 385.650000 ;
      RECT 707.500000 384.350000 708.500000 385.650000 ;
      RECT 666.500000 384.350000 699.500000 385.650000 ;
      RECT 657.500000 384.350000 658.500000 385.650000 ;
      RECT 616.500000 384.350000 649.500000 385.650000 ;
      RECT 607.500000 384.350000 608.500000 385.650000 ;
      RECT 566.500000 384.350000 599.500000 385.650000 ;
      RECT 557.500000 384.350000 558.500000 385.650000 ;
      RECT 516.500000 384.350000 549.500000 385.650000 ;
      RECT 507.500000 384.350000 508.500000 385.650000 ;
      RECT 466.500000 384.350000 499.500000 385.650000 ;
      RECT 457.500000 384.350000 458.500000 385.650000 ;
      RECT 416.500000 384.350000 449.500000 385.650000 ;
      RECT 407.500000 384.350000 408.500000 385.650000 ;
      RECT 366.500000 384.350000 399.500000 385.650000 ;
      RECT 357.500000 384.350000 358.500000 385.650000 ;
      RECT 316.500000 384.350000 349.500000 385.650000 ;
      RECT 307.500000 384.350000 308.500000 385.650000 ;
      RECT 266.500000 384.350000 299.500000 385.650000 ;
      RECT 257.500000 384.350000 258.500000 385.650000 ;
      RECT 216.500000 384.350000 249.500000 385.650000 ;
      RECT 207.500000 384.350000 208.500000 385.650000 ;
      RECT 166.500000 384.350000 199.500000 385.650000 ;
      RECT 157.500000 384.350000 158.500000 385.650000 ;
      RECT 116.500000 384.350000 149.500000 385.650000 ;
      RECT 107.500000 384.350000 108.500000 385.650000 ;
      RECT 66.500000 384.350000 99.500000 385.650000 ;
      RECT 57.500000 384.350000 58.500000 385.650000 ;
      RECT 29.500000 384.350000 49.500000 385.650000 ;
      RECT 15.500000 384.350000 16.500000 385.650000 ;
      RECT 0.000000 384.350000 2.500000 387.650000 ;
      RECT 1169.500000 383.650000 1186.000000 384.350000 ;
      RECT 1116.500000 383.650000 1156.500000 384.350000 ;
      RECT 1066.500000 383.650000 1108.500000 384.350000 ;
      RECT 1016.500000 383.650000 1058.500000 384.350000 ;
      RECT 966.500000 383.650000 1008.500000 384.350000 ;
      RECT 916.500000 383.650000 958.500000 384.350000 ;
      RECT 866.500000 383.650000 908.500000 384.350000 ;
      RECT 816.500000 383.650000 858.500000 384.350000 ;
      RECT 766.500000 383.650000 808.500000 384.350000 ;
      RECT 716.500000 383.650000 758.500000 384.350000 ;
      RECT 666.500000 383.650000 708.500000 384.350000 ;
      RECT 616.500000 383.650000 658.500000 384.350000 ;
      RECT 566.500000 383.650000 608.500000 384.350000 ;
      RECT 516.500000 383.650000 558.500000 384.350000 ;
      RECT 466.500000 383.650000 508.500000 384.350000 ;
      RECT 416.500000 383.650000 458.500000 384.350000 ;
      RECT 366.500000 383.650000 408.500000 384.350000 ;
      RECT 316.500000 383.650000 358.500000 384.350000 ;
      RECT 266.500000 383.650000 308.500000 384.350000 ;
      RECT 216.500000 383.650000 258.500000 384.350000 ;
      RECT 166.500000 383.650000 208.500000 384.350000 ;
      RECT 116.500000 383.650000 158.500000 384.350000 ;
      RECT 66.500000 383.650000 108.500000 384.350000 ;
      RECT 29.500000 383.650000 58.500000 384.350000 ;
      RECT 0.000000 383.650000 16.500000 384.350000 ;
      RECT 1169.500000 382.350000 1170.500000 383.650000 ;
      RECT 1116.500000 382.350000 1149.500000 383.650000 ;
      RECT 1107.500000 382.350000 1108.500000 383.650000 ;
      RECT 1066.500000 382.350000 1099.500000 383.650000 ;
      RECT 1057.500000 382.350000 1058.500000 383.650000 ;
      RECT 1016.500000 382.350000 1049.500000 383.650000 ;
      RECT 1007.500000 382.350000 1008.500000 383.650000 ;
      RECT 966.500000 382.350000 999.500000 383.650000 ;
      RECT 957.500000 382.350000 958.500000 383.650000 ;
      RECT 916.500000 382.350000 949.500000 383.650000 ;
      RECT 907.500000 382.350000 908.500000 383.650000 ;
      RECT 866.500000 382.350000 899.500000 383.650000 ;
      RECT 857.500000 382.350000 858.500000 383.650000 ;
      RECT 816.500000 382.350000 849.500000 383.650000 ;
      RECT 807.500000 382.350000 808.500000 383.650000 ;
      RECT 766.500000 382.350000 799.500000 383.650000 ;
      RECT 757.500000 382.350000 758.500000 383.650000 ;
      RECT 716.500000 382.350000 749.500000 383.650000 ;
      RECT 707.500000 382.350000 708.500000 383.650000 ;
      RECT 666.500000 382.350000 699.500000 383.650000 ;
      RECT 657.500000 382.350000 658.500000 383.650000 ;
      RECT 616.500000 382.350000 649.500000 383.650000 ;
      RECT 607.500000 382.350000 608.500000 383.650000 ;
      RECT 566.500000 382.350000 599.500000 383.650000 ;
      RECT 557.500000 382.350000 558.500000 383.650000 ;
      RECT 516.500000 382.350000 549.500000 383.650000 ;
      RECT 507.500000 382.350000 508.500000 383.650000 ;
      RECT 466.500000 382.350000 499.500000 383.650000 ;
      RECT 457.500000 382.350000 458.500000 383.650000 ;
      RECT 416.500000 382.350000 449.500000 383.650000 ;
      RECT 407.500000 382.350000 408.500000 383.650000 ;
      RECT 366.500000 382.350000 399.500000 383.650000 ;
      RECT 357.500000 382.350000 358.500000 383.650000 ;
      RECT 316.500000 382.350000 349.500000 383.650000 ;
      RECT 307.500000 382.350000 308.500000 383.650000 ;
      RECT 266.500000 382.350000 299.500000 383.650000 ;
      RECT 257.500000 382.350000 258.500000 383.650000 ;
      RECT 216.500000 382.350000 249.500000 383.650000 ;
      RECT 207.500000 382.350000 208.500000 383.650000 ;
      RECT 166.500000 382.350000 199.500000 383.650000 ;
      RECT 157.500000 382.350000 158.500000 383.650000 ;
      RECT 116.500000 382.350000 149.500000 383.650000 ;
      RECT 107.500000 382.350000 108.500000 383.650000 ;
      RECT 66.500000 382.350000 99.500000 383.650000 ;
      RECT 57.500000 382.350000 58.500000 383.650000 ;
      RECT 29.500000 382.350000 49.500000 383.650000 ;
      RECT 15.500000 382.350000 16.500000 383.650000 ;
      RECT 1157.500000 381.650000 1170.500000 382.350000 ;
      RECT 1107.500000 381.650000 1149.500000 382.350000 ;
      RECT 1057.500000 381.650000 1099.500000 382.350000 ;
      RECT 1007.500000 381.650000 1049.500000 382.350000 ;
      RECT 957.500000 381.650000 999.500000 382.350000 ;
      RECT 907.500000 381.650000 949.500000 382.350000 ;
      RECT 857.500000 381.650000 899.500000 382.350000 ;
      RECT 807.500000 381.650000 849.500000 382.350000 ;
      RECT 757.500000 381.650000 799.500000 382.350000 ;
      RECT 707.500000 381.650000 749.500000 382.350000 ;
      RECT 657.500000 381.650000 699.500000 382.350000 ;
      RECT 607.500000 381.650000 649.500000 382.350000 ;
      RECT 557.500000 381.650000 599.500000 382.350000 ;
      RECT 507.500000 381.650000 549.500000 382.350000 ;
      RECT 457.500000 381.650000 499.500000 382.350000 ;
      RECT 407.500000 381.650000 449.500000 382.350000 ;
      RECT 357.500000 381.650000 399.500000 382.350000 ;
      RECT 307.500000 381.650000 349.500000 382.350000 ;
      RECT 257.500000 381.650000 299.500000 382.350000 ;
      RECT 207.500000 381.650000 249.500000 382.350000 ;
      RECT 157.500000 381.650000 199.500000 382.350000 ;
      RECT 107.500000 381.650000 149.500000 382.350000 ;
      RECT 57.500000 381.650000 99.500000 382.350000 ;
      RECT 15.500000 381.650000 49.500000 382.350000 ;
      RECT 1183.500000 380.350000 1186.000000 383.650000 ;
      RECT 1169.500000 380.350000 1170.500000 381.650000 ;
      RECT 1116.500000 380.350000 1149.500000 381.650000 ;
      RECT 1107.500000 380.350000 1108.500000 381.650000 ;
      RECT 1066.500000 380.350000 1099.500000 381.650000 ;
      RECT 1057.500000 380.350000 1058.500000 381.650000 ;
      RECT 1016.500000 380.350000 1049.500000 381.650000 ;
      RECT 1007.500000 380.350000 1008.500000 381.650000 ;
      RECT 966.500000 380.350000 999.500000 381.650000 ;
      RECT 957.500000 380.350000 958.500000 381.650000 ;
      RECT 916.500000 380.350000 949.500000 381.650000 ;
      RECT 907.500000 380.350000 908.500000 381.650000 ;
      RECT 866.500000 380.350000 899.500000 381.650000 ;
      RECT 857.500000 380.350000 858.500000 381.650000 ;
      RECT 816.500000 380.350000 849.500000 381.650000 ;
      RECT 807.500000 380.350000 808.500000 381.650000 ;
      RECT 766.500000 380.350000 799.500000 381.650000 ;
      RECT 757.500000 380.350000 758.500000 381.650000 ;
      RECT 716.500000 380.350000 749.500000 381.650000 ;
      RECT 707.500000 380.350000 708.500000 381.650000 ;
      RECT 666.500000 380.350000 699.500000 381.650000 ;
      RECT 657.500000 380.350000 658.500000 381.650000 ;
      RECT 616.500000 380.350000 649.500000 381.650000 ;
      RECT 607.500000 380.350000 608.500000 381.650000 ;
      RECT 566.500000 380.350000 599.500000 381.650000 ;
      RECT 557.500000 380.350000 558.500000 381.650000 ;
      RECT 516.500000 380.350000 549.500000 381.650000 ;
      RECT 507.500000 380.350000 508.500000 381.650000 ;
      RECT 466.500000 380.350000 499.500000 381.650000 ;
      RECT 457.500000 380.350000 458.500000 381.650000 ;
      RECT 416.500000 380.350000 449.500000 381.650000 ;
      RECT 407.500000 380.350000 408.500000 381.650000 ;
      RECT 366.500000 380.350000 399.500000 381.650000 ;
      RECT 357.500000 380.350000 358.500000 381.650000 ;
      RECT 316.500000 380.350000 349.500000 381.650000 ;
      RECT 307.500000 380.350000 308.500000 381.650000 ;
      RECT 266.500000 380.350000 299.500000 381.650000 ;
      RECT 257.500000 380.350000 258.500000 381.650000 ;
      RECT 216.500000 380.350000 249.500000 381.650000 ;
      RECT 207.500000 380.350000 208.500000 381.650000 ;
      RECT 166.500000 380.350000 199.500000 381.650000 ;
      RECT 157.500000 380.350000 158.500000 381.650000 ;
      RECT 116.500000 380.350000 149.500000 381.650000 ;
      RECT 107.500000 380.350000 108.500000 381.650000 ;
      RECT 66.500000 380.350000 99.500000 381.650000 ;
      RECT 57.500000 380.350000 58.500000 381.650000 ;
      RECT 29.500000 380.350000 49.500000 381.650000 ;
      RECT 15.500000 380.350000 16.500000 381.650000 ;
      RECT 0.000000 380.350000 2.500000 383.650000 ;
      RECT 1169.500000 379.650000 1186.000000 380.350000 ;
      RECT 1116.500000 379.650000 1156.500000 380.350000 ;
      RECT 1066.500000 379.650000 1108.500000 380.350000 ;
      RECT 1016.500000 379.650000 1058.500000 380.350000 ;
      RECT 966.500000 379.650000 1008.500000 380.350000 ;
      RECT 916.500000 379.650000 958.500000 380.350000 ;
      RECT 866.500000 379.650000 908.500000 380.350000 ;
      RECT 816.500000 379.650000 858.500000 380.350000 ;
      RECT 766.500000 379.650000 808.500000 380.350000 ;
      RECT 716.500000 379.650000 758.500000 380.350000 ;
      RECT 666.500000 379.650000 708.500000 380.350000 ;
      RECT 616.500000 379.650000 658.500000 380.350000 ;
      RECT 566.500000 379.650000 608.500000 380.350000 ;
      RECT 516.500000 379.650000 558.500000 380.350000 ;
      RECT 466.500000 379.650000 508.500000 380.350000 ;
      RECT 416.500000 379.650000 458.500000 380.350000 ;
      RECT 366.500000 379.650000 408.500000 380.350000 ;
      RECT 316.500000 379.650000 358.500000 380.350000 ;
      RECT 266.500000 379.650000 308.500000 380.350000 ;
      RECT 216.500000 379.650000 258.500000 380.350000 ;
      RECT 166.500000 379.650000 208.500000 380.350000 ;
      RECT 116.500000 379.650000 158.500000 380.350000 ;
      RECT 66.500000 379.650000 108.500000 380.350000 ;
      RECT 29.500000 379.650000 58.500000 380.350000 ;
      RECT 0.000000 379.650000 16.500000 380.350000 ;
      RECT 1169.500000 378.350000 1170.500000 379.650000 ;
      RECT 1116.500000 378.350000 1149.500000 379.650000 ;
      RECT 1107.500000 378.350000 1108.500000 379.650000 ;
      RECT 1066.500000 378.350000 1099.500000 379.650000 ;
      RECT 1057.500000 378.350000 1058.500000 379.650000 ;
      RECT 1016.500000 378.350000 1049.500000 379.650000 ;
      RECT 1007.500000 378.350000 1008.500000 379.650000 ;
      RECT 966.500000 378.350000 999.500000 379.650000 ;
      RECT 957.500000 378.350000 958.500000 379.650000 ;
      RECT 916.500000 378.350000 949.500000 379.650000 ;
      RECT 907.500000 378.350000 908.500000 379.650000 ;
      RECT 866.500000 378.350000 899.500000 379.650000 ;
      RECT 857.500000 378.350000 858.500000 379.650000 ;
      RECT 816.500000 378.350000 849.500000 379.650000 ;
      RECT 807.500000 378.350000 808.500000 379.650000 ;
      RECT 766.500000 378.350000 799.500000 379.650000 ;
      RECT 757.500000 378.350000 758.500000 379.650000 ;
      RECT 716.500000 378.350000 749.500000 379.650000 ;
      RECT 707.500000 378.350000 708.500000 379.650000 ;
      RECT 666.500000 378.350000 699.500000 379.650000 ;
      RECT 657.500000 378.350000 658.500000 379.650000 ;
      RECT 616.500000 378.350000 649.500000 379.650000 ;
      RECT 607.500000 378.350000 608.500000 379.650000 ;
      RECT 566.500000 378.350000 599.500000 379.650000 ;
      RECT 557.500000 378.350000 558.500000 379.650000 ;
      RECT 516.500000 378.350000 549.500000 379.650000 ;
      RECT 507.500000 378.350000 508.500000 379.650000 ;
      RECT 466.500000 378.350000 499.500000 379.650000 ;
      RECT 457.500000 378.350000 458.500000 379.650000 ;
      RECT 416.500000 378.350000 449.500000 379.650000 ;
      RECT 407.500000 378.350000 408.500000 379.650000 ;
      RECT 366.500000 378.350000 399.500000 379.650000 ;
      RECT 357.500000 378.350000 358.500000 379.650000 ;
      RECT 316.500000 378.350000 349.500000 379.650000 ;
      RECT 307.500000 378.350000 308.500000 379.650000 ;
      RECT 266.500000 378.350000 299.500000 379.650000 ;
      RECT 257.500000 378.350000 258.500000 379.650000 ;
      RECT 216.500000 378.350000 249.500000 379.650000 ;
      RECT 207.500000 378.350000 208.500000 379.650000 ;
      RECT 166.500000 378.350000 199.500000 379.650000 ;
      RECT 157.500000 378.350000 158.500000 379.650000 ;
      RECT 116.500000 378.350000 149.500000 379.650000 ;
      RECT 107.500000 378.350000 108.500000 379.650000 ;
      RECT 66.500000 378.350000 99.500000 379.650000 ;
      RECT 57.500000 378.350000 58.500000 379.650000 ;
      RECT 29.500000 378.350000 49.500000 379.650000 ;
      RECT 15.500000 378.350000 16.500000 379.650000 ;
      RECT 1157.500000 377.650000 1170.500000 378.350000 ;
      RECT 1107.500000 377.650000 1149.500000 378.350000 ;
      RECT 1057.500000 377.650000 1099.500000 378.350000 ;
      RECT 1007.500000 377.650000 1049.500000 378.350000 ;
      RECT 957.500000 377.650000 999.500000 378.350000 ;
      RECT 907.500000 377.650000 949.500000 378.350000 ;
      RECT 857.500000 377.650000 899.500000 378.350000 ;
      RECT 807.500000 377.650000 849.500000 378.350000 ;
      RECT 757.500000 377.650000 799.500000 378.350000 ;
      RECT 707.500000 377.650000 749.500000 378.350000 ;
      RECT 657.500000 377.650000 699.500000 378.350000 ;
      RECT 607.500000 377.650000 649.500000 378.350000 ;
      RECT 557.500000 377.650000 599.500000 378.350000 ;
      RECT 507.500000 377.650000 549.500000 378.350000 ;
      RECT 457.500000 377.650000 499.500000 378.350000 ;
      RECT 407.500000 377.650000 449.500000 378.350000 ;
      RECT 357.500000 377.650000 399.500000 378.350000 ;
      RECT 307.500000 377.650000 349.500000 378.350000 ;
      RECT 257.500000 377.650000 299.500000 378.350000 ;
      RECT 207.500000 377.650000 249.500000 378.350000 ;
      RECT 157.500000 377.650000 199.500000 378.350000 ;
      RECT 107.500000 377.650000 149.500000 378.350000 ;
      RECT 57.500000 377.650000 99.500000 378.350000 ;
      RECT 15.500000 377.650000 49.500000 378.350000 ;
      RECT 1183.500000 376.350000 1186.000000 379.650000 ;
      RECT 1169.500000 376.350000 1170.500000 377.650000 ;
      RECT 1116.500000 376.350000 1149.500000 377.650000 ;
      RECT 1107.500000 376.350000 1108.500000 377.650000 ;
      RECT 1066.500000 376.350000 1099.500000 377.650000 ;
      RECT 1057.500000 376.350000 1058.500000 377.650000 ;
      RECT 1016.500000 376.350000 1049.500000 377.650000 ;
      RECT 1007.500000 376.350000 1008.500000 377.650000 ;
      RECT 966.500000 376.350000 999.500000 377.650000 ;
      RECT 957.500000 376.350000 958.500000 377.650000 ;
      RECT 916.500000 376.350000 949.500000 377.650000 ;
      RECT 907.500000 376.350000 908.500000 377.650000 ;
      RECT 866.500000 376.350000 899.500000 377.650000 ;
      RECT 857.500000 376.350000 858.500000 377.650000 ;
      RECT 816.500000 376.350000 849.500000 377.650000 ;
      RECT 807.500000 376.350000 808.500000 377.650000 ;
      RECT 766.500000 376.350000 799.500000 377.650000 ;
      RECT 757.500000 376.350000 758.500000 377.650000 ;
      RECT 716.500000 376.350000 749.500000 377.650000 ;
      RECT 707.500000 376.350000 708.500000 377.650000 ;
      RECT 666.500000 376.350000 699.500000 377.650000 ;
      RECT 657.500000 376.350000 658.500000 377.650000 ;
      RECT 616.500000 376.350000 649.500000 377.650000 ;
      RECT 607.500000 376.350000 608.500000 377.650000 ;
      RECT 566.500000 376.350000 599.500000 377.650000 ;
      RECT 557.500000 376.350000 558.500000 377.650000 ;
      RECT 516.500000 376.350000 549.500000 377.650000 ;
      RECT 507.500000 376.350000 508.500000 377.650000 ;
      RECT 466.500000 376.350000 499.500000 377.650000 ;
      RECT 457.500000 376.350000 458.500000 377.650000 ;
      RECT 416.500000 376.350000 449.500000 377.650000 ;
      RECT 407.500000 376.350000 408.500000 377.650000 ;
      RECT 366.500000 376.350000 399.500000 377.650000 ;
      RECT 357.500000 376.350000 358.500000 377.650000 ;
      RECT 316.500000 376.350000 349.500000 377.650000 ;
      RECT 307.500000 376.350000 308.500000 377.650000 ;
      RECT 266.500000 376.350000 299.500000 377.650000 ;
      RECT 257.500000 376.350000 258.500000 377.650000 ;
      RECT 216.500000 376.350000 249.500000 377.650000 ;
      RECT 207.500000 376.350000 208.500000 377.650000 ;
      RECT 166.500000 376.350000 199.500000 377.650000 ;
      RECT 157.500000 376.350000 158.500000 377.650000 ;
      RECT 116.500000 376.350000 149.500000 377.650000 ;
      RECT 107.500000 376.350000 108.500000 377.650000 ;
      RECT 66.500000 376.350000 99.500000 377.650000 ;
      RECT 57.500000 376.350000 58.500000 377.650000 ;
      RECT 29.500000 376.350000 49.500000 377.650000 ;
      RECT 15.500000 376.350000 16.500000 377.650000 ;
      RECT 0.000000 376.350000 2.500000 379.650000 ;
      RECT 1169.500000 375.650000 1186.000000 376.350000 ;
      RECT 1116.500000 375.650000 1156.500000 376.350000 ;
      RECT 1066.500000 375.650000 1108.500000 376.350000 ;
      RECT 1016.500000 375.650000 1058.500000 376.350000 ;
      RECT 966.500000 375.650000 1008.500000 376.350000 ;
      RECT 916.500000 375.650000 958.500000 376.350000 ;
      RECT 866.500000 375.650000 908.500000 376.350000 ;
      RECT 816.500000 375.650000 858.500000 376.350000 ;
      RECT 766.500000 375.650000 808.500000 376.350000 ;
      RECT 716.500000 375.650000 758.500000 376.350000 ;
      RECT 666.500000 375.650000 708.500000 376.350000 ;
      RECT 616.500000 375.650000 658.500000 376.350000 ;
      RECT 566.500000 375.650000 608.500000 376.350000 ;
      RECT 516.500000 375.650000 558.500000 376.350000 ;
      RECT 466.500000 375.650000 508.500000 376.350000 ;
      RECT 416.500000 375.650000 458.500000 376.350000 ;
      RECT 366.500000 375.650000 408.500000 376.350000 ;
      RECT 316.500000 375.650000 358.500000 376.350000 ;
      RECT 266.500000 375.650000 308.500000 376.350000 ;
      RECT 216.500000 375.650000 258.500000 376.350000 ;
      RECT 166.500000 375.650000 208.500000 376.350000 ;
      RECT 116.500000 375.650000 158.500000 376.350000 ;
      RECT 66.500000 375.650000 108.500000 376.350000 ;
      RECT 29.500000 375.650000 58.500000 376.350000 ;
      RECT 0.000000 375.650000 16.500000 376.350000 ;
      RECT 1169.500000 374.350000 1170.500000 375.650000 ;
      RECT 1116.500000 374.350000 1149.500000 375.650000 ;
      RECT 1107.500000 374.350000 1108.500000 375.650000 ;
      RECT 1066.500000 374.350000 1099.500000 375.650000 ;
      RECT 1057.500000 374.350000 1058.500000 375.650000 ;
      RECT 1016.500000 374.350000 1049.500000 375.650000 ;
      RECT 1007.500000 374.350000 1008.500000 375.650000 ;
      RECT 966.500000 374.350000 999.500000 375.650000 ;
      RECT 957.500000 374.350000 958.500000 375.650000 ;
      RECT 916.500000 374.350000 949.500000 375.650000 ;
      RECT 907.500000 374.350000 908.500000 375.650000 ;
      RECT 866.500000 374.350000 899.500000 375.650000 ;
      RECT 857.500000 374.350000 858.500000 375.650000 ;
      RECT 816.500000 374.350000 849.500000 375.650000 ;
      RECT 807.500000 374.350000 808.500000 375.650000 ;
      RECT 766.500000 374.350000 799.500000 375.650000 ;
      RECT 757.500000 374.350000 758.500000 375.650000 ;
      RECT 716.500000 374.350000 749.500000 375.650000 ;
      RECT 707.500000 374.350000 708.500000 375.650000 ;
      RECT 666.500000 374.350000 699.500000 375.650000 ;
      RECT 657.500000 374.350000 658.500000 375.650000 ;
      RECT 616.500000 374.350000 649.500000 375.650000 ;
      RECT 607.500000 374.350000 608.500000 375.650000 ;
      RECT 566.500000 374.350000 599.500000 375.650000 ;
      RECT 557.500000 374.350000 558.500000 375.650000 ;
      RECT 516.500000 374.350000 549.500000 375.650000 ;
      RECT 507.500000 374.350000 508.500000 375.650000 ;
      RECT 466.500000 374.350000 499.500000 375.650000 ;
      RECT 457.500000 374.350000 458.500000 375.650000 ;
      RECT 416.500000 374.350000 449.500000 375.650000 ;
      RECT 407.500000 374.350000 408.500000 375.650000 ;
      RECT 366.500000 374.350000 399.500000 375.650000 ;
      RECT 357.500000 374.350000 358.500000 375.650000 ;
      RECT 316.500000 374.350000 349.500000 375.650000 ;
      RECT 307.500000 374.350000 308.500000 375.650000 ;
      RECT 266.500000 374.350000 299.500000 375.650000 ;
      RECT 257.500000 374.350000 258.500000 375.650000 ;
      RECT 216.500000 374.350000 249.500000 375.650000 ;
      RECT 207.500000 374.350000 208.500000 375.650000 ;
      RECT 166.500000 374.350000 199.500000 375.650000 ;
      RECT 157.500000 374.350000 158.500000 375.650000 ;
      RECT 116.500000 374.350000 149.500000 375.650000 ;
      RECT 107.500000 374.350000 108.500000 375.650000 ;
      RECT 66.500000 374.350000 99.500000 375.650000 ;
      RECT 57.500000 374.350000 58.500000 375.650000 ;
      RECT 29.500000 374.350000 49.500000 375.650000 ;
      RECT 15.500000 374.350000 16.500000 375.650000 ;
      RECT 1157.500000 373.650000 1170.500000 374.350000 ;
      RECT 1107.500000 373.650000 1149.500000 374.350000 ;
      RECT 1057.500000 373.650000 1099.500000 374.350000 ;
      RECT 1007.500000 373.650000 1049.500000 374.350000 ;
      RECT 957.500000 373.650000 999.500000 374.350000 ;
      RECT 907.500000 373.650000 949.500000 374.350000 ;
      RECT 857.500000 373.650000 899.500000 374.350000 ;
      RECT 807.500000 373.650000 849.500000 374.350000 ;
      RECT 757.500000 373.650000 799.500000 374.350000 ;
      RECT 707.500000 373.650000 749.500000 374.350000 ;
      RECT 657.500000 373.650000 699.500000 374.350000 ;
      RECT 607.500000 373.650000 649.500000 374.350000 ;
      RECT 557.500000 373.650000 599.500000 374.350000 ;
      RECT 507.500000 373.650000 549.500000 374.350000 ;
      RECT 457.500000 373.650000 499.500000 374.350000 ;
      RECT 407.500000 373.650000 449.500000 374.350000 ;
      RECT 357.500000 373.650000 399.500000 374.350000 ;
      RECT 307.500000 373.650000 349.500000 374.350000 ;
      RECT 257.500000 373.650000 299.500000 374.350000 ;
      RECT 207.500000 373.650000 249.500000 374.350000 ;
      RECT 157.500000 373.650000 199.500000 374.350000 ;
      RECT 107.500000 373.650000 149.500000 374.350000 ;
      RECT 57.500000 373.650000 99.500000 374.350000 ;
      RECT 15.500000 373.650000 49.500000 374.350000 ;
      RECT 1183.500000 372.350000 1186.000000 375.650000 ;
      RECT 1169.500000 372.350000 1170.500000 373.650000 ;
      RECT 1116.500000 372.350000 1149.500000 373.650000 ;
      RECT 1107.500000 372.350000 1108.500000 373.650000 ;
      RECT 1066.500000 372.350000 1099.500000 373.650000 ;
      RECT 1057.500000 372.350000 1058.500000 373.650000 ;
      RECT 1016.500000 372.350000 1049.500000 373.650000 ;
      RECT 1007.500000 372.350000 1008.500000 373.650000 ;
      RECT 966.500000 372.350000 999.500000 373.650000 ;
      RECT 957.500000 372.350000 958.500000 373.650000 ;
      RECT 916.500000 372.350000 949.500000 373.650000 ;
      RECT 907.500000 372.350000 908.500000 373.650000 ;
      RECT 866.500000 372.350000 899.500000 373.650000 ;
      RECT 857.500000 372.350000 858.500000 373.650000 ;
      RECT 816.500000 372.350000 849.500000 373.650000 ;
      RECT 807.500000 372.350000 808.500000 373.650000 ;
      RECT 766.500000 372.350000 799.500000 373.650000 ;
      RECT 757.500000 372.350000 758.500000 373.650000 ;
      RECT 716.500000 372.350000 749.500000 373.650000 ;
      RECT 707.500000 372.350000 708.500000 373.650000 ;
      RECT 666.500000 372.350000 699.500000 373.650000 ;
      RECT 657.500000 372.350000 658.500000 373.650000 ;
      RECT 616.500000 372.350000 649.500000 373.650000 ;
      RECT 607.500000 372.350000 608.500000 373.650000 ;
      RECT 566.500000 372.350000 599.500000 373.650000 ;
      RECT 557.500000 372.350000 558.500000 373.650000 ;
      RECT 516.500000 372.350000 549.500000 373.650000 ;
      RECT 507.500000 372.350000 508.500000 373.650000 ;
      RECT 466.500000 372.350000 499.500000 373.650000 ;
      RECT 457.500000 372.350000 458.500000 373.650000 ;
      RECT 416.500000 372.350000 449.500000 373.650000 ;
      RECT 407.500000 372.350000 408.500000 373.650000 ;
      RECT 366.500000 372.350000 399.500000 373.650000 ;
      RECT 357.500000 372.350000 358.500000 373.650000 ;
      RECT 316.500000 372.350000 349.500000 373.650000 ;
      RECT 307.500000 372.350000 308.500000 373.650000 ;
      RECT 266.500000 372.350000 299.500000 373.650000 ;
      RECT 257.500000 372.350000 258.500000 373.650000 ;
      RECT 216.500000 372.350000 249.500000 373.650000 ;
      RECT 207.500000 372.350000 208.500000 373.650000 ;
      RECT 166.500000 372.350000 199.500000 373.650000 ;
      RECT 157.500000 372.350000 158.500000 373.650000 ;
      RECT 116.500000 372.350000 149.500000 373.650000 ;
      RECT 107.500000 372.350000 108.500000 373.650000 ;
      RECT 66.500000 372.350000 99.500000 373.650000 ;
      RECT 57.500000 372.350000 58.500000 373.650000 ;
      RECT 29.500000 372.350000 49.500000 373.650000 ;
      RECT 15.500000 372.350000 16.500000 373.650000 ;
      RECT 0.000000 372.350000 2.500000 375.650000 ;
      RECT 1169.500000 371.650000 1186.000000 372.350000 ;
      RECT 1116.500000 371.650000 1156.500000 372.350000 ;
      RECT 1066.500000 371.650000 1108.500000 372.350000 ;
      RECT 1016.500000 371.650000 1058.500000 372.350000 ;
      RECT 966.500000 371.650000 1008.500000 372.350000 ;
      RECT 916.500000 371.650000 958.500000 372.350000 ;
      RECT 866.500000 371.650000 908.500000 372.350000 ;
      RECT 816.500000 371.650000 858.500000 372.350000 ;
      RECT 766.500000 371.650000 808.500000 372.350000 ;
      RECT 716.500000 371.650000 758.500000 372.350000 ;
      RECT 666.500000 371.650000 708.500000 372.350000 ;
      RECT 616.500000 371.650000 658.500000 372.350000 ;
      RECT 566.500000 371.650000 608.500000 372.350000 ;
      RECT 516.500000 371.650000 558.500000 372.350000 ;
      RECT 466.500000 371.650000 508.500000 372.350000 ;
      RECT 416.500000 371.650000 458.500000 372.350000 ;
      RECT 366.500000 371.650000 408.500000 372.350000 ;
      RECT 316.500000 371.650000 358.500000 372.350000 ;
      RECT 266.500000 371.650000 308.500000 372.350000 ;
      RECT 216.500000 371.650000 258.500000 372.350000 ;
      RECT 166.500000 371.650000 208.500000 372.350000 ;
      RECT 116.500000 371.650000 158.500000 372.350000 ;
      RECT 66.500000 371.650000 108.500000 372.350000 ;
      RECT 29.500000 371.650000 58.500000 372.350000 ;
      RECT 0.000000 371.650000 16.500000 372.350000 ;
      RECT 1169.500000 370.350000 1170.500000 371.650000 ;
      RECT 1116.500000 370.350000 1149.500000 371.650000 ;
      RECT 1107.500000 370.350000 1108.500000 371.650000 ;
      RECT 1066.500000 370.350000 1099.500000 371.650000 ;
      RECT 1057.500000 370.350000 1058.500000 371.650000 ;
      RECT 1016.500000 370.350000 1049.500000 371.650000 ;
      RECT 1007.500000 370.350000 1008.500000 371.650000 ;
      RECT 966.500000 370.350000 999.500000 371.650000 ;
      RECT 957.500000 370.350000 958.500000 371.650000 ;
      RECT 916.500000 370.350000 949.500000 371.650000 ;
      RECT 907.500000 370.350000 908.500000 371.650000 ;
      RECT 866.500000 370.350000 899.500000 371.650000 ;
      RECT 857.500000 370.350000 858.500000 371.650000 ;
      RECT 816.500000 370.350000 849.500000 371.650000 ;
      RECT 807.500000 370.350000 808.500000 371.650000 ;
      RECT 766.500000 370.350000 799.500000 371.650000 ;
      RECT 757.500000 370.350000 758.500000 371.650000 ;
      RECT 716.500000 370.350000 749.500000 371.650000 ;
      RECT 707.500000 370.350000 708.500000 371.650000 ;
      RECT 666.500000 370.350000 699.500000 371.650000 ;
      RECT 657.500000 370.350000 658.500000 371.650000 ;
      RECT 616.500000 370.350000 649.500000 371.650000 ;
      RECT 607.500000 370.350000 608.500000 371.650000 ;
      RECT 566.500000 370.350000 599.500000 371.650000 ;
      RECT 557.500000 370.350000 558.500000 371.650000 ;
      RECT 516.500000 370.350000 549.500000 371.650000 ;
      RECT 507.500000 370.350000 508.500000 371.650000 ;
      RECT 466.500000 370.350000 499.500000 371.650000 ;
      RECT 457.500000 370.350000 458.500000 371.650000 ;
      RECT 416.500000 370.350000 449.500000 371.650000 ;
      RECT 407.500000 370.350000 408.500000 371.650000 ;
      RECT 366.500000 370.350000 399.500000 371.650000 ;
      RECT 357.500000 370.350000 358.500000 371.650000 ;
      RECT 316.500000 370.350000 349.500000 371.650000 ;
      RECT 307.500000 370.350000 308.500000 371.650000 ;
      RECT 266.500000 370.350000 299.500000 371.650000 ;
      RECT 257.500000 370.350000 258.500000 371.650000 ;
      RECT 216.500000 370.350000 249.500000 371.650000 ;
      RECT 207.500000 370.350000 208.500000 371.650000 ;
      RECT 166.500000 370.350000 199.500000 371.650000 ;
      RECT 157.500000 370.350000 158.500000 371.650000 ;
      RECT 116.500000 370.350000 149.500000 371.650000 ;
      RECT 107.500000 370.350000 108.500000 371.650000 ;
      RECT 66.500000 370.350000 99.500000 371.650000 ;
      RECT 57.500000 370.350000 58.500000 371.650000 ;
      RECT 29.500000 370.350000 49.500000 371.650000 ;
      RECT 15.500000 370.350000 16.500000 371.650000 ;
      RECT 1157.500000 369.650000 1170.500000 370.350000 ;
      RECT 1107.500000 369.650000 1149.500000 370.350000 ;
      RECT 1057.500000 369.650000 1099.500000 370.350000 ;
      RECT 1007.500000 369.650000 1049.500000 370.350000 ;
      RECT 957.500000 369.650000 999.500000 370.350000 ;
      RECT 907.500000 369.650000 949.500000 370.350000 ;
      RECT 857.500000 369.650000 899.500000 370.350000 ;
      RECT 807.500000 369.650000 849.500000 370.350000 ;
      RECT 757.500000 369.650000 799.500000 370.350000 ;
      RECT 707.500000 369.650000 749.500000 370.350000 ;
      RECT 657.500000 369.650000 699.500000 370.350000 ;
      RECT 607.500000 369.650000 649.500000 370.350000 ;
      RECT 557.500000 369.650000 599.500000 370.350000 ;
      RECT 507.500000 369.650000 549.500000 370.350000 ;
      RECT 407.500000 369.650000 449.500000 370.350000 ;
      RECT 357.500000 369.650000 399.500000 370.350000 ;
      RECT 307.500000 369.650000 349.500000 370.350000 ;
      RECT 257.500000 369.650000 299.500000 370.350000 ;
      RECT 207.500000 369.650000 249.500000 370.350000 ;
      RECT 157.500000 369.650000 199.500000 370.350000 ;
      RECT 107.500000 369.650000 149.500000 370.350000 ;
      RECT 57.500000 369.650000 99.500000 370.350000 ;
      RECT 15.500000 369.650000 49.500000 370.350000 ;
      RECT 1183.500000 368.350000 1186.000000 371.650000 ;
      RECT 1169.500000 368.350000 1170.500000 369.650000 ;
      RECT 1116.500000 368.350000 1149.500000 369.650000 ;
      RECT 1107.500000 368.350000 1108.500000 369.650000 ;
      RECT 1066.500000 368.350000 1099.500000 369.650000 ;
      RECT 1057.500000 368.350000 1058.500000 369.650000 ;
      RECT 1016.500000 368.350000 1049.500000 369.650000 ;
      RECT 1007.500000 368.350000 1008.500000 369.650000 ;
      RECT 966.500000 368.350000 999.500000 369.650000 ;
      RECT 957.500000 368.350000 958.500000 369.650000 ;
      RECT 916.500000 368.350000 949.500000 369.650000 ;
      RECT 907.500000 368.350000 908.500000 369.650000 ;
      RECT 866.500000 368.350000 899.500000 369.650000 ;
      RECT 857.500000 368.350000 858.500000 369.650000 ;
      RECT 816.500000 368.350000 849.500000 369.650000 ;
      RECT 807.500000 368.350000 808.500000 369.650000 ;
      RECT 766.500000 368.350000 799.500000 369.650000 ;
      RECT 757.500000 368.350000 758.500000 369.650000 ;
      RECT 716.500000 368.350000 749.500000 369.650000 ;
      RECT 707.500000 368.350000 708.500000 369.650000 ;
      RECT 666.500000 368.350000 699.500000 369.650000 ;
      RECT 657.500000 368.350000 658.500000 369.650000 ;
      RECT 616.500000 368.350000 649.500000 369.650000 ;
      RECT 607.500000 368.350000 608.500000 369.650000 ;
      RECT 566.500000 368.350000 599.500000 369.650000 ;
      RECT 557.500000 368.350000 558.500000 369.650000 ;
      RECT 516.500000 368.350000 549.500000 369.650000 ;
      RECT 507.500000 368.350000 508.500000 369.650000 ;
      RECT 457.500000 368.350000 499.500000 370.350000 ;
      RECT 407.500000 368.350000 408.500000 369.650000 ;
      RECT 366.500000 368.350000 399.500000 369.650000 ;
      RECT 357.500000 368.350000 358.500000 369.650000 ;
      RECT 316.500000 368.350000 349.500000 369.650000 ;
      RECT 307.500000 368.350000 308.500000 369.650000 ;
      RECT 266.500000 368.350000 299.500000 369.650000 ;
      RECT 257.500000 368.350000 258.500000 369.650000 ;
      RECT 216.500000 368.350000 249.500000 369.650000 ;
      RECT 207.500000 368.350000 208.500000 369.650000 ;
      RECT 166.500000 368.350000 199.500000 369.650000 ;
      RECT 157.500000 368.350000 158.500000 369.650000 ;
      RECT 116.500000 368.350000 149.500000 369.650000 ;
      RECT 107.500000 368.350000 108.500000 369.650000 ;
      RECT 66.500000 368.350000 99.500000 369.650000 ;
      RECT 57.500000 368.350000 58.500000 369.650000 ;
      RECT 29.500000 368.350000 49.500000 369.650000 ;
      RECT 15.500000 368.350000 16.500000 369.650000 ;
      RECT 0.000000 368.350000 2.500000 371.650000 ;
      RECT 1169.500000 367.650000 1186.000000 368.350000 ;
      RECT 1116.500000 367.650000 1156.500000 368.350000 ;
      RECT 1066.500000 367.650000 1108.500000 368.350000 ;
      RECT 1016.500000 367.650000 1058.500000 368.350000 ;
      RECT 966.500000 367.650000 1008.500000 368.350000 ;
      RECT 916.500000 367.650000 958.500000 368.350000 ;
      RECT 866.500000 367.650000 908.500000 368.350000 ;
      RECT 816.500000 367.650000 858.500000 368.350000 ;
      RECT 766.500000 367.650000 808.500000 368.350000 ;
      RECT 716.500000 367.650000 758.500000 368.350000 ;
      RECT 666.500000 367.650000 708.500000 368.350000 ;
      RECT 616.500000 367.650000 658.500000 368.350000 ;
      RECT 566.500000 367.650000 608.500000 368.350000 ;
      RECT 516.500000 367.650000 558.500000 368.350000 ;
      RECT 457.500000 367.650000 508.500000 368.350000 ;
      RECT 366.500000 367.650000 408.500000 368.350000 ;
      RECT 316.500000 367.650000 358.500000 368.350000 ;
      RECT 266.500000 367.650000 308.500000 368.350000 ;
      RECT 216.500000 367.650000 258.500000 368.350000 ;
      RECT 166.500000 367.650000 208.500000 368.350000 ;
      RECT 116.500000 367.650000 158.500000 368.350000 ;
      RECT 66.500000 367.650000 108.500000 368.350000 ;
      RECT 29.500000 367.650000 58.500000 368.350000 ;
      RECT 0.000000 367.650000 16.500000 368.350000 ;
      RECT 1169.500000 366.350000 1170.500000 367.650000 ;
      RECT 1116.500000 366.350000 1149.500000 367.650000 ;
      RECT 1107.500000 366.350000 1108.500000 367.650000 ;
      RECT 1066.500000 366.350000 1099.500000 367.650000 ;
      RECT 1057.500000 366.350000 1058.500000 367.650000 ;
      RECT 1016.500000 366.350000 1049.500000 367.650000 ;
      RECT 1007.500000 366.350000 1008.500000 367.650000 ;
      RECT 966.500000 366.350000 999.500000 367.650000 ;
      RECT 957.500000 366.350000 958.500000 367.650000 ;
      RECT 916.500000 366.350000 949.500000 367.650000 ;
      RECT 907.500000 366.350000 908.500000 367.650000 ;
      RECT 866.500000 366.350000 899.500000 367.650000 ;
      RECT 857.500000 366.350000 858.500000 367.650000 ;
      RECT 816.500000 366.350000 849.500000 367.650000 ;
      RECT 807.500000 366.350000 808.500000 367.650000 ;
      RECT 766.500000 366.350000 799.500000 367.650000 ;
      RECT 757.500000 366.350000 758.500000 367.650000 ;
      RECT 716.500000 366.350000 749.500000 367.650000 ;
      RECT 707.500000 366.350000 708.500000 367.650000 ;
      RECT 666.500000 366.350000 699.500000 367.650000 ;
      RECT 657.500000 366.350000 658.500000 367.650000 ;
      RECT 616.500000 366.350000 649.500000 367.650000 ;
      RECT 607.500000 366.350000 608.500000 367.650000 ;
      RECT 566.500000 366.350000 599.500000 367.650000 ;
      RECT 557.500000 366.350000 558.500000 367.650000 ;
      RECT 516.500000 366.350000 549.500000 367.650000 ;
      RECT 507.500000 366.350000 508.500000 367.650000 ;
      RECT 416.500000 366.350000 449.500000 369.650000 ;
      RECT 407.500000 366.350000 408.500000 367.650000 ;
      RECT 366.500000 366.350000 399.500000 367.650000 ;
      RECT 357.500000 366.350000 358.500000 367.650000 ;
      RECT 316.500000 366.350000 349.500000 367.650000 ;
      RECT 307.500000 366.350000 308.500000 367.650000 ;
      RECT 266.500000 366.350000 299.500000 367.650000 ;
      RECT 257.500000 366.350000 258.500000 367.650000 ;
      RECT 216.500000 366.350000 249.500000 367.650000 ;
      RECT 207.500000 366.350000 208.500000 367.650000 ;
      RECT 166.500000 366.350000 199.500000 367.650000 ;
      RECT 157.500000 366.350000 158.500000 367.650000 ;
      RECT 116.500000 366.350000 149.500000 367.650000 ;
      RECT 107.500000 366.350000 108.500000 367.650000 ;
      RECT 66.500000 366.350000 99.500000 367.650000 ;
      RECT 57.500000 366.350000 58.500000 367.650000 ;
      RECT 29.500000 366.350000 49.500000 367.650000 ;
      RECT 15.500000 366.350000 16.500000 367.650000 ;
      RECT 1157.500000 365.650000 1170.500000 366.350000 ;
      RECT 1107.500000 365.650000 1149.500000 366.350000 ;
      RECT 1057.500000 365.650000 1099.500000 366.350000 ;
      RECT 1007.500000 365.650000 1049.500000 366.350000 ;
      RECT 957.500000 365.650000 999.500000 366.350000 ;
      RECT 907.500000 365.650000 949.500000 366.350000 ;
      RECT 857.500000 365.650000 899.500000 366.350000 ;
      RECT 807.500000 365.650000 849.500000 366.350000 ;
      RECT 757.500000 365.650000 799.500000 366.350000 ;
      RECT 707.500000 365.650000 749.500000 366.350000 ;
      RECT 657.500000 365.650000 699.500000 366.350000 ;
      RECT 607.500000 365.650000 649.500000 366.350000 ;
      RECT 557.500000 365.650000 599.500000 366.350000 ;
      RECT 507.500000 365.650000 549.500000 366.350000 ;
      RECT 407.500000 365.650000 449.500000 366.350000 ;
      RECT 357.500000 365.650000 399.500000 366.350000 ;
      RECT 307.500000 365.650000 349.500000 366.350000 ;
      RECT 257.500000 365.650000 299.500000 366.350000 ;
      RECT 207.500000 365.650000 249.500000 366.350000 ;
      RECT 157.500000 365.650000 199.500000 366.350000 ;
      RECT 107.500000 365.650000 149.500000 366.350000 ;
      RECT 57.500000 365.650000 99.500000 366.350000 ;
      RECT 15.500000 365.650000 49.500000 366.350000 ;
      RECT 457.500000 364.605000 499.500000 367.650000 ;
      RECT 416.500000 364.605000 449.500000 365.650000 ;
      RECT 1183.500000 364.350000 1186.000000 367.650000 ;
      RECT 1169.500000 364.350000 1170.500000 365.650000 ;
      RECT 1116.500000 364.350000 1149.500000 365.650000 ;
      RECT 1107.500000 364.350000 1108.500000 365.650000 ;
      RECT 1066.500000 364.350000 1099.500000 365.650000 ;
      RECT 1057.500000 364.350000 1058.500000 365.650000 ;
      RECT 1016.500000 364.350000 1049.500000 365.650000 ;
      RECT 1007.500000 364.350000 1008.500000 365.650000 ;
      RECT 966.500000 364.350000 999.500000 365.650000 ;
      RECT 957.500000 364.350000 958.500000 365.650000 ;
      RECT 916.500000 364.350000 949.500000 365.650000 ;
      RECT 907.500000 364.350000 908.500000 365.650000 ;
      RECT 866.500000 364.350000 899.500000 365.650000 ;
      RECT 857.500000 364.350000 858.500000 365.650000 ;
      RECT 816.500000 364.350000 849.500000 365.650000 ;
      RECT 807.500000 364.350000 808.500000 365.650000 ;
      RECT 766.500000 364.350000 799.500000 365.650000 ;
      RECT 757.500000 364.350000 758.500000 365.650000 ;
      RECT 716.500000 364.350000 749.500000 365.650000 ;
      RECT 707.500000 364.350000 708.500000 365.650000 ;
      RECT 666.500000 364.350000 699.500000 365.650000 ;
      RECT 657.500000 364.350000 658.500000 365.650000 ;
      RECT 616.500000 364.350000 649.500000 365.650000 ;
      RECT 607.500000 364.350000 608.500000 365.650000 ;
      RECT 566.500000 364.350000 599.500000 365.650000 ;
      RECT 557.500000 364.350000 558.500000 365.650000 ;
      RECT 516.500000 364.350000 549.500000 365.650000 ;
      RECT 507.500000 364.350000 508.500000 365.650000 ;
      RECT 416.500000 364.350000 499.500000 364.605000 ;
      RECT 407.500000 364.350000 408.500000 365.650000 ;
      RECT 366.500000 364.350000 399.500000 365.650000 ;
      RECT 357.500000 364.350000 358.500000 365.650000 ;
      RECT 316.500000 364.350000 349.500000 365.650000 ;
      RECT 307.500000 364.350000 308.500000 365.650000 ;
      RECT 266.500000 364.350000 299.500000 365.650000 ;
      RECT 257.500000 364.350000 258.500000 365.650000 ;
      RECT 216.500000 364.350000 249.500000 365.650000 ;
      RECT 207.500000 364.350000 208.500000 365.650000 ;
      RECT 166.500000 364.350000 199.500000 365.650000 ;
      RECT 157.500000 364.350000 158.500000 365.650000 ;
      RECT 116.500000 364.350000 149.500000 365.650000 ;
      RECT 107.500000 364.350000 108.500000 365.650000 ;
      RECT 66.500000 364.350000 99.500000 365.650000 ;
      RECT 57.500000 364.350000 58.500000 365.650000 ;
      RECT 29.500000 364.350000 49.500000 365.650000 ;
      RECT 15.500000 364.350000 16.500000 365.650000 ;
      RECT 0.000000 364.350000 2.500000 367.650000 ;
      RECT 1169.500000 363.650000 1186.000000 364.350000 ;
      RECT 1116.500000 363.650000 1156.500000 364.350000 ;
      RECT 1066.500000 363.650000 1108.500000 364.350000 ;
      RECT 1016.500000 363.650000 1058.500000 364.350000 ;
      RECT 966.500000 363.650000 1008.500000 364.350000 ;
      RECT 916.500000 363.650000 958.500000 364.350000 ;
      RECT 866.500000 363.650000 908.500000 364.350000 ;
      RECT 816.500000 363.650000 858.500000 364.350000 ;
      RECT 766.500000 363.650000 808.500000 364.350000 ;
      RECT 716.500000 363.650000 758.500000 364.350000 ;
      RECT 666.500000 363.650000 708.500000 364.350000 ;
      RECT 616.500000 363.650000 658.500000 364.350000 ;
      RECT 566.500000 363.650000 608.500000 364.350000 ;
      RECT 516.500000 363.650000 558.500000 364.350000 ;
      RECT 416.500000 363.650000 508.500000 364.350000 ;
      RECT 366.500000 363.650000 408.500000 364.350000 ;
      RECT 316.500000 363.650000 358.500000 364.350000 ;
      RECT 266.500000 363.650000 308.500000 364.350000 ;
      RECT 216.500000 363.650000 258.500000 364.350000 ;
      RECT 166.500000 363.650000 208.500000 364.350000 ;
      RECT 116.500000 363.650000 158.500000 364.350000 ;
      RECT 66.500000 363.650000 108.500000 364.350000 ;
      RECT 29.500000 363.650000 58.500000 364.350000 ;
      RECT 0.000000 363.650000 16.500000 364.350000 ;
      RECT 1169.500000 362.350000 1170.500000 363.650000 ;
      RECT 1116.500000 362.350000 1149.500000 363.650000 ;
      RECT 1107.500000 362.350000 1108.500000 363.650000 ;
      RECT 1066.500000 362.350000 1099.500000 363.650000 ;
      RECT 1057.500000 362.350000 1058.500000 363.650000 ;
      RECT 1016.500000 362.350000 1049.500000 363.650000 ;
      RECT 1007.500000 362.350000 1008.500000 363.650000 ;
      RECT 966.500000 362.350000 999.500000 363.650000 ;
      RECT 957.500000 362.350000 958.500000 363.650000 ;
      RECT 916.500000 362.350000 949.500000 363.650000 ;
      RECT 907.500000 362.350000 908.500000 363.650000 ;
      RECT 866.500000 362.350000 899.500000 363.650000 ;
      RECT 857.500000 362.350000 858.500000 363.650000 ;
      RECT 816.500000 362.350000 849.500000 363.650000 ;
      RECT 807.500000 362.350000 808.500000 363.650000 ;
      RECT 766.500000 362.350000 799.500000 363.650000 ;
      RECT 757.500000 362.350000 758.500000 363.650000 ;
      RECT 716.500000 362.350000 749.500000 363.650000 ;
      RECT 707.500000 362.350000 708.500000 363.650000 ;
      RECT 666.500000 362.350000 699.500000 363.650000 ;
      RECT 657.500000 362.350000 658.500000 363.650000 ;
      RECT 616.500000 362.350000 649.500000 363.650000 ;
      RECT 607.500000 362.350000 608.500000 363.650000 ;
      RECT 566.500000 362.350000 599.500000 363.650000 ;
      RECT 557.500000 362.350000 558.500000 363.650000 ;
      RECT 516.500000 362.350000 549.500000 363.650000 ;
      RECT 507.500000 362.350000 508.500000 363.650000 ;
      RECT 416.500000 362.350000 499.500000 363.650000 ;
      RECT 407.500000 362.350000 408.500000 363.650000 ;
      RECT 366.500000 362.350000 399.500000 363.650000 ;
      RECT 357.500000 362.350000 358.500000 363.650000 ;
      RECT 316.500000 362.350000 349.500000 363.650000 ;
      RECT 307.500000 362.350000 308.500000 363.650000 ;
      RECT 266.500000 362.350000 299.500000 363.650000 ;
      RECT 257.500000 362.350000 258.500000 363.650000 ;
      RECT 216.500000 362.350000 249.500000 363.650000 ;
      RECT 207.500000 362.350000 208.500000 363.650000 ;
      RECT 166.500000 362.350000 199.500000 363.650000 ;
      RECT 157.500000 362.350000 158.500000 363.650000 ;
      RECT 116.500000 362.350000 149.500000 363.650000 ;
      RECT 107.500000 362.350000 108.500000 363.650000 ;
      RECT 66.500000 362.350000 99.500000 363.650000 ;
      RECT 57.500000 362.350000 58.500000 363.650000 ;
      RECT 29.500000 362.350000 49.500000 363.650000 ;
      RECT 15.500000 362.350000 16.500000 363.650000 ;
      RECT 1157.500000 361.650000 1170.500000 362.350000 ;
      RECT 1107.500000 361.650000 1149.500000 362.350000 ;
      RECT 1057.500000 361.650000 1099.500000 362.350000 ;
      RECT 1007.500000 361.650000 1049.500000 362.350000 ;
      RECT 957.500000 361.650000 999.500000 362.350000 ;
      RECT 907.500000 361.650000 949.500000 362.350000 ;
      RECT 857.500000 361.650000 899.500000 362.350000 ;
      RECT 807.500000 361.650000 849.500000 362.350000 ;
      RECT 757.500000 361.650000 799.500000 362.350000 ;
      RECT 707.500000 361.650000 749.500000 362.350000 ;
      RECT 657.500000 361.650000 699.500000 362.350000 ;
      RECT 607.500000 361.650000 649.500000 362.350000 ;
      RECT 557.500000 361.650000 599.500000 362.350000 ;
      RECT 507.500000 361.650000 549.500000 362.350000 ;
      RECT 407.500000 361.650000 499.500000 362.350000 ;
      RECT 357.500000 361.650000 399.500000 362.350000 ;
      RECT 307.500000 361.650000 349.500000 362.350000 ;
      RECT 257.500000 361.650000 299.500000 362.350000 ;
      RECT 207.500000 361.650000 249.500000 362.350000 ;
      RECT 157.500000 361.650000 199.500000 362.350000 ;
      RECT 107.500000 361.650000 149.500000 362.350000 ;
      RECT 15.500000 361.650000 49.500000 362.350000 ;
      RECT 1183.500000 360.350000 1186.000000 363.650000 ;
      RECT 1169.500000 360.350000 1170.500000 361.650000 ;
      RECT 1116.500000 360.350000 1149.500000 361.650000 ;
      RECT 1107.500000 360.350000 1108.500000 361.650000 ;
      RECT 1066.500000 360.350000 1099.500000 361.650000 ;
      RECT 1057.500000 360.350000 1058.500000 361.650000 ;
      RECT 1016.500000 360.350000 1049.500000 361.650000 ;
      RECT 1007.500000 360.350000 1008.500000 361.650000 ;
      RECT 966.500000 360.350000 999.500000 361.650000 ;
      RECT 957.500000 360.350000 958.500000 361.650000 ;
      RECT 916.500000 360.350000 949.500000 361.650000 ;
      RECT 907.500000 360.350000 908.500000 361.650000 ;
      RECT 866.500000 360.350000 899.500000 361.650000 ;
      RECT 857.500000 360.350000 858.500000 361.650000 ;
      RECT 816.500000 360.350000 849.500000 361.650000 ;
      RECT 807.500000 360.350000 808.500000 361.650000 ;
      RECT 766.500000 360.350000 799.500000 361.650000 ;
      RECT 757.500000 360.350000 758.500000 361.650000 ;
      RECT 716.500000 360.350000 749.500000 361.650000 ;
      RECT 707.500000 360.350000 708.500000 361.650000 ;
      RECT 666.500000 360.350000 699.500000 361.650000 ;
      RECT 657.500000 360.350000 658.500000 361.650000 ;
      RECT 616.500000 360.350000 649.500000 361.650000 ;
      RECT 607.500000 360.350000 608.500000 361.650000 ;
      RECT 566.500000 360.350000 599.500000 361.650000 ;
      RECT 557.500000 360.350000 558.500000 361.650000 ;
      RECT 516.500000 360.350000 549.500000 361.650000 ;
      RECT 507.500000 360.350000 508.500000 361.650000 ;
      RECT 416.500000 360.350000 499.500000 361.650000 ;
      RECT 407.500000 360.350000 408.500000 361.650000 ;
      RECT 366.500000 360.350000 399.500000 361.650000 ;
      RECT 357.500000 360.350000 358.500000 361.650000 ;
      RECT 316.500000 360.350000 349.500000 361.650000 ;
      RECT 307.500000 360.350000 308.500000 361.650000 ;
      RECT 266.500000 360.350000 299.500000 361.650000 ;
      RECT 257.500000 360.350000 258.500000 361.650000 ;
      RECT 216.500000 360.350000 249.500000 361.650000 ;
      RECT 207.500000 360.350000 208.500000 361.650000 ;
      RECT 166.500000 360.350000 199.500000 361.650000 ;
      RECT 157.500000 360.350000 158.500000 361.650000 ;
      RECT 116.500000 360.350000 149.500000 361.650000 ;
      RECT 107.500000 360.350000 108.500000 361.650000 ;
      RECT 57.500000 360.350000 99.500000 362.350000 ;
      RECT 29.500000 360.350000 49.500000 361.650000 ;
      RECT 15.500000 360.350000 16.500000 361.650000 ;
      RECT 0.000000 360.350000 2.500000 363.650000 ;
      RECT 1169.500000 359.650000 1186.000000 360.350000 ;
      RECT 1116.500000 359.650000 1156.500000 360.350000 ;
      RECT 1066.500000 359.650000 1108.500000 360.350000 ;
      RECT 1016.500000 359.650000 1058.500000 360.350000 ;
      RECT 966.500000 359.650000 1008.500000 360.350000 ;
      RECT 916.500000 359.650000 958.500000 360.350000 ;
      RECT 866.500000 359.650000 908.500000 360.350000 ;
      RECT 816.500000 359.650000 858.500000 360.350000 ;
      RECT 766.500000 359.650000 808.500000 360.350000 ;
      RECT 716.500000 359.650000 758.500000 360.350000 ;
      RECT 666.500000 359.650000 708.500000 360.350000 ;
      RECT 616.500000 359.650000 658.500000 360.350000 ;
      RECT 566.500000 359.650000 608.500000 360.350000 ;
      RECT 516.500000 359.650000 558.500000 360.350000 ;
      RECT 416.500000 359.650000 508.500000 360.350000 ;
      RECT 366.500000 359.650000 408.500000 360.350000 ;
      RECT 316.500000 359.650000 358.500000 360.350000 ;
      RECT 266.500000 359.650000 308.500000 360.350000 ;
      RECT 216.500000 359.650000 258.500000 360.350000 ;
      RECT 166.500000 359.650000 208.500000 360.350000 ;
      RECT 116.500000 359.650000 158.500000 360.350000 ;
      RECT 29.500000 359.650000 108.500000 360.350000 ;
      RECT 0.000000 359.650000 16.500000 360.350000 ;
      RECT 1169.500000 358.350000 1170.500000 359.650000 ;
      RECT 1116.500000 358.350000 1149.500000 359.650000 ;
      RECT 1107.500000 358.350000 1108.500000 359.650000 ;
      RECT 1066.500000 358.350000 1099.500000 359.650000 ;
      RECT 1057.500000 358.350000 1058.500000 359.650000 ;
      RECT 1016.500000 358.350000 1049.500000 359.650000 ;
      RECT 1007.500000 358.350000 1008.500000 359.650000 ;
      RECT 966.500000 358.350000 999.500000 359.650000 ;
      RECT 957.500000 358.350000 958.500000 359.650000 ;
      RECT 916.500000 358.350000 949.500000 359.650000 ;
      RECT 907.500000 358.350000 908.500000 359.650000 ;
      RECT 866.500000 358.350000 899.500000 359.650000 ;
      RECT 857.500000 358.350000 858.500000 359.650000 ;
      RECT 816.500000 358.350000 849.500000 359.650000 ;
      RECT 807.500000 358.350000 808.500000 359.650000 ;
      RECT 766.500000 358.350000 799.500000 359.650000 ;
      RECT 757.500000 358.350000 758.500000 359.650000 ;
      RECT 716.500000 358.350000 749.500000 359.650000 ;
      RECT 707.500000 358.350000 708.500000 359.650000 ;
      RECT 666.500000 358.350000 699.500000 359.650000 ;
      RECT 657.500000 358.350000 658.500000 359.650000 ;
      RECT 616.500000 358.350000 649.500000 359.650000 ;
      RECT 607.500000 358.350000 608.500000 359.650000 ;
      RECT 566.500000 358.350000 599.500000 359.650000 ;
      RECT 557.500000 358.350000 558.500000 359.650000 ;
      RECT 516.500000 358.350000 549.500000 359.650000 ;
      RECT 507.500000 358.350000 508.500000 359.650000 ;
      RECT 416.500000 358.350000 499.500000 359.650000 ;
      RECT 407.500000 358.350000 408.500000 359.650000 ;
      RECT 366.500000 358.350000 399.500000 359.650000 ;
      RECT 357.500000 358.350000 358.500000 359.650000 ;
      RECT 316.500000 358.350000 349.500000 359.650000 ;
      RECT 307.500000 358.350000 308.500000 359.650000 ;
      RECT 266.500000 358.350000 299.500000 359.650000 ;
      RECT 257.500000 358.350000 258.500000 359.650000 ;
      RECT 216.500000 358.350000 249.500000 359.650000 ;
      RECT 207.500000 358.350000 208.500000 359.650000 ;
      RECT 166.500000 358.350000 199.500000 359.650000 ;
      RECT 157.500000 358.350000 158.500000 359.650000 ;
      RECT 116.500000 358.350000 149.500000 359.650000 ;
      RECT 107.500000 358.350000 108.500000 359.650000 ;
      RECT 29.500000 358.350000 99.500000 359.650000 ;
      RECT 15.500000 358.350000 16.500000 359.650000 ;
      RECT 1157.500000 357.650000 1170.500000 358.350000 ;
      RECT 1107.500000 357.650000 1149.500000 358.350000 ;
      RECT 1057.500000 357.650000 1099.500000 358.350000 ;
      RECT 1007.500000 357.650000 1049.500000 358.350000 ;
      RECT 957.500000 357.650000 999.500000 358.350000 ;
      RECT 907.500000 357.650000 949.500000 358.350000 ;
      RECT 857.500000 357.650000 899.500000 358.350000 ;
      RECT 807.500000 357.650000 849.500000 358.350000 ;
      RECT 757.500000 357.650000 799.500000 358.350000 ;
      RECT 707.500000 357.650000 749.500000 358.350000 ;
      RECT 657.500000 357.650000 699.500000 358.350000 ;
      RECT 607.500000 357.650000 649.500000 358.350000 ;
      RECT 557.500000 357.650000 599.500000 358.350000 ;
      RECT 507.500000 357.650000 549.500000 358.350000 ;
      RECT 407.500000 357.650000 499.500000 358.350000 ;
      RECT 357.500000 357.650000 399.500000 358.350000 ;
      RECT 307.500000 357.650000 349.500000 358.350000 ;
      RECT 257.500000 357.650000 299.500000 358.350000 ;
      RECT 207.500000 357.650000 249.500000 358.350000 ;
      RECT 157.500000 357.650000 199.500000 358.350000 ;
      RECT 107.500000 357.650000 149.500000 358.350000 ;
      RECT 15.500000 357.650000 99.500000 358.350000 ;
      RECT 1183.500000 356.350000 1186.000000 359.650000 ;
      RECT 1169.500000 356.350000 1170.500000 357.650000 ;
      RECT 1116.500000 356.350000 1149.500000 357.650000 ;
      RECT 1107.500000 356.350000 1108.500000 357.650000 ;
      RECT 1066.500000 356.350000 1099.500000 357.650000 ;
      RECT 1057.500000 356.350000 1058.500000 357.650000 ;
      RECT 1016.500000 356.350000 1049.500000 357.650000 ;
      RECT 1007.500000 356.350000 1008.500000 357.650000 ;
      RECT 966.500000 356.350000 999.500000 357.650000 ;
      RECT 957.500000 356.350000 958.500000 357.650000 ;
      RECT 916.500000 356.350000 949.500000 357.650000 ;
      RECT 907.500000 356.350000 908.500000 357.650000 ;
      RECT 866.500000 356.350000 899.500000 357.650000 ;
      RECT 857.500000 356.350000 858.500000 357.650000 ;
      RECT 816.500000 356.350000 849.500000 357.650000 ;
      RECT 807.500000 356.350000 808.500000 357.650000 ;
      RECT 766.500000 356.350000 799.500000 357.650000 ;
      RECT 757.500000 356.350000 758.500000 357.650000 ;
      RECT 716.500000 356.350000 749.500000 357.650000 ;
      RECT 707.500000 356.350000 708.500000 357.650000 ;
      RECT 666.500000 356.350000 699.500000 357.650000 ;
      RECT 657.500000 356.350000 658.500000 357.650000 ;
      RECT 616.500000 356.350000 649.500000 357.650000 ;
      RECT 607.500000 356.350000 608.500000 357.650000 ;
      RECT 566.500000 356.350000 599.500000 357.650000 ;
      RECT 557.500000 356.350000 558.500000 357.650000 ;
      RECT 516.500000 356.350000 549.500000 357.650000 ;
      RECT 507.500000 356.350000 508.500000 357.650000 ;
      RECT 416.500000 356.350000 499.500000 357.650000 ;
      RECT 407.500000 356.350000 408.500000 357.650000 ;
      RECT 366.500000 356.350000 399.500000 357.650000 ;
      RECT 357.500000 356.350000 358.500000 357.650000 ;
      RECT 316.500000 356.350000 349.500000 357.650000 ;
      RECT 307.500000 356.350000 308.500000 357.650000 ;
      RECT 266.500000 356.350000 299.500000 357.650000 ;
      RECT 257.500000 356.350000 258.500000 357.650000 ;
      RECT 216.500000 356.350000 249.500000 357.650000 ;
      RECT 207.500000 356.350000 208.500000 357.650000 ;
      RECT 166.500000 356.350000 199.500000 357.650000 ;
      RECT 157.500000 356.350000 158.500000 357.650000 ;
      RECT 116.500000 356.350000 149.500000 357.650000 ;
      RECT 107.500000 356.350000 108.500000 357.650000 ;
      RECT 29.500000 356.350000 99.500000 357.650000 ;
      RECT 15.500000 356.350000 16.500000 357.650000 ;
      RECT 0.000000 356.350000 2.500000 359.650000 ;
      RECT 29.500000 356.245000 108.500000 356.350000 ;
      RECT 1169.500000 355.650000 1186.000000 356.350000 ;
      RECT 1116.500000 355.650000 1156.500000 356.350000 ;
      RECT 1066.500000 355.650000 1108.500000 356.350000 ;
      RECT 1016.500000 355.650000 1058.500000 356.350000 ;
      RECT 966.500000 355.650000 1008.500000 356.350000 ;
      RECT 916.500000 355.650000 958.500000 356.350000 ;
      RECT 866.500000 355.650000 908.500000 356.350000 ;
      RECT 816.500000 355.650000 858.500000 356.350000 ;
      RECT 766.500000 355.650000 808.500000 356.350000 ;
      RECT 716.500000 355.650000 758.500000 356.350000 ;
      RECT 666.500000 355.650000 708.500000 356.350000 ;
      RECT 616.500000 355.650000 658.500000 356.350000 ;
      RECT 566.500000 355.650000 608.500000 356.350000 ;
      RECT 516.500000 355.650000 558.500000 356.350000 ;
      RECT 416.500000 355.650000 508.500000 356.350000 ;
      RECT 366.500000 355.650000 408.500000 356.350000 ;
      RECT 316.500000 355.650000 358.500000 356.350000 ;
      RECT 266.500000 355.650000 308.500000 356.350000 ;
      RECT 216.500000 355.650000 258.500000 356.350000 ;
      RECT 166.500000 355.650000 208.500000 356.350000 ;
      RECT 116.500000 355.650000 158.500000 356.350000 ;
      RECT 57.500000 355.650000 108.500000 356.245000 ;
      RECT 0.000000 355.650000 16.500000 356.350000 ;
      RECT 1169.500000 354.350000 1170.500000 355.650000 ;
      RECT 1116.500000 354.350000 1149.500000 355.650000 ;
      RECT 1107.500000 354.350000 1108.500000 355.650000 ;
      RECT 1066.500000 354.350000 1099.500000 355.650000 ;
      RECT 1057.500000 354.350000 1058.500000 355.650000 ;
      RECT 1016.500000 354.350000 1049.500000 355.650000 ;
      RECT 1007.500000 354.350000 1008.500000 355.650000 ;
      RECT 966.500000 354.350000 999.500000 355.650000 ;
      RECT 957.500000 354.350000 958.500000 355.650000 ;
      RECT 916.500000 354.350000 949.500000 355.650000 ;
      RECT 907.500000 354.350000 908.500000 355.650000 ;
      RECT 866.500000 354.350000 899.500000 355.650000 ;
      RECT 857.500000 354.350000 858.500000 355.650000 ;
      RECT 816.500000 354.350000 849.500000 355.650000 ;
      RECT 807.500000 354.350000 808.500000 355.650000 ;
      RECT 766.500000 354.350000 799.500000 355.650000 ;
      RECT 757.500000 354.350000 758.500000 355.650000 ;
      RECT 716.500000 354.350000 749.500000 355.650000 ;
      RECT 707.500000 354.350000 708.500000 355.650000 ;
      RECT 666.500000 354.350000 699.500000 355.650000 ;
      RECT 657.500000 354.350000 658.500000 355.650000 ;
      RECT 616.500000 354.350000 649.500000 355.650000 ;
      RECT 607.500000 354.350000 608.500000 355.650000 ;
      RECT 566.500000 354.350000 599.500000 355.650000 ;
      RECT 557.500000 354.350000 558.500000 355.650000 ;
      RECT 516.500000 354.350000 549.500000 355.650000 ;
      RECT 507.500000 354.350000 508.500000 355.650000 ;
      RECT 416.500000 354.350000 499.500000 355.650000 ;
      RECT 407.500000 354.350000 408.500000 355.650000 ;
      RECT 366.500000 354.350000 399.500000 355.650000 ;
      RECT 357.500000 354.350000 358.500000 355.650000 ;
      RECT 316.500000 354.350000 349.500000 355.650000 ;
      RECT 307.500000 354.350000 308.500000 355.650000 ;
      RECT 266.500000 354.350000 299.500000 355.650000 ;
      RECT 257.500000 354.350000 258.500000 355.650000 ;
      RECT 216.500000 354.350000 249.500000 355.650000 ;
      RECT 207.500000 354.350000 208.500000 355.650000 ;
      RECT 166.500000 354.350000 199.500000 355.650000 ;
      RECT 157.500000 354.350000 158.500000 355.650000 ;
      RECT 116.500000 354.350000 149.500000 355.650000 ;
      RECT 107.500000 354.350000 108.500000 355.650000 ;
      RECT 29.500000 354.350000 49.500000 356.245000 ;
      RECT 15.500000 354.350000 16.500000 355.650000 ;
      RECT 57.500000 354.245000 99.500000 355.650000 ;
      RECT 407.500000 353.730000 499.500000 354.350000 ;
      RECT 1157.500000 353.650000 1170.500000 354.350000 ;
      RECT 1107.500000 353.650000 1149.500000 354.350000 ;
      RECT 1057.500000 353.650000 1099.500000 354.350000 ;
      RECT 1007.500000 353.650000 1049.500000 354.350000 ;
      RECT 957.500000 353.650000 999.500000 354.350000 ;
      RECT 907.500000 353.650000 949.500000 354.350000 ;
      RECT 857.500000 353.650000 899.500000 354.350000 ;
      RECT 807.500000 353.650000 849.500000 354.350000 ;
      RECT 757.500000 353.650000 799.500000 354.350000 ;
      RECT 707.500000 353.650000 749.500000 354.350000 ;
      RECT 657.500000 353.650000 699.500000 354.350000 ;
      RECT 607.500000 353.650000 649.500000 354.350000 ;
      RECT 557.500000 353.650000 599.500000 354.350000 ;
      RECT 507.500000 353.650000 549.500000 354.350000 ;
      RECT 407.500000 353.650000 458.500000 353.730000 ;
      RECT 357.500000 353.650000 399.500000 354.350000 ;
      RECT 307.500000 353.650000 349.500000 354.350000 ;
      RECT 257.500000 353.650000 299.500000 354.350000 ;
      RECT 207.500000 353.650000 249.500000 354.350000 ;
      RECT 157.500000 353.650000 199.500000 354.350000 ;
      RECT 107.500000 353.650000 149.500000 354.350000 ;
      RECT 15.500000 353.650000 49.500000 354.350000 ;
      RECT 57.500000 352.945000 58.500000 354.245000 ;
      RECT 29.500000 352.945000 49.500000 353.650000 ;
      RECT 1183.500000 352.350000 1186.000000 355.650000 ;
      RECT 1169.500000 352.350000 1170.500000 353.650000 ;
      RECT 1116.500000 352.350000 1149.500000 353.650000 ;
      RECT 1107.500000 352.350000 1108.500000 353.650000 ;
      RECT 1066.500000 352.350000 1099.500000 353.650000 ;
      RECT 1057.500000 352.350000 1058.500000 353.650000 ;
      RECT 1016.500000 352.350000 1049.500000 353.650000 ;
      RECT 1007.500000 352.350000 1008.500000 353.650000 ;
      RECT 966.500000 352.350000 999.500000 353.650000 ;
      RECT 957.500000 352.350000 958.500000 353.650000 ;
      RECT 916.500000 352.350000 949.500000 353.650000 ;
      RECT 907.500000 352.350000 908.500000 353.650000 ;
      RECT 866.500000 352.350000 899.500000 353.650000 ;
      RECT 857.500000 352.350000 858.500000 353.650000 ;
      RECT 816.500000 352.350000 849.500000 353.650000 ;
      RECT 807.500000 352.350000 808.500000 353.650000 ;
      RECT 766.500000 352.350000 799.500000 353.650000 ;
      RECT 757.500000 352.350000 758.500000 353.650000 ;
      RECT 716.500000 352.350000 749.500000 353.650000 ;
      RECT 707.500000 352.350000 708.500000 353.650000 ;
      RECT 666.500000 352.350000 699.500000 353.650000 ;
      RECT 657.500000 352.350000 658.500000 353.650000 ;
      RECT 616.500000 352.350000 649.500000 353.650000 ;
      RECT 607.500000 352.350000 608.500000 353.650000 ;
      RECT 566.500000 352.350000 599.500000 353.650000 ;
      RECT 557.500000 352.350000 558.500000 353.650000 ;
      RECT 516.500000 352.350000 549.500000 353.650000 ;
      RECT 507.500000 352.350000 508.500000 353.650000 ;
      RECT 466.500000 352.350000 499.500000 353.730000 ;
      RECT 407.500000 352.350000 408.500000 353.650000 ;
      RECT 366.500000 352.350000 399.500000 353.650000 ;
      RECT 357.500000 352.350000 358.500000 353.650000 ;
      RECT 316.500000 352.350000 349.500000 353.650000 ;
      RECT 307.500000 352.350000 308.500000 353.650000 ;
      RECT 266.500000 352.350000 299.500000 353.650000 ;
      RECT 257.500000 352.350000 258.500000 353.650000 ;
      RECT 216.500000 352.350000 249.500000 353.650000 ;
      RECT 207.500000 352.350000 208.500000 353.650000 ;
      RECT 166.500000 352.350000 199.500000 353.650000 ;
      RECT 157.500000 352.350000 158.500000 353.650000 ;
      RECT 116.500000 352.350000 149.500000 353.650000 ;
      RECT 107.500000 352.350000 108.500000 353.650000 ;
      RECT 65.580000 352.350000 99.500000 354.245000 ;
      RECT 15.500000 352.350000 16.500000 353.650000 ;
      RECT 0.000000 352.350000 2.500000 355.650000 ;
      RECT 1169.500000 351.650000 1186.000000 352.350000 ;
      RECT 1116.500000 351.650000 1156.500000 352.350000 ;
      RECT 1066.500000 351.650000 1108.500000 352.350000 ;
      RECT 1016.500000 351.650000 1058.500000 352.350000 ;
      RECT 966.500000 351.650000 1008.500000 352.350000 ;
      RECT 916.500000 351.650000 958.500000 352.350000 ;
      RECT 866.500000 351.650000 908.500000 352.350000 ;
      RECT 816.500000 351.650000 858.500000 352.350000 ;
      RECT 766.500000 351.650000 808.500000 352.350000 ;
      RECT 716.500000 351.650000 758.500000 352.350000 ;
      RECT 666.500000 351.650000 708.500000 352.350000 ;
      RECT 616.500000 351.650000 658.500000 352.350000 ;
      RECT 566.500000 351.650000 608.500000 352.350000 ;
      RECT 516.500000 351.650000 558.500000 352.350000 ;
      RECT 466.500000 351.650000 508.500000 352.350000 ;
      RECT 366.500000 351.650000 408.500000 352.350000 ;
      RECT 316.500000 351.650000 358.500000 352.350000 ;
      RECT 266.500000 351.650000 308.500000 352.350000 ;
      RECT 216.500000 351.650000 258.500000 352.350000 ;
      RECT 166.500000 351.650000 208.500000 352.350000 ;
      RECT 116.500000 351.650000 158.500000 352.350000 ;
      RECT 65.580000 351.650000 108.500000 352.350000 ;
      RECT 0.000000 351.650000 16.500000 352.350000 ;
      RECT 65.580000 350.945000 99.500000 351.650000 ;
      RECT 29.500000 350.945000 58.500000 352.945000 ;
      RECT 1169.500000 350.350000 1170.500000 351.650000 ;
      RECT 1116.500000 350.350000 1149.500000 351.650000 ;
      RECT 1107.500000 350.350000 1108.500000 351.650000 ;
      RECT 1066.500000 350.350000 1099.500000 351.650000 ;
      RECT 1057.500000 350.350000 1058.500000 351.650000 ;
      RECT 1016.500000 350.350000 1049.500000 351.650000 ;
      RECT 1007.500000 350.350000 1008.500000 351.650000 ;
      RECT 966.500000 350.350000 999.500000 351.650000 ;
      RECT 957.500000 350.350000 958.500000 351.650000 ;
      RECT 916.500000 350.350000 949.500000 351.650000 ;
      RECT 907.500000 350.350000 908.500000 351.650000 ;
      RECT 866.500000 350.350000 899.500000 351.650000 ;
      RECT 857.500000 350.350000 858.500000 351.650000 ;
      RECT 816.500000 350.350000 849.500000 351.650000 ;
      RECT 807.500000 350.350000 808.500000 351.650000 ;
      RECT 766.500000 350.350000 799.500000 351.650000 ;
      RECT 757.500000 350.350000 758.500000 351.650000 ;
      RECT 716.500000 350.350000 749.500000 351.650000 ;
      RECT 707.500000 350.350000 708.500000 351.650000 ;
      RECT 666.500000 350.350000 699.500000 351.650000 ;
      RECT 657.500000 350.350000 658.500000 351.650000 ;
      RECT 616.500000 350.350000 649.500000 351.650000 ;
      RECT 607.500000 350.350000 608.500000 351.650000 ;
      RECT 566.500000 350.350000 599.500000 351.650000 ;
      RECT 557.500000 350.350000 558.500000 351.650000 ;
      RECT 516.500000 350.350000 549.500000 351.650000 ;
      RECT 507.500000 350.350000 508.500000 351.650000 ;
      RECT 416.500000 350.350000 458.500000 353.650000 ;
      RECT 407.500000 350.350000 408.500000 351.650000 ;
      RECT 366.500000 350.350000 399.500000 351.650000 ;
      RECT 357.500000 350.350000 358.500000 351.650000 ;
      RECT 316.500000 350.350000 349.500000 351.650000 ;
      RECT 307.500000 350.350000 308.500000 351.650000 ;
      RECT 266.500000 350.350000 299.500000 351.650000 ;
      RECT 257.500000 350.350000 258.500000 351.650000 ;
      RECT 216.500000 350.350000 249.500000 351.650000 ;
      RECT 207.500000 350.350000 208.500000 351.650000 ;
      RECT 166.500000 350.350000 199.500000 351.650000 ;
      RECT 157.500000 350.350000 158.500000 351.650000 ;
      RECT 116.500000 350.350000 149.500000 351.650000 ;
      RECT 107.500000 350.350000 108.500000 351.650000 ;
      RECT 29.500000 350.350000 99.500000 350.945000 ;
      RECT 15.500000 350.350000 16.500000 351.650000 ;
      RECT 466.500000 349.730000 499.500000 351.650000 ;
      RECT 407.500000 349.730000 458.500000 350.350000 ;
      RECT 1157.500000 349.650000 1170.500000 350.350000 ;
      RECT 1107.500000 349.650000 1149.500000 350.350000 ;
      RECT 1057.500000 349.650000 1099.500000 350.350000 ;
      RECT 1007.500000 349.650000 1049.500000 350.350000 ;
      RECT 957.500000 349.650000 999.500000 350.350000 ;
      RECT 907.500000 349.650000 949.500000 350.350000 ;
      RECT 857.500000 349.650000 899.500000 350.350000 ;
      RECT 807.500000 349.650000 849.500000 350.350000 ;
      RECT 757.500000 349.650000 799.500000 350.350000 ;
      RECT 707.500000 349.650000 749.500000 350.350000 ;
      RECT 657.500000 349.650000 699.500000 350.350000 ;
      RECT 607.500000 349.650000 649.500000 350.350000 ;
      RECT 557.500000 349.650000 599.500000 350.350000 ;
      RECT 507.500000 349.650000 549.500000 350.350000 ;
      RECT 407.500000 349.650000 499.500000 349.730000 ;
      RECT 357.500000 349.650000 399.500000 350.350000 ;
      RECT 307.500000 349.650000 349.500000 350.350000 ;
      RECT 257.500000 349.650000 299.500000 350.350000 ;
      RECT 207.500000 349.650000 249.500000 350.350000 ;
      RECT 157.500000 349.650000 199.500000 350.350000 ;
      RECT 107.500000 349.650000 149.500000 350.350000 ;
      RECT 15.500000 349.650000 99.500000 350.350000 ;
      RECT 1183.500000 348.350000 1186.000000 351.650000 ;
      RECT 1169.500000 348.350000 1170.500000 349.650000 ;
      RECT 1116.500000 348.350000 1149.500000 349.650000 ;
      RECT 1107.500000 348.350000 1108.500000 349.650000 ;
      RECT 1066.500000 348.350000 1099.500000 349.650000 ;
      RECT 1057.500000 348.350000 1058.500000 349.650000 ;
      RECT 1016.500000 348.350000 1049.500000 349.650000 ;
      RECT 1007.500000 348.350000 1008.500000 349.650000 ;
      RECT 966.500000 348.350000 999.500000 349.650000 ;
      RECT 957.500000 348.350000 958.500000 349.650000 ;
      RECT 916.500000 348.350000 949.500000 349.650000 ;
      RECT 907.500000 348.350000 908.500000 349.650000 ;
      RECT 866.500000 348.350000 899.500000 349.650000 ;
      RECT 857.500000 348.350000 858.500000 349.650000 ;
      RECT 816.500000 348.350000 849.500000 349.650000 ;
      RECT 807.500000 348.350000 808.500000 349.650000 ;
      RECT 766.500000 348.350000 799.500000 349.650000 ;
      RECT 757.500000 348.350000 758.500000 349.650000 ;
      RECT 716.500000 348.350000 749.500000 349.650000 ;
      RECT 707.500000 348.350000 708.500000 349.650000 ;
      RECT 666.500000 348.350000 699.500000 349.650000 ;
      RECT 657.500000 348.350000 658.500000 349.650000 ;
      RECT 616.500000 348.350000 649.500000 349.650000 ;
      RECT 607.500000 348.350000 608.500000 349.650000 ;
      RECT 566.500000 348.350000 599.500000 349.650000 ;
      RECT 557.500000 348.350000 558.500000 349.650000 ;
      RECT 516.500000 348.350000 549.500000 349.650000 ;
      RECT 507.500000 348.350000 508.500000 349.650000 ;
      RECT 466.500000 348.350000 499.500000 349.650000 ;
      RECT 407.500000 348.350000 408.500000 349.650000 ;
      RECT 366.500000 348.350000 399.500000 349.650000 ;
      RECT 357.500000 348.350000 358.500000 349.650000 ;
      RECT 316.500000 348.350000 349.500000 349.650000 ;
      RECT 307.500000 348.350000 308.500000 349.650000 ;
      RECT 266.500000 348.350000 299.500000 349.650000 ;
      RECT 257.500000 348.350000 258.500000 349.650000 ;
      RECT 216.500000 348.350000 249.500000 349.650000 ;
      RECT 207.500000 348.350000 208.500000 349.650000 ;
      RECT 166.500000 348.350000 199.500000 349.650000 ;
      RECT 157.500000 348.350000 158.500000 349.650000 ;
      RECT 116.500000 348.350000 149.500000 349.650000 ;
      RECT 107.500000 348.350000 108.500000 349.650000 ;
      RECT 66.500000 348.350000 99.500000 349.650000 ;
      RECT 15.500000 348.350000 16.500000 349.650000 ;
      RECT 0.000000 348.350000 2.500000 351.650000 ;
      RECT 1169.500000 347.650000 1186.000000 348.350000 ;
      RECT 1116.500000 347.650000 1156.500000 348.350000 ;
      RECT 1066.500000 347.650000 1108.500000 348.350000 ;
      RECT 1016.500000 347.650000 1058.500000 348.350000 ;
      RECT 966.500000 347.650000 1008.500000 348.350000 ;
      RECT 916.500000 347.650000 958.500000 348.350000 ;
      RECT 866.500000 347.650000 908.500000 348.350000 ;
      RECT 816.500000 347.650000 858.500000 348.350000 ;
      RECT 766.500000 347.650000 808.500000 348.350000 ;
      RECT 716.500000 347.650000 758.500000 348.350000 ;
      RECT 666.500000 347.650000 708.500000 348.350000 ;
      RECT 616.500000 347.650000 658.500000 348.350000 ;
      RECT 566.500000 347.650000 608.500000 348.350000 ;
      RECT 516.500000 347.650000 558.500000 348.350000 ;
      RECT 466.500000 347.650000 508.500000 348.350000 ;
      RECT 416.500000 347.650000 458.500000 349.650000 ;
      RECT 366.500000 347.650000 408.500000 348.350000 ;
      RECT 316.500000 347.650000 358.500000 348.350000 ;
      RECT 266.500000 347.650000 308.500000 348.350000 ;
      RECT 216.500000 347.650000 258.500000 348.350000 ;
      RECT 166.500000 347.650000 208.500000 348.350000 ;
      RECT 116.500000 347.650000 158.500000 348.350000 ;
      RECT 66.500000 347.650000 108.500000 348.350000 ;
      RECT 29.500000 347.650000 58.500000 349.650000 ;
      RECT 0.000000 347.650000 16.500000 348.350000 ;
      RECT 1169.500000 346.350000 1170.500000 347.650000 ;
      RECT 1116.500000 346.350000 1149.500000 347.650000 ;
      RECT 1107.500000 346.350000 1108.500000 347.650000 ;
      RECT 1066.500000 346.350000 1099.500000 347.650000 ;
      RECT 1057.500000 346.350000 1058.500000 347.650000 ;
      RECT 1016.500000 346.350000 1049.500000 347.650000 ;
      RECT 1007.500000 346.350000 1008.500000 347.650000 ;
      RECT 966.500000 346.350000 999.500000 347.650000 ;
      RECT 957.500000 346.350000 958.500000 347.650000 ;
      RECT 916.500000 346.350000 949.500000 347.650000 ;
      RECT 907.500000 346.350000 908.500000 347.650000 ;
      RECT 866.500000 346.350000 899.500000 347.650000 ;
      RECT 857.500000 346.350000 858.500000 347.650000 ;
      RECT 816.500000 346.350000 849.500000 347.650000 ;
      RECT 807.500000 346.350000 808.500000 347.650000 ;
      RECT 766.500000 346.350000 799.500000 347.650000 ;
      RECT 757.500000 346.350000 758.500000 347.650000 ;
      RECT 716.500000 346.350000 749.500000 347.650000 ;
      RECT 707.500000 346.350000 708.500000 347.650000 ;
      RECT 666.500000 346.350000 699.500000 347.650000 ;
      RECT 657.500000 346.350000 658.500000 347.650000 ;
      RECT 616.500000 346.350000 649.500000 347.650000 ;
      RECT 607.500000 346.350000 608.500000 347.650000 ;
      RECT 566.500000 346.350000 599.500000 347.650000 ;
      RECT 557.500000 346.350000 558.500000 347.650000 ;
      RECT 516.500000 346.350000 549.500000 347.650000 ;
      RECT 507.500000 346.350000 508.500000 347.650000 ;
      RECT 466.500000 346.350000 499.500000 347.650000 ;
      RECT 457.500000 346.350000 458.500000 347.650000 ;
      RECT 416.500000 346.350000 449.500000 347.650000 ;
      RECT 407.500000 346.350000 408.500000 347.650000 ;
      RECT 366.500000 346.350000 399.500000 347.650000 ;
      RECT 357.500000 346.350000 358.500000 347.650000 ;
      RECT 316.500000 346.350000 349.500000 347.650000 ;
      RECT 307.500000 346.350000 308.500000 347.650000 ;
      RECT 266.500000 346.350000 299.500000 347.650000 ;
      RECT 257.500000 346.350000 258.500000 347.650000 ;
      RECT 216.500000 346.350000 249.500000 347.650000 ;
      RECT 207.500000 346.350000 208.500000 347.650000 ;
      RECT 166.500000 346.350000 199.500000 347.650000 ;
      RECT 157.500000 346.350000 158.500000 347.650000 ;
      RECT 116.500000 346.350000 149.500000 347.650000 ;
      RECT 107.500000 346.350000 108.500000 347.650000 ;
      RECT 66.500000 346.350000 99.500000 347.650000 ;
      RECT 57.500000 346.350000 58.500000 347.650000 ;
      RECT 29.500000 346.350000 49.500000 347.650000 ;
      RECT 15.500000 346.350000 16.500000 347.650000 ;
      RECT 1157.500000 345.650000 1170.500000 346.350000 ;
      RECT 1107.500000 345.650000 1149.500000 346.350000 ;
      RECT 1057.500000 345.650000 1099.500000 346.350000 ;
      RECT 1007.500000 345.650000 1049.500000 346.350000 ;
      RECT 957.500000 345.650000 999.500000 346.350000 ;
      RECT 907.500000 345.650000 949.500000 346.350000 ;
      RECT 857.500000 345.650000 899.500000 346.350000 ;
      RECT 807.500000 345.650000 849.500000 346.350000 ;
      RECT 757.500000 345.650000 799.500000 346.350000 ;
      RECT 707.500000 345.650000 749.500000 346.350000 ;
      RECT 657.500000 345.650000 699.500000 346.350000 ;
      RECT 607.500000 345.650000 649.500000 346.350000 ;
      RECT 557.500000 345.650000 599.500000 346.350000 ;
      RECT 507.500000 345.650000 549.500000 346.350000 ;
      RECT 457.500000 345.650000 499.500000 346.350000 ;
      RECT 407.500000 345.650000 449.500000 346.350000 ;
      RECT 357.500000 345.650000 399.500000 346.350000 ;
      RECT 307.500000 345.650000 349.500000 346.350000 ;
      RECT 257.500000 345.650000 299.500000 346.350000 ;
      RECT 207.500000 345.650000 249.500000 346.350000 ;
      RECT 157.500000 345.650000 199.500000 346.350000 ;
      RECT 107.500000 345.650000 149.500000 346.350000 ;
      RECT 57.500000 345.650000 99.500000 346.350000 ;
      RECT 15.500000 345.650000 49.500000 346.350000 ;
      RECT 1183.500000 344.350000 1186.000000 347.650000 ;
      RECT 1169.500000 344.350000 1170.500000 345.650000 ;
      RECT 1116.500000 344.350000 1149.500000 345.650000 ;
      RECT 1107.500000 344.350000 1108.500000 345.650000 ;
      RECT 1066.500000 344.350000 1099.500000 345.650000 ;
      RECT 1057.500000 344.350000 1058.500000 345.650000 ;
      RECT 1016.500000 344.350000 1049.500000 345.650000 ;
      RECT 1007.500000 344.350000 1008.500000 345.650000 ;
      RECT 966.500000 344.350000 999.500000 345.650000 ;
      RECT 957.500000 344.350000 958.500000 345.650000 ;
      RECT 916.500000 344.350000 949.500000 345.650000 ;
      RECT 907.500000 344.350000 908.500000 345.650000 ;
      RECT 866.500000 344.350000 899.500000 345.650000 ;
      RECT 857.500000 344.350000 858.500000 345.650000 ;
      RECT 816.500000 344.350000 849.500000 345.650000 ;
      RECT 807.500000 344.350000 808.500000 345.650000 ;
      RECT 766.500000 344.350000 799.500000 345.650000 ;
      RECT 757.500000 344.350000 758.500000 345.650000 ;
      RECT 716.500000 344.350000 749.500000 345.650000 ;
      RECT 707.500000 344.350000 708.500000 345.650000 ;
      RECT 666.500000 344.350000 699.500000 345.650000 ;
      RECT 657.500000 344.350000 658.500000 345.650000 ;
      RECT 616.500000 344.350000 649.500000 345.650000 ;
      RECT 607.500000 344.350000 608.500000 345.650000 ;
      RECT 566.500000 344.350000 599.500000 345.650000 ;
      RECT 557.500000 344.350000 558.500000 345.650000 ;
      RECT 516.500000 344.350000 549.500000 345.650000 ;
      RECT 507.500000 344.350000 508.500000 345.650000 ;
      RECT 466.500000 344.350000 499.500000 345.650000 ;
      RECT 457.500000 344.350000 458.500000 345.650000 ;
      RECT 416.500000 344.350000 449.500000 345.650000 ;
      RECT 407.500000 344.350000 408.500000 345.650000 ;
      RECT 366.500000 344.350000 399.500000 345.650000 ;
      RECT 357.500000 344.350000 358.500000 345.650000 ;
      RECT 316.500000 344.350000 349.500000 345.650000 ;
      RECT 307.500000 344.350000 308.500000 345.650000 ;
      RECT 266.500000 344.350000 299.500000 345.650000 ;
      RECT 257.500000 344.350000 258.500000 345.650000 ;
      RECT 216.500000 344.350000 249.500000 345.650000 ;
      RECT 207.500000 344.350000 208.500000 345.650000 ;
      RECT 166.500000 344.350000 199.500000 345.650000 ;
      RECT 157.500000 344.350000 158.500000 345.650000 ;
      RECT 116.500000 344.350000 149.500000 345.650000 ;
      RECT 107.500000 344.350000 108.500000 345.650000 ;
      RECT 66.500000 344.350000 99.500000 345.650000 ;
      RECT 57.500000 344.350000 58.500000 345.650000 ;
      RECT 29.500000 344.350000 49.500000 345.650000 ;
      RECT 15.500000 344.350000 16.500000 345.650000 ;
      RECT 0.000000 344.350000 2.500000 347.650000 ;
      RECT 1169.500000 343.650000 1186.000000 344.350000 ;
      RECT 1116.500000 343.650000 1156.500000 344.350000 ;
      RECT 1066.500000 343.650000 1108.500000 344.350000 ;
      RECT 1016.500000 343.650000 1058.500000 344.350000 ;
      RECT 966.500000 343.650000 1008.500000 344.350000 ;
      RECT 916.500000 343.650000 958.500000 344.350000 ;
      RECT 866.500000 343.650000 908.500000 344.350000 ;
      RECT 816.500000 343.650000 858.500000 344.350000 ;
      RECT 766.500000 343.650000 808.500000 344.350000 ;
      RECT 716.500000 343.650000 758.500000 344.350000 ;
      RECT 666.500000 343.650000 708.500000 344.350000 ;
      RECT 616.500000 343.650000 658.500000 344.350000 ;
      RECT 566.500000 343.650000 608.500000 344.350000 ;
      RECT 516.500000 343.650000 558.500000 344.350000 ;
      RECT 466.500000 343.650000 508.500000 344.350000 ;
      RECT 416.500000 343.650000 458.500000 344.350000 ;
      RECT 366.500000 343.650000 408.500000 344.350000 ;
      RECT 316.500000 343.650000 358.500000 344.350000 ;
      RECT 266.500000 343.650000 308.500000 344.350000 ;
      RECT 216.500000 343.650000 258.500000 344.350000 ;
      RECT 166.500000 343.650000 208.500000 344.350000 ;
      RECT 116.500000 343.650000 158.500000 344.350000 ;
      RECT 66.500000 343.650000 108.500000 344.350000 ;
      RECT 29.500000 343.650000 58.500000 344.350000 ;
      RECT 0.000000 343.650000 16.500000 344.350000 ;
      RECT 1169.500000 342.350000 1170.500000 343.650000 ;
      RECT 1116.500000 342.350000 1149.500000 343.650000 ;
      RECT 1107.500000 342.350000 1108.500000 343.650000 ;
      RECT 1066.500000 342.350000 1099.500000 343.650000 ;
      RECT 1057.500000 342.350000 1058.500000 343.650000 ;
      RECT 1016.500000 342.350000 1049.500000 343.650000 ;
      RECT 1007.500000 342.350000 1008.500000 343.650000 ;
      RECT 966.500000 342.350000 999.500000 343.650000 ;
      RECT 957.500000 342.350000 958.500000 343.650000 ;
      RECT 916.500000 342.350000 949.500000 343.650000 ;
      RECT 907.500000 342.350000 908.500000 343.650000 ;
      RECT 866.500000 342.350000 899.500000 343.650000 ;
      RECT 857.500000 342.350000 858.500000 343.650000 ;
      RECT 816.500000 342.350000 849.500000 343.650000 ;
      RECT 807.500000 342.350000 808.500000 343.650000 ;
      RECT 766.500000 342.350000 799.500000 343.650000 ;
      RECT 757.500000 342.350000 758.500000 343.650000 ;
      RECT 716.500000 342.350000 749.500000 343.650000 ;
      RECT 707.500000 342.350000 708.500000 343.650000 ;
      RECT 666.500000 342.350000 699.500000 343.650000 ;
      RECT 657.500000 342.350000 658.500000 343.650000 ;
      RECT 616.500000 342.350000 649.500000 343.650000 ;
      RECT 607.500000 342.350000 608.500000 343.650000 ;
      RECT 566.500000 342.350000 599.500000 343.650000 ;
      RECT 557.500000 342.350000 558.500000 343.650000 ;
      RECT 516.500000 342.350000 549.500000 343.650000 ;
      RECT 507.500000 342.350000 508.500000 343.650000 ;
      RECT 466.500000 342.350000 499.500000 343.650000 ;
      RECT 457.500000 342.350000 458.500000 343.650000 ;
      RECT 416.500000 342.350000 449.500000 343.650000 ;
      RECT 407.500000 342.350000 408.500000 343.650000 ;
      RECT 366.500000 342.350000 399.500000 343.650000 ;
      RECT 357.500000 342.350000 358.500000 343.650000 ;
      RECT 316.500000 342.350000 349.500000 343.650000 ;
      RECT 307.500000 342.350000 308.500000 343.650000 ;
      RECT 266.500000 342.350000 299.500000 343.650000 ;
      RECT 257.500000 342.350000 258.500000 343.650000 ;
      RECT 216.500000 342.350000 249.500000 343.650000 ;
      RECT 207.500000 342.350000 208.500000 343.650000 ;
      RECT 166.500000 342.350000 199.500000 343.650000 ;
      RECT 157.500000 342.350000 158.500000 343.650000 ;
      RECT 116.500000 342.350000 149.500000 343.650000 ;
      RECT 107.500000 342.350000 108.500000 343.650000 ;
      RECT 66.500000 342.350000 99.500000 343.650000 ;
      RECT 57.500000 342.350000 58.500000 343.650000 ;
      RECT 29.500000 342.350000 49.500000 343.650000 ;
      RECT 15.500000 342.350000 16.500000 343.650000 ;
      RECT 1157.500000 341.650000 1170.500000 342.350000 ;
      RECT 1107.500000 341.650000 1149.500000 342.350000 ;
      RECT 1057.500000 341.650000 1099.500000 342.350000 ;
      RECT 1007.500000 341.650000 1049.500000 342.350000 ;
      RECT 957.500000 341.650000 999.500000 342.350000 ;
      RECT 907.500000 341.650000 949.500000 342.350000 ;
      RECT 857.500000 341.650000 899.500000 342.350000 ;
      RECT 807.500000 341.650000 849.500000 342.350000 ;
      RECT 757.500000 341.650000 799.500000 342.350000 ;
      RECT 707.500000 341.650000 749.500000 342.350000 ;
      RECT 657.500000 341.650000 699.500000 342.350000 ;
      RECT 607.500000 341.650000 649.500000 342.350000 ;
      RECT 557.500000 341.650000 599.500000 342.350000 ;
      RECT 507.500000 341.650000 549.500000 342.350000 ;
      RECT 457.500000 341.650000 499.500000 342.350000 ;
      RECT 407.500000 341.650000 449.500000 342.350000 ;
      RECT 357.500000 341.650000 399.500000 342.350000 ;
      RECT 307.500000 341.650000 349.500000 342.350000 ;
      RECT 257.500000 341.650000 299.500000 342.350000 ;
      RECT 207.500000 341.650000 249.500000 342.350000 ;
      RECT 157.500000 341.650000 199.500000 342.350000 ;
      RECT 107.500000 341.650000 149.500000 342.350000 ;
      RECT 57.500000 341.650000 99.500000 342.350000 ;
      RECT 15.500000 341.650000 49.500000 342.350000 ;
      RECT 1183.500000 340.350000 1186.000000 343.650000 ;
      RECT 1169.500000 340.350000 1170.500000 341.650000 ;
      RECT 1116.500000 340.350000 1149.500000 341.650000 ;
      RECT 1107.500000 340.350000 1108.500000 341.650000 ;
      RECT 1066.500000 340.350000 1099.500000 341.650000 ;
      RECT 1057.500000 340.350000 1058.500000 341.650000 ;
      RECT 1016.500000 340.350000 1049.500000 341.650000 ;
      RECT 1007.500000 340.350000 1008.500000 341.650000 ;
      RECT 966.500000 340.350000 999.500000 341.650000 ;
      RECT 957.500000 340.350000 958.500000 341.650000 ;
      RECT 916.500000 340.350000 949.500000 341.650000 ;
      RECT 907.500000 340.350000 908.500000 341.650000 ;
      RECT 866.500000 340.350000 899.500000 341.650000 ;
      RECT 857.500000 340.350000 858.500000 341.650000 ;
      RECT 816.500000 340.350000 849.500000 341.650000 ;
      RECT 807.500000 340.350000 808.500000 341.650000 ;
      RECT 766.500000 340.350000 799.500000 341.650000 ;
      RECT 757.500000 340.350000 758.500000 341.650000 ;
      RECT 716.500000 340.350000 749.500000 341.650000 ;
      RECT 707.500000 340.350000 708.500000 341.650000 ;
      RECT 666.500000 340.350000 699.500000 341.650000 ;
      RECT 657.500000 340.350000 658.500000 341.650000 ;
      RECT 616.500000 340.350000 649.500000 341.650000 ;
      RECT 607.500000 340.350000 608.500000 341.650000 ;
      RECT 566.500000 340.350000 599.500000 341.650000 ;
      RECT 557.500000 340.350000 558.500000 341.650000 ;
      RECT 516.500000 340.350000 549.500000 341.650000 ;
      RECT 507.500000 340.350000 508.500000 341.650000 ;
      RECT 466.500000 340.350000 499.500000 341.650000 ;
      RECT 457.500000 340.350000 458.500000 341.650000 ;
      RECT 416.500000 340.350000 449.500000 341.650000 ;
      RECT 407.500000 340.350000 408.500000 341.650000 ;
      RECT 366.500000 340.350000 399.500000 341.650000 ;
      RECT 357.500000 340.350000 358.500000 341.650000 ;
      RECT 316.500000 340.350000 349.500000 341.650000 ;
      RECT 307.500000 340.350000 308.500000 341.650000 ;
      RECT 266.500000 340.350000 299.500000 341.650000 ;
      RECT 257.500000 340.350000 258.500000 341.650000 ;
      RECT 216.500000 340.350000 249.500000 341.650000 ;
      RECT 207.500000 340.350000 208.500000 341.650000 ;
      RECT 166.500000 340.350000 199.500000 341.650000 ;
      RECT 157.500000 340.350000 158.500000 341.650000 ;
      RECT 116.500000 340.350000 149.500000 341.650000 ;
      RECT 107.500000 340.350000 108.500000 341.650000 ;
      RECT 66.500000 340.350000 99.500000 341.650000 ;
      RECT 57.500000 340.350000 58.500000 341.650000 ;
      RECT 29.500000 340.350000 49.500000 341.650000 ;
      RECT 15.500000 340.350000 16.500000 341.650000 ;
      RECT 0.000000 340.350000 2.500000 343.650000 ;
      RECT 1169.500000 339.650000 1186.000000 340.350000 ;
      RECT 1116.500000 339.650000 1156.500000 340.350000 ;
      RECT 1066.500000 339.650000 1108.500000 340.350000 ;
      RECT 1016.500000 339.650000 1058.500000 340.350000 ;
      RECT 966.500000 339.650000 1008.500000 340.350000 ;
      RECT 916.500000 339.650000 958.500000 340.350000 ;
      RECT 866.500000 339.650000 908.500000 340.350000 ;
      RECT 816.500000 339.650000 858.500000 340.350000 ;
      RECT 766.500000 339.650000 808.500000 340.350000 ;
      RECT 716.500000 339.650000 758.500000 340.350000 ;
      RECT 666.500000 339.650000 708.500000 340.350000 ;
      RECT 616.500000 339.650000 658.500000 340.350000 ;
      RECT 566.500000 339.650000 608.500000 340.350000 ;
      RECT 516.500000 339.650000 558.500000 340.350000 ;
      RECT 466.500000 339.650000 508.500000 340.350000 ;
      RECT 416.500000 339.650000 458.500000 340.350000 ;
      RECT 366.500000 339.650000 408.500000 340.350000 ;
      RECT 316.500000 339.650000 358.500000 340.350000 ;
      RECT 266.500000 339.650000 308.500000 340.350000 ;
      RECT 216.500000 339.650000 258.500000 340.350000 ;
      RECT 166.500000 339.650000 208.500000 340.350000 ;
      RECT 116.500000 339.650000 158.500000 340.350000 ;
      RECT 66.500000 339.650000 108.500000 340.350000 ;
      RECT 29.500000 339.650000 58.500000 340.350000 ;
      RECT 0.000000 339.650000 16.500000 340.350000 ;
      RECT 1169.500000 338.350000 1170.500000 339.650000 ;
      RECT 1116.500000 338.350000 1149.500000 339.650000 ;
      RECT 1107.500000 338.350000 1108.500000 339.650000 ;
      RECT 1066.500000 338.350000 1099.500000 339.650000 ;
      RECT 1057.500000 338.350000 1058.500000 339.650000 ;
      RECT 1016.500000 338.350000 1049.500000 339.650000 ;
      RECT 1007.500000 338.350000 1008.500000 339.650000 ;
      RECT 966.500000 338.350000 999.500000 339.650000 ;
      RECT 957.500000 338.350000 958.500000 339.650000 ;
      RECT 916.500000 338.350000 949.500000 339.650000 ;
      RECT 907.500000 338.350000 908.500000 339.650000 ;
      RECT 866.500000 338.350000 899.500000 339.650000 ;
      RECT 857.500000 338.350000 858.500000 339.650000 ;
      RECT 816.500000 338.350000 849.500000 339.650000 ;
      RECT 807.500000 338.350000 808.500000 339.650000 ;
      RECT 766.500000 338.350000 799.500000 339.650000 ;
      RECT 757.500000 338.350000 758.500000 339.650000 ;
      RECT 716.500000 338.350000 749.500000 339.650000 ;
      RECT 707.500000 338.350000 708.500000 339.650000 ;
      RECT 666.500000 338.350000 699.500000 339.650000 ;
      RECT 657.500000 338.350000 658.500000 339.650000 ;
      RECT 616.500000 338.350000 649.500000 339.650000 ;
      RECT 607.500000 338.350000 608.500000 339.650000 ;
      RECT 566.500000 338.350000 599.500000 339.650000 ;
      RECT 557.500000 338.350000 558.500000 339.650000 ;
      RECT 516.500000 338.350000 549.500000 339.650000 ;
      RECT 507.500000 338.350000 508.500000 339.650000 ;
      RECT 466.500000 338.350000 499.500000 339.650000 ;
      RECT 457.500000 338.350000 458.500000 339.650000 ;
      RECT 416.500000 338.350000 449.500000 339.650000 ;
      RECT 407.500000 338.350000 408.500000 339.650000 ;
      RECT 366.500000 338.350000 399.500000 339.650000 ;
      RECT 357.500000 338.350000 358.500000 339.650000 ;
      RECT 316.500000 338.350000 349.500000 339.650000 ;
      RECT 307.500000 338.350000 308.500000 339.650000 ;
      RECT 266.500000 338.350000 299.500000 339.650000 ;
      RECT 257.500000 338.350000 258.500000 339.650000 ;
      RECT 216.500000 338.350000 249.500000 339.650000 ;
      RECT 207.500000 338.350000 208.500000 339.650000 ;
      RECT 166.500000 338.350000 199.500000 339.650000 ;
      RECT 157.500000 338.350000 158.500000 339.650000 ;
      RECT 116.500000 338.350000 149.500000 339.650000 ;
      RECT 107.500000 338.350000 108.500000 339.650000 ;
      RECT 66.500000 338.350000 99.500000 339.650000 ;
      RECT 57.500000 338.350000 58.500000 339.650000 ;
      RECT 29.500000 338.350000 49.500000 339.650000 ;
      RECT 15.500000 338.350000 16.500000 339.650000 ;
      RECT 1157.500000 337.650000 1170.500000 338.350000 ;
      RECT 1107.500000 337.650000 1149.500000 338.350000 ;
      RECT 1057.500000 337.650000 1099.500000 338.350000 ;
      RECT 1007.500000 337.650000 1049.500000 338.350000 ;
      RECT 957.500000 337.650000 999.500000 338.350000 ;
      RECT 907.500000 337.650000 949.500000 338.350000 ;
      RECT 857.500000 337.650000 899.500000 338.350000 ;
      RECT 807.500000 337.650000 849.500000 338.350000 ;
      RECT 757.500000 337.650000 799.500000 338.350000 ;
      RECT 707.500000 337.650000 749.500000 338.350000 ;
      RECT 657.500000 337.650000 699.500000 338.350000 ;
      RECT 607.500000 337.650000 649.500000 338.350000 ;
      RECT 557.500000 337.650000 599.500000 338.350000 ;
      RECT 507.500000 337.650000 549.500000 338.350000 ;
      RECT 457.500000 337.650000 499.500000 338.350000 ;
      RECT 407.500000 337.650000 449.500000 338.350000 ;
      RECT 357.500000 337.650000 399.500000 338.350000 ;
      RECT 307.500000 337.650000 349.500000 338.350000 ;
      RECT 257.500000 337.650000 299.500000 338.350000 ;
      RECT 207.500000 337.650000 249.500000 338.350000 ;
      RECT 157.500000 337.650000 199.500000 338.350000 ;
      RECT 107.500000 337.650000 149.500000 338.350000 ;
      RECT 57.500000 337.650000 99.500000 338.350000 ;
      RECT 15.500000 337.650000 49.500000 338.350000 ;
      RECT 1183.500000 336.350000 1186.000000 339.650000 ;
      RECT 1169.500000 336.350000 1170.500000 337.650000 ;
      RECT 1116.500000 336.350000 1149.500000 337.650000 ;
      RECT 1107.500000 336.350000 1108.500000 337.650000 ;
      RECT 1066.500000 336.350000 1099.500000 337.650000 ;
      RECT 1057.500000 336.350000 1058.500000 337.650000 ;
      RECT 1016.500000 336.350000 1049.500000 337.650000 ;
      RECT 1007.500000 336.350000 1008.500000 337.650000 ;
      RECT 966.500000 336.350000 999.500000 337.650000 ;
      RECT 957.500000 336.350000 958.500000 337.650000 ;
      RECT 916.500000 336.350000 949.500000 337.650000 ;
      RECT 907.500000 336.350000 908.500000 337.650000 ;
      RECT 866.500000 336.350000 899.500000 337.650000 ;
      RECT 857.500000 336.350000 858.500000 337.650000 ;
      RECT 816.500000 336.350000 849.500000 337.650000 ;
      RECT 807.500000 336.350000 808.500000 337.650000 ;
      RECT 766.500000 336.350000 799.500000 337.650000 ;
      RECT 757.500000 336.350000 758.500000 337.650000 ;
      RECT 716.500000 336.350000 749.500000 337.650000 ;
      RECT 707.500000 336.350000 708.500000 337.650000 ;
      RECT 666.500000 336.350000 699.500000 337.650000 ;
      RECT 657.500000 336.350000 658.500000 337.650000 ;
      RECT 616.500000 336.350000 649.500000 337.650000 ;
      RECT 607.500000 336.350000 608.500000 337.650000 ;
      RECT 566.500000 336.350000 599.500000 337.650000 ;
      RECT 557.500000 336.350000 558.500000 337.650000 ;
      RECT 516.500000 336.350000 549.500000 337.650000 ;
      RECT 507.500000 336.350000 508.500000 337.650000 ;
      RECT 466.500000 336.350000 499.500000 337.650000 ;
      RECT 457.500000 336.350000 458.500000 337.650000 ;
      RECT 416.500000 336.350000 449.500000 337.650000 ;
      RECT 407.500000 336.350000 408.500000 337.650000 ;
      RECT 366.500000 336.350000 399.500000 337.650000 ;
      RECT 357.500000 336.350000 358.500000 337.650000 ;
      RECT 316.500000 336.350000 349.500000 337.650000 ;
      RECT 307.500000 336.350000 308.500000 337.650000 ;
      RECT 266.500000 336.350000 299.500000 337.650000 ;
      RECT 257.500000 336.350000 258.500000 337.650000 ;
      RECT 216.500000 336.350000 249.500000 337.650000 ;
      RECT 207.500000 336.350000 208.500000 337.650000 ;
      RECT 166.500000 336.350000 199.500000 337.650000 ;
      RECT 157.500000 336.350000 158.500000 337.650000 ;
      RECT 116.500000 336.350000 149.500000 337.650000 ;
      RECT 107.500000 336.350000 108.500000 337.650000 ;
      RECT 66.500000 336.350000 99.500000 337.650000 ;
      RECT 57.500000 336.350000 58.500000 337.650000 ;
      RECT 29.500000 336.350000 49.500000 337.650000 ;
      RECT 15.500000 336.350000 16.500000 337.650000 ;
      RECT 0.000000 336.350000 2.500000 339.650000 ;
      RECT 1169.500000 335.650000 1186.000000 336.350000 ;
      RECT 1116.500000 335.650000 1156.500000 336.350000 ;
      RECT 1066.500000 335.650000 1108.500000 336.350000 ;
      RECT 1016.500000 335.650000 1058.500000 336.350000 ;
      RECT 966.500000 335.650000 1008.500000 336.350000 ;
      RECT 916.500000 335.650000 958.500000 336.350000 ;
      RECT 866.500000 335.650000 908.500000 336.350000 ;
      RECT 816.500000 335.650000 858.500000 336.350000 ;
      RECT 766.500000 335.650000 808.500000 336.350000 ;
      RECT 716.500000 335.650000 758.500000 336.350000 ;
      RECT 666.500000 335.650000 708.500000 336.350000 ;
      RECT 616.500000 335.650000 658.500000 336.350000 ;
      RECT 566.500000 335.650000 608.500000 336.350000 ;
      RECT 516.500000 335.650000 558.500000 336.350000 ;
      RECT 466.500000 335.650000 508.500000 336.350000 ;
      RECT 416.500000 335.650000 458.500000 336.350000 ;
      RECT 366.500000 335.650000 408.500000 336.350000 ;
      RECT 316.500000 335.650000 358.500000 336.350000 ;
      RECT 266.500000 335.650000 308.500000 336.350000 ;
      RECT 216.500000 335.650000 258.500000 336.350000 ;
      RECT 166.500000 335.650000 208.500000 336.350000 ;
      RECT 116.500000 335.650000 158.500000 336.350000 ;
      RECT 66.500000 335.650000 108.500000 336.350000 ;
      RECT 29.500000 335.650000 58.500000 336.350000 ;
      RECT 0.000000 335.650000 16.500000 336.350000 ;
      RECT 1169.500000 334.350000 1170.500000 335.650000 ;
      RECT 1116.500000 334.350000 1149.500000 335.650000 ;
      RECT 1107.500000 334.350000 1108.500000 335.650000 ;
      RECT 1066.500000 334.350000 1099.500000 335.650000 ;
      RECT 1057.500000 334.350000 1058.500000 335.650000 ;
      RECT 1016.500000 334.350000 1049.500000 335.650000 ;
      RECT 1007.500000 334.350000 1008.500000 335.650000 ;
      RECT 966.500000 334.350000 999.500000 335.650000 ;
      RECT 957.500000 334.350000 958.500000 335.650000 ;
      RECT 916.500000 334.350000 949.500000 335.650000 ;
      RECT 907.500000 334.350000 908.500000 335.650000 ;
      RECT 866.500000 334.350000 899.500000 335.650000 ;
      RECT 857.500000 334.350000 858.500000 335.650000 ;
      RECT 816.500000 334.350000 849.500000 335.650000 ;
      RECT 807.500000 334.350000 808.500000 335.650000 ;
      RECT 766.500000 334.350000 799.500000 335.650000 ;
      RECT 757.500000 334.350000 758.500000 335.650000 ;
      RECT 716.500000 334.350000 749.500000 335.650000 ;
      RECT 707.500000 334.350000 708.500000 335.650000 ;
      RECT 666.500000 334.350000 699.500000 335.650000 ;
      RECT 657.500000 334.350000 658.500000 335.650000 ;
      RECT 616.500000 334.350000 649.500000 335.650000 ;
      RECT 607.500000 334.350000 608.500000 335.650000 ;
      RECT 566.500000 334.350000 599.500000 335.650000 ;
      RECT 557.500000 334.350000 558.500000 335.650000 ;
      RECT 516.500000 334.350000 549.500000 335.650000 ;
      RECT 507.500000 334.350000 508.500000 335.650000 ;
      RECT 466.500000 334.350000 499.500000 335.650000 ;
      RECT 457.500000 334.350000 458.500000 335.650000 ;
      RECT 416.500000 334.350000 449.500000 335.650000 ;
      RECT 407.500000 334.350000 408.500000 335.650000 ;
      RECT 366.500000 334.350000 399.500000 335.650000 ;
      RECT 357.500000 334.350000 358.500000 335.650000 ;
      RECT 316.500000 334.350000 349.500000 335.650000 ;
      RECT 307.500000 334.350000 308.500000 335.650000 ;
      RECT 266.500000 334.350000 299.500000 335.650000 ;
      RECT 257.500000 334.350000 258.500000 335.650000 ;
      RECT 216.500000 334.350000 249.500000 335.650000 ;
      RECT 207.500000 334.350000 208.500000 335.650000 ;
      RECT 166.500000 334.350000 199.500000 335.650000 ;
      RECT 157.500000 334.350000 158.500000 335.650000 ;
      RECT 116.500000 334.350000 149.500000 335.650000 ;
      RECT 107.500000 334.350000 108.500000 335.650000 ;
      RECT 66.500000 334.350000 99.500000 335.650000 ;
      RECT 57.500000 334.350000 58.500000 335.650000 ;
      RECT 29.500000 334.350000 49.500000 335.650000 ;
      RECT 15.500000 334.350000 16.500000 335.650000 ;
      RECT 1157.500000 333.650000 1170.500000 334.350000 ;
      RECT 1107.500000 333.650000 1149.500000 334.350000 ;
      RECT 1057.500000 333.650000 1099.500000 334.350000 ;
      RECT 1007.500000 333.650000 1049.500000 334.350000 ;
      RECT 957.500000 333.650000 999.500000 334.350000 ;
      RECT 907.500000 333.650000 949.500000 334.350000 ;
      RECT 857.500000 333.650000 899.500000 334.350000 ;
      RECT 807.500000 333.650000 849.500000 334.350000 ;
      RECT 757.500000 333.650000 799.500000 334.350000 ;
      RECT 707.500000 333.650000 749.500000 334.350000 ;
      RECT 657.500000 333.650000 699.500000 334.350000 ;
      RECT 607.500000 333.650000 649.500000 334.350000 ;
      RECT 557.500000 333.650000 599.500000 334.350000 ;
      RECT 507.500000 333.650000 549.500000 334.350000 ;
      RECT 457.500000 333.650000 499.500000 334.350000 ;
      RECT 407.500000 333.650000 449.500000 334.350000 ;
      RECT 357.500000 333.650000 399.500000 334.350000 ;
      RECT 307.500000 333.650000 349.500000 334.350000 ;
      RECT 257.500000 333.650000 299.500000 334.350000 ;
      RECT 207.500000 333.650000 249.500000 334.350000 ;
      RECT 157.500000 333.650000 199.500000 334.350000 ;
      RECT 107.500000 333.650000 149.500000 334.350000 ;
      RECT 57.500000 333.650000 99.500000 334.350000 ;
      RECT 15.500000 333.650000 49.500000 334.350000 ;
      RECT 1183.500000 332.350000 1186.000000 335.650000 ;
      RECT 1169.500000 332.350000 1170.500000 333.650000 ;
      RECT 1116.500000 332.350000 1149.500000 333.650000 ;
      RECT 1107.500000 332.350000 1108.500000 333.650000 ;
      RECT 1066.500000 332.350000 1099.500000 333.650000 ;
      RECT 1057.500000 332.350000 1058.500000 333.650000 ;
      RECT 1016.500000 332.350000 1049.500000 333.650000 ;
      RECT 1007.500000 332.350000 1008.500000 333.650000 ;
      RECT 966.500000 332.350000 999.500000 333.650000 ;
      RECT 957.500000 332.350000 958.500000 333.650000 ;
      RECT 916.500000 332.350000 949.500000 333.650000 ;
      RECT 907.500000 332.350000 908.500000 333.650000 ;
      RECT 866.500000 332.350000 899.500000 333.650000 ;
      RECT 857.500000 332.350000 858.500000 333.650000 ;
      RECT 816.500000 332.350000 849.500000 333.650000 ;
      RECT 807.500000 332.350000 808.500000 333.650000 ;
      RECT 766.500000 332.350000 799.500000 333.650000 ;
      RECT 757.500000 332.350000 758.500000 333.650000 ;
      RECT 716.500000 332.350000 749.500000 333.650000 ;
      RECT 707.500000 332.350000 708.500000 333.650000 ;
      RECT 666.500000 332.350000 699.500000 333.650000 ;
      RECT 657.500000 332.350000 658.500000 333.650000 ;
      RECT 616.500000 332.350000 649.500000 333.650000 ;
      RECT 607.500000 332.350000 608.500000 333.650000 ;
      RECT 566.500000 332.350000 599.500000 333.650000 ;
      RECT 557.500000 332.350000 558.500000 333.650000 ;
      RECT 516.500000 332.350000 549.500000 333.650000 ;
      RECT 507.500000 332.350000 508.500000 333.650000 ;
      RECT 466.500000 332.350000 499.500000 333.650000 ;
      RECT 457.500000 332.350000 458.500000 333.650000 ;
      RECT 416.500000 332.350000 449.500000 333.650000 ;
      RECT 407.500000 332.350000 408.500000 333.650000 ;
      RECT 366.500000 332.350000 399.500000 333.650000 ;
      RECT 357.500000 332.350000 358.500000 333.650000 ;
      RECT 316.500000 332.350000 349.500000 333.650000 ;
      RECT 307.500000 332.350000 308.500000 333.650000 ;
      RECT 266.500000 332.350000 299.500000 333.650000 ;
      RECT 257.500000 332.350000 258.500000 333.650000 ;
      RECT 216.500000 332.350000 249.500000 333.650000 ;
      RECT 207.500000 332.350000 208.500000 333.650000 ;
      RECT 166.500000 332.350000 199.500000 333.650000 ;
      RECT 157.500000 332.350000 158.500000 333.650000 ;
      RECT 116.500000 332.350000 149.500000 333.650000 ;
      RECT 107.500000 332.350000 108.500000 333.650000 ;
      RECT 66.500000 332.350000 99.500000 333.650000 ;
      RECT 57.500000 332.350000 58.500000 333.650000 ;
      RECT 29.500000 332.350000 49.500000 333.650000 ;
      RECT 15.500000 332.350000 16.500000 333.650000 ;
      RECT 0.000000 332.350000 2.500000 335.650000 ;
      RECT 1169.500000 331.650000 1186.000000 332.350000 ;
      RECT 1116.500000 331.650000 1156.500000 332.350000 ;
      RECT 1066.500000 331.650000 1108.500000 332.350000 ;
      RECT 1016.500000 331.650000 1058.500000 332.350000 ;
      RECT 966.500000 331.650000 1008.500000 332.350000 ;
      RECT 916.500000 331.650000 958.500000 332.350000 ;
      RECT 866.500000 331.650000 908.500000 332.350000 ;
      RECT 816.500000 331.650000 858.500000 332.350000 ;
      RECT 766.500000 331.650000 808.500000 332.350000 ;
      RECT 716.500000 331.650000 758.500000 332.350000 ;
      RECT 666.500000 331.650000 708.500000 332.350000 ;
      RECT 616.500000 331.650000 658.500000 332.350000 ;
      RECT 566.500000 331.650000 608.500000 332.350000 ;
      RECT 516.500000 331.650000 558.500000 332.350000 ;
      RECT 466.500000 331.650000 508.500000 332.350000 ;
      RECT 416.500000 331.650000 458.500000 332.350000 ;
      RECT 366.500000 331.650000 408.500000 332.350000 ;
      RECT 316.500000 331.650000 358.500000 332.350000 ;
      RECT 266.500000 331.650000 308.500000 332.350000 ;
      RECT 216.500000 331.650000 258.500000 332.350000 ;
      RECT 166.500000 331.650000 208.500000 332.350000 ;
      RECT 116.500000 331.650000 158.500000 332.350000 ;
      RECT 66.500000 331.650000 108.500000 332.350000 ;
      RECT 29.500000 331.650000 58.500000 332.350000 ;
      RECT 0.000000 331.650000 16.500000 332.350000 ;
      RECT 1169.500000 330.350000 1170.500000 331.650000 ;
      RECT 1116.500000 330.350000 1149.500000 331.650000 ;
      RECT 1107.500000 330.350000 1108.500000 331.650000 ;
      RECT 1066.500000 330.350000 1099.500000 331.650000 ;
      RECT 1057.500000 330.350000 1058.500000 331.650000 ;
      RECT 1016.500000 330.350000 1049.500000 331.650000 ;
      RECT 1007.500000 330.350000 1008.500000 331.650000 ;
      RECT 966.500000 330.350000 999.500000 331.650000 ;
      RECT 957.500000 330.350000 958.500000 331.650000 ;
      RECT 916.500000 330.350000 949.500000 331.650000 ;
      RECT 907.500000 330.350000 908.500000 331.650000 ;
      RECT 866.500000 330.350000 899.500000 331.650000 ;
      RECT 857.500000 330.350000 858.500000 331.650000 ;
      RECT 816.500000 330.350000 849.500000 331.650000 ;
      RECT 807.500000 330.350000 808.500000 331.650000 ;
      RECT 766.500000 330.350000 799.500000 331.650000 ;
      RECT 757.500000 330.350000 758.500000 331.650000 ;
      RECT 716.500000 330.350000 749.500000 331.650000 ;
      RECT 707.500000 330.350000 708.500000 331.650000 ;
      RECT 666.500000 330.350000 699.500000 331.650000 ;
      RECT 657.500000 330.350000 658.500000 331.650000 ;
      RECT 616.500000 330.350000 649.500000 331.650000 ;
      RECT 607.500000 330.350000 608.500000 331.650000 ;
      RECT 566.500000 330.350000 599.500000 331.650000 ;
      RECT 557.500000 330.350000 558.500000 331.650000 ;
      RECT 516.500000 330.350000 549.500000 331.650000 ;
      RECT 507.500000 330.350000 508.500000 331.650000 ;
      RECT 466.500000 330.350000 499.500000 331.650000 ;
      RECT 457.500000 330.350000 458.500000 331.650000 ;
      RECT 416.500000 330.350000 449.500000 331.650000 ;
      RECT 407.500000 330.350000 408.500000 331.650000 ;
      RECT 366.500000 330.350000 399.500000 331.650000 ;
      RECT 357.500000 330.350000 358.500000 331.650000 ;
      RECT 316.500000 330.350000 349.500000 331.650000 ;
      RECT 307.500000 330.350000 308.500000 331.650000 ;
      RECT 266.500000 330.350000 299.500000 331.650000 ;
      RECT 257.500000 330.350000 258.500000 331.650000 ;
      RECT 216.500000 330.350000 249.500000 331.650000 ;
      RECT 207.500000 330.350000 208.500000 331.650000 ;
      RECT 166.500000 330.350000 199.500000 331.650000 ;
      RECT 157.500000 330.350000 158.500000 331.650000 ;
      RECT 116.500000 330.350000 149.500000 331.650000 ;
      RECT 107.500000 330.350000 108.500000 331.650000 ;
      RECT 66.500000 330.350000 99.500000 331.650000 ;
      RECT 57.500000 330.350000 58.500000 331.650000 ;
      RECT 29.500000 330.350000 49.500000 331.650000 ;
      RECT 15.500000 330.350000 16.500000 331.650000 ;
      RECT 1157.500000 329.650000 1170.500000 330.350000 ;
      RECT 1107.500000 329.650000 1149.500000 330.350000 ;
      RECT 1057.500000 329.650000 1099.500000 330.350000 ;
      RECT 1007.500000 329.650000 1049.500000 330.350000 ;
      RECT 957.500000 329.650000 999.500000 330.350000 ;
      RECT 907.500000 329.650000 949.500000 330.350000 ;
      RECT 857.500000 329.650000 899.500000 330.350000 ;
      RECT 807.500000 329.650000 849.500000 330.350000 ;
      RECT 757.500000 329.650000 799.500000 330.350000 ;
      RECT 707.500000 329.650000 749.500000 330.350000 ;
      RECT 657.500000 329.650000 699.500000 330.350000 ;
      RECT 607.500000 329.650000 649.500000 330.350000 ;
      RECT 557.500000 329.650000 599.500000 330.350000 ;
      RECT 507.500000 329.650000 549.500000 330.350000 ;
      RECT 457.500000 329.650000 499.500000 330.350000 ;
      RECT 407.500000 329.650000 449.500000 330.350000 ;
      RECT 357.500000 329.650000 399.500000 330.350000 ;
      RECT 307.500000 329.650000 349.500000 330.350000 ;
      RECT 257.500000 329.650000 299.500000 330.350000 ;
      RECT 207.500000 329.650000 249.500000 330.350000 ;
      RECT 157.500000 329.650000 199.500000 330.350000 ;
      RECT 107.500000 329.650000 149.500000 330.350000 ;
      RECT 57.500000 329.650000 99.500000 330.350000 ;
      RECT 15.500000 329.650000 49.500000 330.350000 ;
      RECT 1183.500000 328.350000 1186.000000 331.650000 ;
      RECT 1169.500000 328.350000 1170.500000 329.650000 ;
      RECT 1116.500000 328.350000 1149.500000 329.650000 ;
      RECT 1107.500000 328.350000 1108.500000 329.650000 ;
      RECT 1066.500000 328.350000 1099.500000 329.650000 ;
      RECT 1057.500000 328.350000 1058.500000 329.650000 ;
      RECT 1016.500000 328.350000 1049.500000 329.650000 ;
      RECT 1007.500000 328.350000 1008.500000 329.650000 ;
      RECT 966.500000 328.350000 999.500000 329.650000 ;
      RECT 957.500000 328.350000 958.500000 329.650000 ;
      RECT 916.500000 328.350000 949.500000 329.650000 ;
      RECT 907.500000 328.350000 908.500000 329.650000 ;
      RECT 866.500000 328.350000 899.500000 329.650000 ;
      RECT 857.500000 328.350000 858.500000 329.650000 ;
      RECT 816.500000 328.350000 849.500000 329.650000 ;
      RECT 807.500000 328.350000 808.500000 329.650000 ;
      RECT 766.500000 328.350000 799.500000 329.650000 ;
      RECT 757.500000 328.350000 758.500000 329.650000 ;
      RECT 716.500000 328.350000 749.500000 329.650000 ;
      RECT 707.500000 328.350000 708.500000 329.650000 ;
      RECT 666.500000 328.350000 699.500000 329.650000 ;
      RECT 657.500000 328.350000 658.500000 329.650000 ;
      RECT 616.500000 328.350000 649.500000 329.650000 ;
      RECT 607.500000 328.350000 608.500000 329.650000 ;
      RECT 566.500000 328.350000 599.500000 329.650000 ;
      RECT 557.500000 328.350000 558.500000 329.650000 ;
      RECT 516.500000 328.350000 549.500000 329.650000 ;
      RECT 507.500000 328.350000 508.500000 329.650000 ;
      RECT 466.500000 328.350000 499.500000 329.650000 ;
      RECT 457.500000 328.350000 458.500000 329.650000 ;
      RECT 416.500000 328.350000 449.500000 329.650000 ;
      RECT 407.500000 328.350000 408.500000 329.650000 ;
      RECT 366.500000 328.350000 399.500000 329.650000 ;
      RECT 357.500000 328.350000 358.500000 329.650000 ;
      RECT 316.500000 328.350000 349.500000 329.650000 ;
      RECT 307.500000 328.350000 308.500000 329.650000 ;
      RECT 266.500000 328.350000 299.500000 329.650000 ;
      RECT 257.500000 328.350000 258.500000 329.650000 ;
      RECT 216.500000 328.350000 249.500000 329.650000 ;
      RECT 207.500000 328.350000 208.500000 329.650000 ;
      RECT 166.500000 328.350000 199.500000 329.650000 ;
      RECT 157.500000 328.350000 158.500000 329.650000 ;
      RECT 116.500000 328.350000 149.500000 329.650000 ;
      RECT 107.500000 328.350000 108.500000 329.650000 ;
      RECT 66.500000 328.350000 99.500000 329.650000 ;
      RECT 57.500000 328.350000 58.500000 329.650000 ;
      RECT 29.500000 328.350000 49.500000 329.650000 ;
      RECT 15.500000 328.350000 16.500000 329.650000 ;
      RECT 0.000000 328.350000 2.500000 331.650000 ;
      RECT 1169.500000 327.650000 1186.000000 328.350000 ;
      RECT 1116.500000 327.650000 1156.500000 328.350000 ;
      RECT 1066.500000 327.650000 1108.500000 328.350000 ;
      RECT 1016.500000 327.650000 1058.500000 328.350000 ;
      RECT 966.500000 327.650000 1008.500000 328.350000 ;
      RECT 916.500000 327.650000 958.500000 328.350000 ;
      RECT 866.500000 327.650000 908.500000 328.350000 ;
      RECT 816.500000 327.650000 858.500000 328.350000 ;
      RECT 766.500000 327.650000 808.500000 328.350000 ;
      RECT 716.500000 327.650000 758.500000 328.350000 ;
      RECT 666.500000 327.650000 708.500000 328.350000 ;
      RECT 616.500000 327.650000 658.500000 328.350000 ;
      RECT 566.500000 327.650000 608.500000 328.350000 ;
      RECT 516.500000 327.650000 558.500000 328.350000 ;
      RECT 466.500000 327.650000 508.500000 328.350000 ;
      RECT 416.500000 327.650000 458.500000 328.350000 ;
      RECT 366.500000 327.650000 408.500000 328.350000 ;
      RECT 316.500000 327.650000 358.500000 328.350000 ;
      RECT 266.500000 327.650000 308.500000 328.350000 ;
      RECT 216.500000 327.650000 258.500000 328.350000 ;
      RECT 166.500000 327.650000 208.500000 328.350000 ;
      RECT 116.500000 327.650000 158.500000 328.350000 ;
      RECT 66.500000 327.650000 108.500000 328.350000 ;
      RECT 29.500000 327.650000 58.500000 328.350000 ;
      RECT 0.000000 327.650000 16.500000 328.350000 ;
      RECT 1169.500000 326.350000 1170.500000 327.650000 ;
      RECT 1116.500000 326.350000 1149.500000 327.650000 ;
      RECT 1107.500000 326.350000 1108.500000 327.650000 ;
      RECT 1066.500000 326.350000 1099.500000 327.650000 ;
      RECT 1057.500000 326.350000 1058.500000 327.650000 ;
      RECT 1016.500000 326.350000 1049.500000 327.650000 ;
      RECT 1007.500000 326.350000 1008.500000 327.650000 ;
      RECT 966.500000 326.350000 999.500000 327.650000 ;
      RECT 957.500000 326.350000 958.500000 327.650000 ;
      RECT 916.500000 326.350000 949.500000 327.650000 ;
      RECT 907.500000 326.350000 908.500000 327.650000 ;
      RECT 866.500000 326.350000 899.500000 327.650000 ;
      RECT 857.500000 326.350000 858.500000 327.650000 ;
      RECT 816.500000 326.350000 849.500000 327.650000 ;
      RECT 807.500000 326.350000 808.500000 327.650000 ;
      RECT 766.500000 326.350000 799.500000 327.650000 ;
      RECT 757.500000 326.350000 758.500000 327.650000 ;
      RECT 716.500000 326.350000 749.500000 327.650000 ;
      RECT 707.500000 326.350000 708.500000 327.650000 ;
      RECT 666.500000 326.350000 699.500000 327.650000 ;
      RECT 657.500000 326.350000 658.500000 327.650000 ;
      RECT 616.500000 326.350000 649.500000 327.650000 ;
      RECT 607.500000 326.350000 608.500000 327.650000 ;
      RECT 566.500000 326.350000 599.500000 327.650000 ;
      RECT 557.500000 326.350000 558.500000 327.650000 ;
      RECT 516.500000 326.350000 549.500000 327.650000 ;
      RECT 507.500000 326.350000 508.500000 327.650000 ;
      RECT 466.500000 326.350000 499.500000 327.650000 ;
      RECT 457.500000 326.350000 458.500000 327.650000 ;
      RECT 416.500000 326.350000 449.500000 327.650000 ;
      RECT 407.500000 326.350000 408.500000 327.650000 ;
      RECT 366.500000 326.350000 399.500000 327.650000 ;
      RECT 357.500000 326.350000 358.500000 327.650000 ;
      RECT 316.500000 326.350000 349.500000 327.650000 ;
      RECT 307.500000 326.350000 308.500000 327.650000 ;
      RECT 266.500000 326.350000 299.500000 327.650000 ;
      RECT 257.500000 326.350000 258.500000 327.650000 ;
      RECT 216.500000 326.350000 249.500000 327.650000 ;
      RECT 207.500000 326.350000 208.500000 327.650000 ;
      RECT 166.500000 326.350000 199.500000 327.650000 ;
      RECT 157.500000 326.350000 158.500000 327.650000 ;
      RECT 116.500000 326.350000 149.500000 327.650000 ;
      RECT 107.500000 326.350000 108.500000 327.650000 ;
      RECT 66.500000 326.350000 99.500000 327.650000 ;
      RECT 57.500000 326.350000 58.500000 327.650000 ;
      RECT 29.500000 326.350000 49.500000 327.650000 ;
      RECT 15.500000 326.350000 16.500000 327.650000 ;
      RECT 1157.500000 325.650000 1170.500000 326.350000 ;
      RECT 1107.500000 325.650000 1149.500000 326.350000 ;
      RECT 1057.500000 325.650000 1099.500000 326.350000 ;
      RECT 1007.500000 325.650000 1049.500000 326.350000 ;
      RECT 957.500000 325.650000 999.500000 326.350000 ;
      RECT 907.500000 325.650000 949.500000 326.350000 ;
      RECT 857.500000 325.650000 899.500000 326.350000 ;
      RECT 807.500000 325.650000 849.500000 326.350000 ;
      RECT 757.500000 325.650000 799.500000 326.350000 ;
      RECT 707.500000 325.650000 749.500000 326.350000 ;
      RECT 657.500000 325.650000 699.500000 326.350000 ;
      RECT 607.500000 325.650000 649.500000 326.350000 ;
      RECT 557.500000 325.650000 599.500000 326.350000 ;
      RECT 507.500000 325.650000 549.500000 326.350000 ;
      RECT 457.500000 325.650000 499.500000 326.350000 ;
      RECT 407.500000 325.650000 449.500000 326.350000 ;
      RECT 357.500000 325.650000 399.500000 326.350000 ;
      RECT 307.500000 325.650000 349.500000 326.350000 ;
      RECT 257.500000 325.650000 299.500000 326.350000 ;
      RECT 207.500000 325.650000 249.500000 326.350000 ;
      RECT 157.500000 325.650000 199.500000 326.350000 ;
      RECT 107.500000 325.650000 149.500000 326.350000 ;
      RECT 57.500000 325.650000 99.500000 326.350000 ;
      RECT 15.500000 325.650000 49.500000 326.350000 ;
      RECT 1183.500000 324.350000 1186.000000 327.650000 ;
      RECT 1169.500000 324.350000 1170.500000 325.650000 ;
      RECT 1116.500000 324.350000 1149.500000 325.650000 ;
      RECT 1107.500000 324.350000 1108.500000 325.650000 ;
      RECT 1066.500000 324.350000 1099.500000 325.650000 ;
      RECT 1057.500000 324.350000 1058.500000 325.650000 ;
      RECT 1016.500000 324.350000 1049.500000 325.650000 ;
      RECT 1007.500000 324.350000 1008.500000 325.650000 ;
      RECT 966.500000 324.350000 999.500000 325.650000 ;
      RECT 957.500000 324.350000 958.500000 325.650000 ;
      RECT 916.500000 324.350000 949.500000 325.650000 ;
      RECT 907.500000 324.350000 908.500000 325.650000 ;
      RECT 866.500000 324.350000 899.500000 325.650000 ;
      RECT 857.500000 324.350000 858.500000 325.650000 ;
      RECT 816.500000 324.350000 849.500000 325.650000 ;
      RECT 807.500000 324.350000 808.500000 325.650000 ;
      RECT 766.500000 324.350000 799.500000 325.650000 ;
      RECT 757.500000 324.350000 758.500000 325.650000 ;
      RECT 716.500000 324.350000 749.500000 325.650000 ;
      RECT 707.500000 324.350000 708.500000 325.650000 ;
      RECT 666.500000 324.350000 699.500000 325.650000 ;
      RECT 657.500000 324.350000 658.500000 325.650000 ;
      RECT 616.500000 324.350000 649.500000 325.650000 ;
      RECT 607.500000 324.350000 608.500000 325.650000 ;
      RECT 566.500000 324.350000 599.500000 325.650000 ;
      RECT 557.500000 324.350000 558.500000 325.650000 ;
      RECT 516.500000 324.350000 549.500000 325.650000 ;
      RECT 507.500000 324.350000 508.500000 325.650000 ;
      RECT 466.500000 324.350000 499.500000 325.650000 ;
      RECT 457.500000 324.350000 458.500000 325.650000 ;
      RECT 416.500000 324.350000 449.500000 325.650000 ;
      RECT 407.500000 324.350000 408.500000 325.650000 ;
      RECT 366.500000 324.350000 399.500000 325.650000 ;
      RECT 357.500000 324.350000 358.500000 325.650000 ;
      RECT 316.500000 324.350000 349.500000 325.650000 ;
      RECT 307.500000 324.350000 308.500000 325.650000 ;
      RECT 266.500000 324.350000 299.500000 325.650000 ;
      RECT 257.500000 324.350000 258.500000 325.650000 ;
      RECT 216.500000 324.350000 249.500000 325.650000 ;
      RECT 207.500000 324.350000 208.500000 325.650000 ;
      RECT 166.500000 324.350000 199.500000 325.650000 ;
      RECT 157.500000 324.350000 158.500000 325.650000 ;
      RECT 116.500000 324.350000 149.500000 325.650000 ;
      RECT 107.500000 324.350000 108.500000 325.650000 ;
      RECT 66.500000 324.350000 99.500000 325.650000 ;
      RECT 57.500000 324.350000 58.500000 325.650000 ;
      RECT 29.500000 324.350000 49.500000 325.650000 ;
      RECT 15.500000 324.350000 16.500000 325.650000 ;
      RECT 0.000000 324.350000 2.500000 327.650000 ;
      RECT 1169.500000 323.650000 1186.000000 324.350000 ;
      RECT 1116.500000 323.650000 1156.500000 324.350000 ;
      RECT 1066.500000 323.650000 1108.500000 324.350000 ;
      RECT 1016.500000 323.650000 1058.500000 324.350000 ;
      RECT 966.500000 323.650000 1008.500000 324.350000 ;
      RECT 916.500000 323.650000 958.500000 324.350000 ;
      RECT 866.500000 323.650000 908.500000 324.350000 ;
      RECT 816.500000 323.650000 858.500000 324.350000 ;
      RECT 766.500000 323.650000 808.500000 324.350000 ;
      RECT 716.500000 323.650000 758.500000 324.350000 ;
      RECT 666.500000 323.650000 708.500000 324.350000 ;
      RECT 616.500000 323.650000 658.500000 324.350000 ;
      RECT 566.500000 323.650000 608.500000 324.350000 ;
      RECT 516.500000 323.650000 558.500000 324.350000 ;
      RECT 466.500000 323.650000 508.500000 324.350000 ;
      RECT 416.500000 323.650000 458.500000 324.350000 ;
      RECT 366.500000 323.650000 408.500000 324.350000 ;
      RECT 316.500000 323.650000 358.500000 324.350000 ;
      RECT 266.500000 323.650000 308.500000 324.350000 ;
      RECT 216.500000 323.650000 258.500000 324.350000 ;
      RECT 166.500000 323.650000 208.500000 324.350000 ;
      RECT 116.500000 323.650000 158.500000 324.350000 ;
      RECT 66.500000 323.650000 108.500000 324.350000 ;
      RECT 29.500000 323.650000 58.500000 324.350000 ;
      RECT 0.000000 323.650000 16.500000 324.350000 ;
      RECT 1169.500000 322.350000 1170.500000 323.650000 ;
      RECT 1116.500000 322.350000 1149.500000 323.650000 ;
      RECT 1107.500000 322.350000 1108.500000 323.650000 ;
      RECT 1066.500000 322.350000 1099.500000 323.650000 ;
      RECT 1057.500000 322.350000 1058.500000 323.650000 ;
      RECT 1016.500000 322.350000 1049.500000 323.650000 ;
      RECT 1007.500000 322.350000 1008.500000 323.650000 ;
      RECT 966.500000 322.350000 999.500000 323.650000 ;
      RECT 957.500000 322.350000 958.500000 323.650000 ;
      RECT 916.500000 322.350000 949.500000 323.650000 ;
      RECT 907.500000 322.350000 908.500000 323.650000 ;
      RECT 866.500000 322.350000 899.500000 323.650000 ;
      RECT 857.500000 322.350000 858.500000 323.650000 ;
      RECT 816.500000 322.350000 849.500000 323.650000 ;
      RECT 807.500000 322.350000 808.500000 323.650000 ;
      RECT 766.500000 322.350000 799.500000 323.650000 ;
      RECT 757.500000 322.350000 758.500000 323.650000 ;
      RECT 716.500000 322.350000 749.500000 323.650000 ;
      RECT 707.500000 322.350000 708.500000 323.650000 ;
      RECT 666.500000 322.350000 699.500000 323.650000 ;
      RECT 657.500000 322.350000 658.500000 323.650000 ;
      RECT 616.500000 322.350000 649.500000 323.650000 ;
      RECT 607.500000 322.350000 608.500000 323.650000 ;
      RECT 566.500000 322.350000 599.500000 323.650000 ;
      RECT 557.500000 322.350000 558.500000 323.650000 ;
      RECT 516.500000 322.350000 549.500000 323.650000 ;
      RECT 507.500000 322.350000 508.500000 323.650000 ;
      RECT 466.500000 322.350000 499.500000 323.650000 ;
      RECT 457.500000 322.350000 458.500000 323.650000 ;
      RECT 416.500000 322.350000 449.500000 323.650000 ;
      RECT 407.500000 322.350000 408.500000 323.650000 ;
      RECT 366.500000 322.350000 399.500000 323.650000 ;
      RECT 357.500000 322.350000 358.500000 323.650000 ;
      RECT 316.500000 322.350000 349.500000 323.650000 ;
      RECT 307.500000 322.350000 308.500000 323.650000 ;
      RECT 266.500000 322.350000 299.500000 323.650000 ;
      RECT 257.500000 322.350000 258.500000 323.650000 ;
      RECT 216.500000 322.350000 249.500000 323.650000 ;
      RECT 207.500000 322.350000 208.500000 323.650000 ;
      RECT 166.500000 322.350000 199.500000 323.650000 ;
      RECT 157.500000 322.350000 158.500000 323.650000 ;
      RECT 116.500000 322.350000 149.500000 323.650000 ;
      RECT 107.500000 322.350000 108.500000 323.650000 ;
      RECT 66.500000 322.350000 99.500000 323.650000 ;
      RECT 57.500000 322.350000 58.500000 323.650000 ;
      RECT 29.500000 322.350000 49.500000 323.650000 ;
      RECT 15.500000 322.350000 16.500000 323.650000 ;
      RECT 1157.500000 321.650000 1170.500000 322.350000 ;
      RECT 1107.500000 321.650000 1149.500000 322.350000 ;
      RECT 1057.500000 321.650000 1099.500000 322.350000 ;
      RECT 1007.500000 321.650000 1049.500000 322.350000 ;
      RECT 957.500000 321.650000 999.500000 322.350000 ;
      RECT 907.500000 321.650000 949.500000 322.350000 ;
      RECT 857.500000 321.650000 899.500000 322.350000 ;
      RECT 807.500000 321.650000 849.500000 322.350000 ;
      RECT 757.500000 321.650000 799.500000 322.350000 ;
      RECT 707.500000 321.650000 749.500000 322.350000 ;
      RECT 657.500000 321.650000 699.500000 322.350000 ;
      RECT 607.500000 321.650000 649.500000 322.350000 ;
      RECT 557.500000 321.650000 599.500000 322.350000 ;
      RECT 507.500000 321.650000 549.500000 322.350000 ;
      RECT 457.500000 321.650000 499.500000 322.350000 ;
      RECT 407.500000 321.650000 449.500000 322.350000 ;
      RECT 357.500000 321.650000 399.500000 322.350000 ;
      RECT 307.500000 321.650000 349.500000 322.350000 ;
      RECT 257.500000 321.650000 299.500000 322.350000 ;
      RECT 207.500000 321.650000 249.500000 322.350000 ;
      RECT 157.500000 321.650000 199.500000 322.350000 ;
      RECT 107.500000 321.650000 149.500000 322.350000 ;
      RECT 57.500000 321.650000 99.500000 322.350000 ;
      RECT 15.500000 321.650000 49.500000 322.350000 ;
      RECT 1183.500000 320.350000 1186.000000 323.650000 ;
      RECT 1169.500000 320.350000 1170.500000 321.650000 ;
      RECT 1116.500000 320.350000 1149.500000 321.650000 ;
      RECT 1107.500000 320.350000 1108.500000 321.650000 ;
      RECT 1066.500000 320.350000 1099.500000 321.650000 ;
      RECT 1057.500000 320.350000 1058.500000 321.650000 ;
      RECT 1016.500000 320.350000 1049.500000 321.650000 ;
      RECT 1007.500000 320.350000 1008.500000 321.650000 ;
      RECT 966.500000 320.350000 999.500000 321.650000 ;
      RECT 957.500000 320.350000 958.500000 321.650000 ;
      RECT 916.500000 320.350000 949.500000 321.650000 ;
      RECT 907.500000 320.350000 908.500000 321.650000 ;
      RECT 866.500000 320.350000 899.500000 321.650000 ;
      RECT 857.500000 320.350000 858.500000 321.650000 ;
      RECT 816.500000 320.350000 849.500000 321.650000 ;
      RECT 807.500000 320.350000 808.500000 321.650000 ;
      RECT 766.500000 320.350000 799.500000 321.650000 ;
      RECT 757.500000 320.350000 758.500000 321.650000 ;
      RECT 716.500000 320.350000 749.500000 321.650000 ;
      RECT 707.500000 320.350000 708.500000 321.650000 ;
      RECT 666.500000 320.350000 699.500000 321.650000 ;
      RECT 657.500000 320.350000 658.500000 321.650000 ;
      RECT 616.500000 320.350000 649.500000 321.650000 ;
      RECT 607.500000 320.350000 608.500000 321.650000 ;
      RECT 566.500000 320.350000 599.500000 321.650000 ;
      RECT 557.500000 320.350000 558.500000 321.650000 ;
      RECT 516.500000 320.350000 549.500000 321.650000 ;
      RECT 507.500000 320.350000 508.500000 321.650000 ;
      RECT 466.500000 320.350000 499.500000 321.650000 ;
      RECT 457.500000 320.350000 458.500000 321.650000 ;
      RECT 416.500000 320.350000 449.500000 321.650000 ;
      RECT 407.500000 320.350000 408.500000 321.650000 ;
      RECT 366.500000 320.350000 399.500000 321.650000 ;
      RECT 357.500000 320.350000 358.500000 321.650000 ;
      RECT 316.500000 320.350000 349.500000 321.650000 ;
      RECT 307.500000 320.350000 308.500000 321.650000 ;
      RECT 266.500000 320.350000 299.500000 321.650000 ;
      RECT 257.500000 320.350000 258.500000 321.650000 ;
      RECT 216.500000 320.350000 249.500000 321.650000 ;
      RECT 207.500000 320.350000 208.500000 321.650000 ;
      RECT 166.500000 320.350000 199.500000 321.650000 ;
      RECT 157.500000 320.350000 158.500000 321.650000 ;
      RECT 116.500000 320.350000 149.500000 321.650000 ;
      RECT 107.500000 320.350000 108.500000 321.650000 ;
      RECT 66.500000 320.350000 99.500000 321.650000 ;
      RECT 57.500000 320.350000 58.500000 321.650000 ;
      RECT 29.500000 320.350000 49.500000 321.650000 ;
      RECT 15.500000 320.350000 16.500000 321.650000 ;
      RECT 0.000000 320.350000 2.500000 323.650000 ;
      RECT 1169.500000 319.650000 1186.000000 320.350000 ;
      RECT 1116.500000 319.650000 1156.500000 320.350000 ;
      RECT 1066.500000 319.650000 1108.500000 320.350000 ;
      RECT 1016.500000 319.650000 1058.500000 320.350000 ;
      RECT 966.500000 319.650000 1008.500000 320.350000 ;
      RECT 916.500000 319.650000 958.500000 320.350000 ;
      RECT 866.500000 319.650000 908.500000 320.350000 ;
      RECT 816.500000 319.650000 858.500000 320.350000 ;
      RECT 766.500000 319.650000 808.500000 320.350000 ;
      RECT 716.500000 319.650000 758.500000 320.350000 ;
      RECT 666.500000 319.650000 708.500000 320.350000 ;
      RECT 616.500000 319.650000 658.500000 320.350000 ;
      RECT 566.500000 319.650000 608.500000 320.350000 ;
      RECT 516.500000 319.650000 558.500000 320.350000 ;
      RECT 466.500000 319.650000 508.500000 320.350000 ;
      RECT 366.500000 319.650000 408.500000 320.350000 ;
      RECT 316.500000 319.650000 358.500000 320.350000 ;
      RECT 266.500000 319.650000 308.500000 320.350000 ;
      RECT 216.500000 319.650000 258.500000 320.350000 ;
      RECT 166.500000 319.650000 208.500000 320.350000 ;
      RECT 116.500000 319.650000 158.500000 320.350000 ;
      RECT 66.500000 319.650000 108.500000 320.350000 ;
      RECT 29.500000 319.650000 58.500000 320.350000 ;
      RECT 0.000000 319.650000 16.500000 320.350000 ;
      RECT 416.500000 318.605000 458.500000 320.350000 ;
      RECT 1169.500000 318.350000 1170.500000 319.650000 ;
      RECT 1116.500000 318.350000 1149.500000 319.650000 ;
      RECT 1107.500000 318.350000 1108.500000 319.650000 ;
      RECT 1066.500000 318.350000 1099.500000 319.650000 ;
      RECT 1057.500000 318.350000 1058.500000 319.650000 ;
      RECT 1016.500000 318.350000 1049.500000 319.650000 ;
      RECT 1007.500000 318.350000 1008.500000 319.650000 ;
      RECT 966.500000 318.350000 999.500000 319.650000 ;
      RECT 957.500000 318.350000 958.500000 319.650000 ;
      RECT 916.500000 318.350000 949.500000 319.650000 ;
      RECT 907.500000 318.350000 908.500000 319.650000 ;
      RECT 866.500000 318.350000 899.500000 319.650000 ;
      RECT 857.500000 318.350000 858.500000 319.650000 ;
      RECT 816.500000 318.350000 849.500000 319.650000 ;
      RECT 807.500000 318.350000 808.500000 319.650000 ;
      RECT 766.500000 318.350000 799.500000 319.650000 ;
      RECT 757.500000 318.350000 758.500000 319.650000 ;
      RECT 716.500000 318.350000 749.500000 319.650000 ;
      RECT 707.500000 318.350000 708.500000 319.650000 ;
      RECT 666.500000 318.350000 699.500000 319.650000 ;
      RECT 657.500000 318.350000 658.500000 319.650000 ;
      RECT 616.500000 318.350000 649.500000 319.650000 ;
      RECT 607.500000 318.350000 608.500000 319.650000 ;
      RECT 566.500000 318.350000 599.500000 319.650000 ;
      RECT 557.500000 318.350000 558.500000 319.650000 ;
      RECT 516.500000 318.350000 549.500000 319.650000 ;
      RECT 507.500000 318.350000 508.500000 319.650000 ;
      RECT 466.500000 318.350000 499.500000 319.650000 ;
      RECT 457.500000 318.350000 458.500000 318.605000 ;
      RECT 416.500000 318.350000 449.500000 318.605000 ;
      RECT 407.500000 318.350000 408.500000 319.650000 ;
      RECT 366.500000 318.350000 399.500000 319.650000 ;
      RECT 357.500000 318.350000 358.500000 319.650000 ;
      RECT 316.500000 318.350000 349.500000 319.650000 ;
      RECT 307.500000 318.350000 308.500000 319.650000 ;
      RECT 266.500000 318.350000 299.500000 319.650000 ;
      RECT 257.500000 318.350000 258.500000 319.650000 ;
      RECT 216.500000 318.350000 249.500000 319.650000 ;
      RECT 207.500000 318.350000 208.500000 319.650000 ;
      RECT 166.500000 318.350000 199.500000 319.650000 ;
      RECT 157.500000 318.350000 158.500000 319.650000 ;
      RECT 116.500000 318.350000 149.500000 319.650000 ;
      RECT 107.500000 318.350000 108.500000 319.650000 ;
      RECT 66.500000 318.350000 99.500000 319.650000 ;
      RECT 57.500000 318.350000 58.500000 319.650000 ;
      RECT 29.500000 318.350000 49.500000 319.650000 ;
      RECT 15.500000 318.350000 16.500000 319.650000 ;
      RECT 1157.500000 317.650000 1170.500000 318.350000 ;
      RECT 1107.500000 317.650000 1149.500000 318.350000 ;
      RECT 1057.500000 317.650000 1099.500000 318.350000 ;
      RECT 1007.500000 317.650000 1049.500000 318.350000 ;
      RECT 957.500000 317.650000 999.500000 318.350000 ;
      RECT 907.500000 317.650000 949.500000 318.350000 ;
      RECT 857.500000 317.650000 899.500000 318.350000 ;
      RECT 807.500000 317.650000 849.500000 318.350000 ;
      RECT 757.500000 317.650000 799.500000 318.350000 ;
      RECT 707.500000 317.650000 749.500000 318.350000 ;
      RECT 657.500000 317.650000 699.500000 318.350000 ;
      RECT 607.500000 317.650000 649.500000 318.350000 ;
      RECT 557.500000 317.650000 599.500000 318.350000 ;
      RECT 507.500000 317.650000 549.500000 318.350000 ;
      RECT 407.500000 317.650000 449.500000 318.350000 ;
      RECT 357.500000 317.650000 399.500000 318.350000 ;
      RECT 307.500000 317.650000 349.500000 318.350000 ;
      RECT 257.500000 317.650000 299.500000 318.350000 ;
      RECT 207.500000 317.650000 249.500000 318.350000 ;
      RECT 157.500000 317.650000 199.500000 318.350000 ;
      RECT 107.500000 317.650000 149.500000 318.350000 ;
      RECT 57.500000 317.650000 99.500000 318.350000 ;
      RECT 15.500000 317.650000 49.500000 318.350000 ;
      RECT 1183.500000 316.350000 1186.000000 319.650000 ;
      RECT 1169.500000 316.350000 1170.500000 317.650000 ;
      RECT 1116.500000 316.350000 1149.500000 317.650000 ;
      RECT 1107.500000 316.350000 1108.500000 317.650000 ;
      RECT 1066.500000 316.350000 1099.500000 317.650000 ;
      RECT 1057.500000 316.350000 1058.500000 317.650000 ;
      RECT 1016.500000 316.350000 1049.500000 317.650000 ;
      RECT 1007.500000 316.350000 1008.500000 317.650000 ;
      RECT 966.500000 316.350000 999.500000 317.650000 ;
      RECT 957.500000 316.350000 958.500000 317.650000 ;
      RECT 916.500000 316.350000 949.500000 317.650000 ;
      RECT 907.500000 316.350000 908.500000 317.650000 ;
      RECT 866.500000 316.350000 899.500000 317.650000 ;
      RECT 857.500000 316.350000 858.500000 317.650000 ;
      RECT 816.500000 316.350000 849.500000 317.650000 ;
      RECT 807.500000 316.350000 808.500000 317.650000 ;
      RECT 766.500000 316.350000 799.500000 317.650000 ;
      RECT 757.500000 316.350000 758.500000 317.650000 ;
      RECT 716.500000 316.350000 749.500000 317.650000 ;
      RECT 707.500000 316.350000 708.500000 317.650000 ;
      RECT 666.500000 316.350000 699.500000 317.650000 ;
      RECT 657.500000 316.350000 658.500000 317.650000 ;
      RECT 616.500000 316.350000 649.500000 317.650000 ;
      RECT 607.500000 316.350000 608.500000 317.650000 ;
      RECT 566.500000 316.350000 599.500000 317.650000 ;
      RECT 557.500000 316.350000 558.500000 317.650000 ;
      RECT 516.500000 316.350000 549.500000 317.650000 ;
      RECT 507.500000 316.350000 508.500000 317.650000 ;
      RECT 457.500000 316.350000 499.500000 318.350000 ;
      RECT 407.500000 316.350000 408.500000 317.650000 ;
      RECT 366.500000 316.350000 399.500000 317.650000 ;
      RECT 357.500000 316.350000 358.500000 317.650000 ;
      RECT 316.500000 316.350000 349.500000 317.650000 ;
      RECT 307.500000 316.350000 308.500000 317.650000 ;
      RECT 266.500000 316.350000 299.500000 317.650000 ;
      RECT 257.500000 316.350000 258.500000 317.650000 ;
      RECT 216.500000 316.350000 249.500000 317.650000 ;
      RECT 207.500000 316.350000 208.500000 317.650000 ;
      RECT 166.500000 316.350000 199.500000 317.650000 ;
      RECT 157.500000 316.350000 158.500000 317.650000 ;
      RECT 116.500000 316.350000 149.500000 317.650000 ;
      RECT 107.500000 316.350000 108.500000 317.650000 ;
      RECT 66.500000 316.350000 99.500000 317.650000 ;
      RECT 57.500000 316.350000 58.500000 317.650000 ;
      RECT 29.500000 316.350000 49.500000 317.650000 ;
      RECT 15.500000 316.350000 16.500000 317.650000 ;
      RECT 0.000000 316.350000 2.500000 319.650000 ;
      RECT 1169.500000 315.650000 1186.000000 316.350000 ;
      RECT 1116.500000 315.650000 1156.500000 316.350000 ;
      RECT 1066.500000 315.650000 1108.500000 316.350000 ;
      RECT 1016.500000 315.650000 1058.500000 316.350000 ;
      RECT 966.500000 315.650000 1008.500000 316.350000 ;
      RECT 916.500000 315.650000 958.500000 316.350000 ;
      RECT 866.500000 315.650000 908.500000 316.350000 ;
      RECT 816.500000 315.650000 858.500000 316.350000 ;
      RECT 766.500000 315.650000 808.500000 316.350000 ;
      RECT 716.500000 315.650000 758.500000 316.350000 ;
      RECT 666.500000 315.650000 708.500000 316.350000 ;
      RECT 616.500000 315.650000 658.500000 316.350000 ;
      RECT 566.500000 315.650000 608.500000 316.350000 ;
      RECT 516.500000 315.650000 558.500000 316.350000 ;
      RECT 457.500000 315.650000 508.500000 316.350000 ;
      RECT 366.500000 315.650000 408.500000 316.350000 ;
      RECT 316.500000 315.650000 358.500000 316.350000 ;
      RECT 266.500000 315.650000 308.500000 316.350000 ;
      RECT 216.500000 315.650000 258.500000 316.350000 ;
      RECT 166.500000 315.650000 208.500000 316.350000 ;
      RECT 116.500000 315.650000 158.500000 316.350000 ;
      RECT 66.500000 315.650000 108.500000 316.350000 ;
      RECT 29.500000 315.650000 58.500000 316.350000 ;
      RECT 0.000000 315.650000 16.500000 316.350000 ;
      RECT 457.500000 314.605000 499.500000 315.650000 ;
      RECT 416.500000 314.605000 449.500000 317.650000 ;
      RECT 1169.500000 314.350000 1170.500000 315.650000 ;
      RECT 1116.500000 314.350000 1149.500000 315.650000 ;
      RECT 1107.500000 314.350000 1108.500000 315.650000 ;
      RECT 1066.500000 314.350000 1099.500000 315.650000 ;
      RECT 1057.500000 314.350000 1058.500000 315.650000 ;
      RECT 1016.500000 314.350000 1049.500000 315.650000 ;
      RECT 1007.500000 314.350000 1008.500000 315.650000 ;
      RECT 966.500000 314.350000 999.500000 315.650000 ;
      RECT 957.500000 314.350000 958.500000 315.650000 ;
      RECT 916.500000 314.350000 949.500000 315.650000 ;
      RECT 907.500000 314.350000 908.500000 315.650000 ;
      RECT 866.500000 314.350000 899.500000 315.650000 ;
      RECT 857.500000 314.350000 858.500000 315.650000 ;
      RECT 816.500000 314.350000 849.500000 315.650000 ;
      RECT 807.500000 314.350000 808.500000 315.650000 ;
      RECT 766.500000 314.350000 799.500000 315.650000 ;
      RECT 757.500000 314.350000 758.500000 315.650000 ;
      RECT 716.500000 314.350000 749.500000 315.650000 ;
      RECT 707.500000 314.350000 708.500000 315.650000 ;
      RECT 666.500000 314.350000 699.500000 315.650000 ;
      RECT 657.500000 314.350000 658.500000 315.650000 ;
      RECT 616.500000 314.350000 649.500000 315.650000 ;
      RECT 607.500000 314.350000 608.500000 315.650000 ;
      RECT 566.500000 314.350000 599.500000 315.650000 ;
      RECT 557.500000 314.350000 558.500000 315.650000 ;
      RECT 516.500000 314.350000 549.500000 315.650000 ;
      RECT 507.500000 314.350000 508.500000 315.650000 ;
      RECT 416.500000 314.350000 499.500000 314.605000 ;
      RECT 407.500000 314.350000 408.500000 315.650000 ;
      RECT 366.500000 314.350000 399.500000 315.650000 ;
      RECT 357.500000 314.350000 358.500000 315.650000 ;
      RECT 316.500000 314.350000 349.500000 315.650000 ;
      RECT 307.500000 314.350000 308.500000 315.650000 ;
      RECT 266.500000 314.350000 299.500000 315.650000 ;
      RECT 257.500000 314.350000 258.500000 315.650000 ;
      RECT 216.500000 314.350000 249.500000 315.650000 ;
      RECT 207.500000 314.350000 208.500000 315.650000 ;
      RECT 166.500000 314.350000 199.500000 315.650000 ;
      RECT 157.500000 314.350000 158.500000 315.650000 ;
      RECT 116.500000 314.350000 149.500000 315.650000 ;
      RECT 107.500000 314.350000 108.500000 315.650000 ;
      RECT 66.500000 314.350000 99.500000 315.650000 ;
      RECT 57.500000 314.350000 58.500000 315.650000 ;
      RECT 29.500000 314.350000 49.500000 315.650000 ;
      RECT 15.500000 314.350000 16.500000 315.650000 ;
      RECT 1157.500000 313.650000 1170.500000 314.350000 ;
      RECT 1107.500000 313.650000 1149.500000 314.350000 ;
      RECT 1057.500000 313.650000 1099.500000 314.350000 ;
      RECT 1007.500000 313.650000 1049.500000 314.350000 ;
      RECT 957.500000 313.650000 999.500000 314.350000 ;
      RECT 907.500000 313.650000 949.500000 314.350000 ;
      RECT 857.500000 313.650000 899.500000 314.350000 ;
      RECT 807.500000 313.650000 849.500000 314.350000 ;
      RECT 757.500000 313.650000 799.500000 314.350000 ;
      RECT 707.500000 313.650000 749.500000 314.350000 ;
      RECT 657.500000 313.650000 699.500000 314.350000 ;
      RECT 607.500000 313.650000 649.500000 314.350000 ;
      RECT 557.500000 313.650000 599.500000 314.350000 ;
      RECT 507.500000 313.650000 549.500000 314.350000 ;
      RECT 407.500000 313.650000 499.500000 314.350000 ;
      RECT 357.500000 313.650000 399.500000 314.350000 ;
      RECT 307.500000 313.650000 349.500000 314.350000 ;
      RECT 257.500000 313.650000 299.500000 314.350000 ;
      RECT 207.500000 313.650000 249.500000 314.350000 ;
      RECT 157.500000 313.650000 199.500000 314.350000 ;
      RECT 107.500000 313.650000 149.500000 314.350000 ;
      RECT 57.500000 313.650000 99.500000 314.350000 ;
      RECT 15.500000 313.650000 49.500000 314.350000 ;
      RECT 1183.500000 312.350000 1186.000000 315.650000 ;
      RECT 1169.500000 312.350000 1170.500000 313.650000 ;
      RECT 1116.500000 312.350000 1149.500000 313.650000 ;
      RECT 1107.500000 312.350000 1108.500000 313.650000 ;
      RECT 1066.500000 312.350000 1099.500000 313.650000 ;
      RECT 1057.500000 312.350000 1058.500000 313.650000 ;
      RECT 1016.500000 312.350000 1049.500000 313.650000 ;
      RECT 1007.500000 312.350000 1008.500000 313.650000 ;
      RECT 966.500000 312.350000 999.500000 313.650000 ;
      RECT 957.500000 312.350000 958.500000 313.650000 ;
      RECT 916.500000 312.350000 949.500000 313.650000 ;
      RECT 907.500000 312.350000 908.500000 313.650000 ;
      RECT 866.500000 312.350000 899.500000 313.650000 ;
      RECT 857.500000 312.350000 858.500000 313.650000 ;
      RECT 816.500000 312.350000 849.500000 313.650000 ;
      RECT 807.500000 312.350000 808.500000 313.650000 ;
      RECT 766.500000 312.350000 799.500000 313.650000 ;
      RECT 757.500000 312.350000 758.500000 313.650000 ;
      RECT 716.500000 312.350000 749.500000 313.650000 ;
      RECT 707.500000 312.350000 708.500000 313.650000 ;
      RECT 666.500000 312.350000 699.500000 313.650000 ;
      RECT 657.500000 312.350000 658.500000 313.650000 ;
      RECT 616.500000 312.350000 649.500000 313.650000 ;
      RECT 607.500000 312.350000 608.500000 313.650000 ;
      RECT 566.500000 312.350000 599.500000 313.650000 ;
      RECT 557.500000 312.350000 558.500000 313.650000 ;
      RECT 516.500000 312.350000 549.500000 313.650000 ;
      RECT 507.500000 312.350000 508.500000 313.650000 ;
      RECT 416.500000 312.350000 499.500000 313.650000 ;
      RECT 407.500000 312.350000 408.500000 313.650000 ;
      RECT 366.500000 312.350000 399.500000 313.650000 ;
      RECT 357.500000 312.350000 358.500000 313.650000 ;
      RECT 316.500000 312.350000 349.500000 313.650000 ;
      RECT 307.500000 312.350000 308.500000 313.650000 ;
      RECT 266.500000 312.350000 299.500000 313.650000 ;
      RECT 257.500000 312.350000 258.500000 313.650000 ;
      RECT 216.500000 312.350000 249.500000 313.650000 ;
      RECT 207.500000 312.350000 208.500000 313.650000 ;
      RECT 166.500000 312.350000 199.500000 313.650000 ;
      RECT 157.500000 312.350000 158.500000 313.650000 ;
      RECT 116.500000 312.350000 149.500000 313.650000 ;
      RECT 107.500000 312.350000 108.500000 313.650000 ;
      RECT 66.500000 312.350000 99.500000 313.650000 ;
      RECT 57.500000 312.350000 58.500000 313.650000 ;
      RECT 29.500000 312.350000 49.500000 313.650000 ;
      RECT 15.500000 312.350000 16.500000 313.650000 ;
      RECT 0.000000 312.350000 2.500000 315.650000 ;
      RECT 1169.500000 311.650000 1186.000000 312.350000 ;
      RECT 1116.500000 311.650000 1156.500000 312.350000 ;
      RECT 1066.500000 311.650000 1108.500000 312.350000 ;
      RECT 1016.500000 311.650000 1058.500000 312.350000 ;
      RECT 966.500000 311.650000 1008.500000 312.350000 ;
      RECT 916.500000 311.650000 958.500000 312.350000 ;
      RECT 866.500000 311.650000 908.500000 312.350000 ;
      RECT 816.500000 311.650000 858.500000 312.350000 ;
      RECT 766.500000 311.650000 808.500000 312.350000 ;
      RECT 716.500000 311.650000 758.500000 312.350000 ;
      RECT 666.500000 311.650000 708.500000 312.350000 ;
      RECT 616.500000 311.650000 658.500000 312.350000 ;
      RECT 566.500000 311.650000 608.500000 312.350000 ;
      RECT 516.500000 311.650000 558.500000 312.350000 ;
      RECT 416.500000 311.650000 508.500000 312.350000 ;
      RECT 366.500000 311.650000 408.500000 312.350000 ;
      RECT 316.500000 311.650000 358.500000 312.350000 ;
      RECT 266.500000 311.650000 308.500000 312.350000 ;
      RECT 216.500000 311.650000 258.500000 312.350000 ;
      RECT 166.500000 311.650000 208.500000 312.350000 ;
      RECT 116.500000 311.650000 158.500000 312.350000 ;
      RECT 66.500000 311.650000 108.500000 312.350000 ;
      RECT 29.500000 311.650000 58.500000 312.350000 ;
      RECT 0.000000 311.650000 16.500000 312.350000 ;
      RECT 1169.500000 310.350000 1170.500000 311.650000 ;
      RECT 1116.500000 310.350000 1149.500000 311.650000 ;
      RECT 1107.500000 310.350000 1108.500000 311.650000 ;
      RECT 1066.500000 310.350000 1099.500000 311.650000 ;
      RECT 1057.500000 310.350000 1058.500000 311.650000 ;
      RECT 1016.500000 310.350000 1049.500000 311.650000 ;
      RECT 1007.500000 310.350000 1008.500000 311.650000 ;
      RECT 966.500000 310.350000 999.500000 311.650000 ;
      RECT 957.500000 310.350000 958.500000 311.650000 ;
      RECT 916.500000 310.350000 949.500000 311.650000 ;
      RECT 907.500000 310.350000 908.500000 311.650000 ;
      RECT 866.500000 310.350000 899.500000 311.650000 ;
      RECT 857.500000 310.350000 858.500000 311.650000 ;
      RECT 816.500000 310.350000 849.500000 311.650000 ;
      RECT 807.500000 310.350000 808.500000 311.650000 ;
      RECT 766.500000 310.350000 799.500000 311.650000 ;
      RECT 757.500000 310.350000 758.500000 311.650000 ;
      RECT 716.500000 310.350000 749.500000 311.650000 ;
      RECT 707.500000 310.350000 708.500000 311.650000 ;
      RECT 666.500000 310.350000 699.500000 311.650000 ;
      RECT 657.500000 310.350000 658.500000 311.650000 ;
      RECT 616.500000 310.350000 649.500000 311.650000 ;
      RECT 607.500000 310.350000 608.500000 311.650000 ;
      RECT 566.500000 310.350000 599.500000 311.650000 ;
      RECT 557.500000 310.350000 558.500000 311.650000 ;
      RECT 516.500000 310.350000 549.500000 311.650000 ;
      RECT 507.500000 310.350000 508.500000 311.650000 ;
      RECT 416.500000 310.350000 499.500000 311.650000 ;
      RECT 407.500000 310.350000 408.500000 311.650000 ;
      RECT 366.500000 310.350000 399.500000 311.650000 ;
      RECT 357.500000 310.350000 358.500000 311.650000 ;
      RECT 316.500000 310.350000 349.500000 311.650000 ;
      RECT 307.500000 310.350000 308.500000 311.650000 ;
      RECT 266.500000 310.350000 299.500000 311.650000 ;
      RECT 257.500000 310.350000 258.500000 311.650000 ;
      RECT 216.500000 310.350000 249.500000 311.650000 ;
      RECT 207.500000 310.350000 208.500000 311.650000 ;
      RECT 166.500000 310.350000 199.500000 311.650000 ;
      RECT 157.500000 310.350000 158.500000 311.650000 ;
      RECT 116.500000 310.350000 149.500000 311.650000 ;
      RECT 107.500000 310.350000 108.500000 311.650000 ;
      RECT 66.500000 310.350000 99.500000 311.650000 ;
      RECT 57.500000 310.350000 58.500000 311.650000 ;
      RECT 29.500000 310.350000 49.500000 311.650000 ;
      RECT 15.500000 310.350000 16.500000 311.650000 ;
      RECT 1157.500000 309.650000 1170.500000 310.350000 ;
      RECT 1107.500000 309.650000 1149.500000 310.350000 ;
      RECT 1057.500000 309.650000 1099.500000 310.350000 ;
      RECT 1007.500000 309.650000 1049.500000 310.350000 ;
      RECT 957.500000 309.650000 999.500000 310.350000 ;
      RECT 907.500000 309.650000 949.500000 310.350000 ;
      RECT 857.500000 309.650000 899.500000 310.350000 ;
      RECT 807.500000 309.650000 849.500000 310.350000 ;
      RECT 757.500000 309.650000 799.500000 310.350000 ;
      RECT 707.500000 309.650000 749.500000 310.350000 ;
      RECT 657.500000 309.650000 699.500000 310.350000 ;
      RECT 607.500000 309.650000 649.500000 310.350000 ;
      RECT 557.500000 309.650000 599.500000 310.350000 ;
      RECT 507.500000 309.650000 549.500000 310.350000 ;
      RECT 407.500000 309.650000 499.500000 310.350000 ;
      RECT 357.500000 309.650000 399.500000 310.350000 ;
      RECT 307.500000 309.650000 349.500000 310.350000 ;
      RECT 257.500000 309.650000 299.500000 310.350000 ;
      RECT 207.500000 309.650000 249.500000 310.350000 ;
      RECT 157.500000 309.650000 199.500000 310.350000 ;
      RECT 107.500000 309.650000 149.500000 310.350000 ;
      RECT 57.500000 309.650000 99.500000 310.350000 ;
      RECT 15.500000 309.650000 49.500000 310.350000 ;
      RECT 1183.500000 308.350000 1186.000000 311.650000 ;
      RECT 1169.500000 308.350000 1170.500000 309.650000 ;
      RECT 1116.500000 308.350000 1149.500000 309.650000 ;
      RECT 1107.500000 308.350000 1108.500000 309.650000 ;
      RECT 1066.500000 308.350000 1099.500000 309.650000 ;
      RECT 1057.500000 308.350000 1058.500000 309.650000 ;
      RECT 1016.500000 308.350000 1049.500000 309.650000 ;
      RECT 1007.500000 308.350000 1008.500000 309.650000 ;
      RECT 966.500000 308.350000 999.500000 309.650000 ;
      RECT 957.500000 308.350000 958.500000 309.650000 ;
      RECT 916.500000 308.350000 949.500000 309.650000 ;
      RECT 907.500000 308.350000 908.500000 309.650000 ;
      RECT 866.500000 308.350000 899.500000 309.650000 ;
      RECT 857.500000 308.350000 858.500000 309.650000 ;
      RECT 816.500000 308.350000 849.500000 309.650000 ;
      RECT 807.500000 308.350000 808.500000 309.650000 ;
      RECT 766.500000 308.350000 799.500000 309.650000 ;
      RECT 757.500000 308.350000 758.500000 309.650000 ;
      RECT 716.500000 308.350000 749.500000 309.650000 ;
      RECT 707.500000 308.350000 708.500000 309.650000 ;
      RECT 666.500000 308.350000 699.500000 309.650000 ;
      RECT 657.500000 308.350000 658.500000 309.650000 ;
      RECT 616.500000 308.350000 649.500000 309.650000 ;
      RECT 607.500000 308.350000 608.500000 309.650000 ;
      RECT 566.500000 308.350000 599.500000 309.650000 ;
      RECT 557.500000 308.350000 558.500000 309.650000 ;
      RECT 516.500000 308.350000 549.500000 309.650000 ;
      RECT 507.500000 308.350000 508.500000 309.650000 ;
      RECT 416.500000 308.350000 499.500000 309.650000 ;
      RECT 407.500000 308.350000 408.500000 309.650000 ;
      RECT 366.500000 308.350000 399.500000 309.650000 ;
      RECT 357.500000 308.350000 358.500000 309.650000 ;
      RECT 316.500000 308.350000 349.500000 309.650000 ;
      RECT 307.500000 308.350000 308.500000 309.650000 ;
      RECT 266.500000 308.350000 299.500000 309.650000 ;
      RECT 257.500000 308.350000 258.500000 309.650000 ;
      RECT 216.500000 308.350000 249.500000 309.650000 ;
      RECT 207.500000 308.350000 208.500000 309.650000 ;
      RECT 166.500000 308.350000 199.500000 309.650000 ;
      RECT 157.500000 308.350000 158.500000 309.650000 ;
      RECT 116.500000 308.350000 149.500000 309.650000 ;
      RECT 107.500000 308.350000 108.500000 309.650000 ;
      RECT 66.500000 308.350000 99.500000 309.650000 ;
      RECT 57.500000 308.350000 58.500000 309.650000 ;
      RECT 29.500000 308.350000 49.500000 309.650000 ;
      RECT 15.500000 308.350000 16.500000 309.650000 ;
      RECT 0.000000 308.350000 2.500000 311.650000 ;
      RECT 1169.500000 307.650000 1186.000000 308.350000 ;
      RECT 1116.500000 307.650000 1156.500000 308.350000 ;
      RECT 1066.500000 307.650000 1108.500000 308.350000 ;
      RECT 1016.500000 307.650000 1058.500000 308.350000 ;
      RECT 966.500000 307.650000 1008.500000 308.350000 ;
      RECT 916.500000 307.650000 958.500000 308.350000 ;
      RECT 866.500000 307.650000 908.500000 308.350000 ;
      RECT 816.500000 307.650000 858.500000 308.350000 ;
      RECT 766.500000 307.650000 808.500000 308.350000 ;
      RECT 716.500000 307.650000 758.500000 308.350000 ;
      RECT 666.500000 307.650000 708.500000 308.350000 ;
      RECT 616.500000 307.650000 658.500000 308.350000 ;
      RECT 566.500000 307.650000 608.500000 308.350000 ;
      RECT 516.500000 307.650000 558.500000 308.350000 ;
      RECT 416.500000 307.650000 508.500000 308.350000 ;
      RECT 366.500000 307.650000 408.500000 308.350000 ;
      RECT 316.500000 307.650000 358.500000 308.350000 ;
      RECT 266.500000 307.650000 308.500000 308.350000 ;
      RECT 216.500000 307.650000 258.500000 308.350000 ;
      RECT 166.500000 307.650000 208.500000 308.350000 ;
      RECT 116.500000 307.650000 158.500000 308.350000 ;
      RECT 66.500000 307.650000 108.500000 308.350000 ;
      RECT 29.500000 307.650000 58.500000 308.350000 ;
      RECT 0.000000 307.650000 16.500000 308.350000 ;
      RECT 1169.500000 306.350000 1170.500000 307.650000 ;
      RECT 1116.500000 306.350000 1149.500000 307.650000 ;
      RECT 1107.500000 306.350000 1108.500000 307.650000 ;
      RECT 1066.500000 306.350000 1099.500000 307.650000 ;
      RECT 1057.500000 306.350000 1058.500000 307.650000 ;
      RECT 1016.500000 306.350000 1049.500000 307.650000 ;
      RECT 1007.500000 306.350000 1008.500000 307.650000 ;
      RECT 966.500000 306.350000 999.500000 307.650000 ;
      RECT 957.500000 306.350000 958.500000 307.650000 ;
      RECT 916.500000 306.350000 949.500000 307.650000 ;
      RECT 907.500000 306.350000 908.500000 307.650000 ;
      RECT 866.500000 306.350000 899.500000 307.650000 ;
      RECT 857.500000 306.350000 858.500000 307.650000 ;
      RECT 816.500000 306.350000 849.500000 307.650000 ;
      RECT 807.500000 306.350000 808.500000 307.650000 ;
      RECT 766.500000 306.350000 799.500000 307.650000 ;
      RECT 757.500000 306.350000 758.500000 307.650000 ;
      RECT 716.500000 306.350000 749.500000 307.650000 ;
      RECT 707.500000 306.350000 708.500000 307.650000 ;
      RECT 666.500000 306.350000 699.500000 307.650000 ;
      RECT 657.500000 306.350000 658.500000 307.650000 ;
      RECT 616.500000 306.350000 649.500000 307.650000 ;
      RECT 607.500000 306.350000 608.500000 307.650000 ;
      RECT 566.500000 306.350000 599.500000 307.650000 ;
      RECT 557.500000 306.350000 558.500000 307.650000 ;
      RECT 516.500000 306.350000 549.500000 307.650000 ;
      RECT 507.500000 306.350000 508.500000 307.650000 ;
      RECT 416.500000 306.350000 499.500000 307.650000 ;
      RECT 407.500000 306.350000 408.500000 307.650000 ;
      RECT 366.500000 306.350000 399.500000 307.650000 ;
      RECT 357.500000 306.350000 358.500000 307.650000 ;
      RECT 316.500000 306.350000 349.500000 307.650000 ;
      RECT 307.500000 306.350000 308.500000 307.650000 ;
      RECT 266.500000 306.350000 299.500000 307.650000 ;
      RECT 257.500000 306.350000 258.500000 307.650000 ;
      RECT 216.500000 306.350000 249.500000 307.650000 ;
      RECT 207.500000 306.350000 208.500000 307.650000 ;
      RECT 166.500000 306.350000 199.500000 307.650000 ;
      RECT 157.500000 306.350000 158.500000 307.650000 ;
      RECT 116.500000 306.350000 149.500000 307.650000 ;
      RECT 107.500000 306.350000 108.500000 307.650000 ;
      RECT 66.500000 306.350000 99.500000 307.650000 ;
      RECT 57.500000 306.350000 58.500000 307.650000 ;
      RECT 29.500000 306.350000 49.500000 307.650000 ;
      RECT 15.500000 306.350000 16.500000 307.650000 ;
      RECT 1157.500000 305.650000 1170.500000 306.350000 ;
      RECT 1107.500000 305.650000 1149.500000 306.350000 ;
      RECT 1057.500000 305.650000 1099.500000 306.350000 ;
      RECT 1007.500000 305.650000 1049.500000 306.350000 ;
      RECT 957.500000 305.650000 999.500000 306.350000 ;
      RECT 907.500000 305.650000 949.500000 306.350000 ;
      RECT 857.500000 305.650000 899.500000 306.350000 ;
      RECT 807.500000 305.650000 849.500000 306.350000 ;
      RECT 757.500000 305.650000 799.500000 306.350000 ;
      RECT 707.500000 305.650000 749.500000 306.350000 ;
      RECT 657.500000 305.650000 699.500000 306.350000 ;
      RECT 607.500000 305.650000 649.500000 306.350000 ;
      RECT 557.500000 305.650000 599.500000 306.350000 ;
      RECT 507.500000 305.650000 549.500000 306.350000 ;
      RECT 407.500000 305.650000 499.500000 306.350000 ;
      RECT 357.500000 305.650000 399.500000 306.350000 ;
      RECT 307.500000 305.650000 349.500000 306.350000 ;
      RECT 257.500000 305.650000 299.500000 306.350000 ;
      RECT 207.500000 305.650000 249.500000 306.350000 ;
      RECT 157.500000 305.650000 199.500000 306.350000 ;
      RECT 107.500000 305.650000 149.500000 306.350000 ;
      RECT 57.500000 305.650000 99.500000 306.350000 ;
      RECT 15.500000 305.650000 49.500000 306.350000 ;
      RECT 1183.500000 304.350000 1186.000000 307.650000 ;
      RECT 1169.500000 304.350000 1170.500000 305.650000 ;
      RECT 1116.500000 304.350000 1149.500000 305.650000 ;
      RECT 1107.500000 304.350000 1108.500000 305.650000 ;
      RECT 1066.500000 304.350000 1099.500000 305.650000 ;
      RECT 1057.500000 304.350000 1058.500000 305.650000 ;
      RECT 1016.500000 304.350000 1049.500000 305.650000 ;
      RECT 1007.500000 304.350000 1008.500000 305.650000 ;
      RECT 966.500000 304.350000 999.500000 305.650000 ;
      RECT 957.500000 304.350000 958.500000 305.650000 ;
      RECT 916.500000 304.350000 949.500000 305.650000 ;
      RECT 907.500000 304.350000 908.500000 305.650000 ;
      RECT 866.500000 304.350000 899.500000 305.650000 ;
      RECT 857.500000 304.350000 858.500000 305.650000 ;
      RECT 816.500000 304.350000 849.500000 305.650000 ;
      RECT 807.500000 304.350000 808.500000 305.650000 ;
      RECT 766.500000 304.350000 799.500000 305.650000 ;
      RECT 757.500000 304.350000 758.500000 305.650000 ;
      RECT 716.500000 304.350000 749.500000 305.650000 ;
      RECT 707.500000 304.350000 708.500000 305.650000 ;
      RECT 666.500000 304.350000 699.500000 305.650000 ;
      RECT 657.500000 304.350000 658.500000 305.650000 ;
      RECT 616.500000 304.350000 649.500000 305.650000 ;
      RECT 607.500000 304.350000 608.500000 305.650000 ;
      RECT 566.500000 304.350000 599.500000 305.650000 ;
      RECT 557.500000 304.350000 558.500000 305.650000 ;
      RECT 516.500000 304.350000 549.500000 305.650000 ;
      RECT 507.500000 304.350000 508.500000 305.650000 ;
      RECT 416.500000 304.350000 499.500000 305.650000 ;
      RECT 407.500000 304.350000 408.500000 305.650000 ;
      RECT 366.500000 304.350000 399.500000 305.650000 ;
      RECT 357.500000 304.350000 358.500000 305.650000 ;
      RECT 316.500000 304.350000 349.500000 305.650000 ;
      RECT 307.500000 304.350000 308.500000 305.650000 ;
      RECT 266.500000 304.350000 299.500000 305.650000 ;
      RECT 257.500000 304.350000 258.500000 305.650000 ;
      RECT 216.500000 304.350000 249.500000 305.650000 ;
      RECT 207.500000 304.350000 208.500000 305.650000 ;
      RECT 166.500000 304.350000 199.500000 305.650000 ;
      RECT 157.500000 304.350000 158.500000 305.650000 ;
      RECT 116.500000 304.350000 149.500000 305.650000 ;
      RECT 107.500000 304.350000 108.500000 305.650000 ;
      RECT 66.500000 304.350000 99.500000 305.650000 ;
      RECT 57.500000 304.350000 58.500000 305.650000 ;
      RECT 29.500000 304.350000 49.500000 305.650000 ;
      RECT 15.500000 304.350000 16.500000 305.650000 ;
      RECT 0.000000 304.350000 2.500000 307.650000 ;
      RECT 416.500000 303.730000 508.500000 304.350000 ;
      RECT 1169.500000 303.650000 1186.000000 304.350000 ;
      RECT 1116.500000 303.650000 1156.500000 304.350000 ;
      RECT 1066.500000 303.650000 1108.500000 304.350000 ;
      RECT 1016.500000 303.650000 1058.500000 304.350000 ;
      RECT 966.500000 303.650000 1008.500000 304.350000 ;
      RECT 916.500000 303.650000 958.500000 304.350000 ;
      RECT 866.500000 303.650000 908.500000 304.350000 ;
      RECT 816.500000 303.650000 858.500000 304.350000 ;
      RECT 766.500000 303.650000 808.500000 304.350000 ;
      RECT 716.500000 303.650000 758.500000 304.350000 ;
      RECT 666.500000 303.650000 708.500000 304.350000 ;
      RECT 616.500000 303.650000 658.500000 304.350000 ;
      RECT 566.500000 303.650000 608.500000 304.350000 ;
      RECT 516.500000 303.650000 558.500000 304.350000 ;
      RECT 466.500000 303.650000 508.500000 303.730000 ;
      RECT 366.500000 303.650000 408.500000 304.350000 ;
      RECT 316.500000 303.650000 358.500000 304.350000 ;
      RECT 266.500000 303.650000 308.500000 304.350000 ;
      RECT 216.500000 303.650000 258.500000 304.350000 ;
      RECT 166.500000 303.650000 208.500000 304.350000 ;
      RECT 116.500000 303.650000 158.500000 304.350000 ;
      RECT 66.500000 303.650000 108.500000 304.350000 ;
      RECT 29.500000 303.650000 58.500000 304.350000 ;
      RECT 0.000000 303.650000 16.500000 304.350000 ;
      RECT 1169.500000 302.350000 1170.500000 303.650000 ;
      RECT 1116.500000 302.350000 1149.500000 303.650000 ;
      RECT 1107.500000 302.350000 1108.500000 303.650000 ;
      RECT 1066.500000 302.350000 1099.500000 303.650000 ;
      RECT 1057.500000 302.350000 1058.500000 303.650000 ;
      RECT 1016.500000 302.350000 1049.500000 303.650000 ;
      RECT 1007.500000 302.350000 1008.500000 303.650000 ;
      RECT 966.500000 302.350000 999.500000 303.650000 ;
      RECT 957.500000 302.350000 958.500000 303.650000 ;
      RECT 916.500000 302.350000 949.500000 303.650000 ;
      RECT 907.500000 302.350000 908.500000 303.650000 ;
      RECT 866.500000 302.350000 899.500000 303.650000 ;
      RECT 857.500000 302.350000 858.500000 303.650000 ;
      RECT 816.500000 302.350000 849.500000 303.650000 ;
      RECT 807.500000 302.350000 808.500000 303.650000 ;
      RECT 766.500000 302.350000 799.500000 303.650000 ;
      RECT 757.500000 302.350000 758.500000 303.650000 ;
      RECT 716.500000 302.350000 749.500000 303.650000 ;
      RECT 707.500000 302.350000 708.500000 303.650000 ;
      RECT 666.500000 302.350000 699.500000 303.650000 ;
      RECT 657.500000 302.350000 658.500000 303.650000 ;
      RECT 616.500000 302.350000 649.500000 303.650000 ;
      RECT 607.500000 302.350000 608.500000 303.650000 ;
      RECT 566.500000 302.350000 599.500000 303.650000 ;
      RECT 557.500000 302.350000 558.500000 303.650000 ;
      RECT 516.500000 302.350000 549.500000 303.650000 ;
      RECT 507.500000 302.350000 508.500000 303.650000 ;
      RECT 416.500000 302.350000 458.500000 303.730000 ;
      RECT 407.500000 302.350000 408.500000 303.650000 ;
      RECT 366.500000 302.350000 399.500000 303.650000 ;
      RECT 357.500000 302.350000 358.500000 303.650000 ;
      RECT 316.500000 302.350000 349.500000 303.650000 ;
      RECT 307.500000 302.350000 308.500000 303.650000 ;
      RECT 266.500000 302.350000 299.500000 303.650000 ;
      RECT 257.500000 302.350000 258.500000 303.650000 ;
      RECT 216.500000 302.350000 249.500000 303.650000 ;
      RECT 207.500000 302.350000 208.500000 303.650000 ;
      RECT 166.500000 302.350000 199.500000 303.650000 ;
      RECT 157.500000 302.350000 158.500000 303.650000 ;
      RECT 116.500000 302.350000 149.500000 303.650000 ;
      RECT 107.500000 302.350000 108.500000 303.650000 ;
      RECT 66.500000 302.350000 99.500000 303.650000 ;
      RECT 57.500000 302.350000 58.500000 303.650000 ;
      RECT 29.500000 302.350000 49.500000 303.650000 ;
      RECT 15.500000 302.350000 16.500000 303.650000 ;
      RECT 1157.500000 301.650000 1170.500000 302.350000 ;
      RECT 1107.500000 301.650000 1149.500000 302.350000 ;
      RECT 1057.500000 301.650000 1099.500000 302.350000 ;
      RECT 1007.500000 301.650000 1049.500000 302.350000 ;
      RECT 957.500000 301.650000 999.500000 302.350000 ;
      RECT 907.500000 301.650000 949.500000 302.350000 ;
      RECT 857.500000 301.650000 899.500000 302.350000 ;
      RECT 807.500000 301.650000 849.500000 302.350000 ;
      RECT 757.500000 301.650000 799.500000 302.350000 ;
      RECT 707.500000 301.650000 749.500000 302.350000 ;
      RECT 657.500000 301.650000 699.500000 302.350000 ;
      RECT 607.500000 301.650000 649.500000 302.350000 ;
      RECT 557.500000 301.650000 599.500000 302.350000 ;
      RECT 507.500000 301.650000 549.500000 302.350000 ;
      RECT 407.500000 301.650000 458.500000 302.350000 ;
      RECT 357.500000 301.650000 399.500000 302.350000 ;
      RECT 307.500000 301.650000 349.500000 302.350000 ;
      RECT 257.500000 301.650000 299.500000 302.350000 ;
      RECT 207.500000 301.650000 249.500000 302.350000 ;
      RECT 157.500000 301.650000 199.500000 302.350000 ;
      RECT 107.500000 301.650000 149.500000 302.350000 ;
      RECT 57.500000 301.650000 99.500000 302.350000 ;
      RECT 15.500000 301.650000 49.500000 302.350000 ;
      RECT 1183.500000 300.350000 1186.000000 303.650000 ;
      RECT 1169.500000 300.350000 1170.500000 301.650000 ;
      RECT 1116.500000 300.350000 1149.500000 301.650000 ;
      RECT 1107.500000 300.350000 1108.500000 301.650000 ;
      RECT 1066.500000 300.350000 1099.500000 301.650000 ;
      RECT 1057.500000 300.350000 1058.500000 301.650000 ;
      RECT 1016.500000 300.350000 1049.500000 301.650000 ;
      RECT 1007.500000 300.350000 1008.500000 301.650000 ;
      RECT 966.500000 300.350000 999.500000 301.650000 ;
      RECT 957.500000 300.350000 958.500000 301.650000 ;
      RECT 916.500000 300.350000 949.500000 301.650000 ;
      RECT 907.500000 300.350000 908.500000 301.650000 ;
      RECT 866.500000 300.350000 899.500000 301.650000 ;
      RECT 857.500000 300.350000 858.500000 301.650000 ;
      RECT 816.500000 300.350000 849.500000 301.650000 ;
      RECT 807.500000 300.350000 808.500000 301.650000 ;
      RECT 766.500000 300.350000 799.500000 301.650000 ;
      RECT 757.500000 300.350000 758.500000 301.650000 ;
      RECT 716.500000 300.350000 749.500000 301.650000 ;
      RECT 707.500000 300.350000 708.500000 301.650000 ;
      RECT 666.500000 300.350000 699.500000 301.650000 ;
      RECT 657.500000 300.350000 658.500000 301.650000 ;
      RECT 616.500000 300.350000 649.500000 301.650000 ;
      RECT 607.500000 300.350000 608.500000 301.650000 ;
      RECT 566.500000 300.350000 599.500000 301.650000 ;
      RECT 557.500000 300.350000 558.500000 301.650000 ;
      RECT 516.500000 300.350000 549.500000 301.650000 ;
      RECT 507.500000 300.350000 508.500000 301.650000 ;
      RECT 466.500000 300.350000 499.500000 303.650000 ;
      RECT 407.500000 300.350000 408.500000 301.650000 ;
      RECT 366.500000 300.350000 399.500000 301.650000 ;
      RECT 357.500000 300.350000 358.500000 301.650000 ;
      RECT 316.500000 300.350000 349.500000 301.650000 ;
      RECT 307.500000 300.350000 308.500000 301.650000 ;
      RECT 266.500000 300.350000 299.500000 301.650000 ;
      RECT 257.500000 300.350000 258.500000 301.650000 ;
      RECT 216.500000 300.350000 249.500000 301.650000 ;
      RECT 207.500000 300.350000 208.500000 301.650000 ;
      RECT 166.500000 300.350000 199.500000 301.650000 ;
      RECT 157.500000 300.350000 158.500000 301.650000 ;
      RECT 116.500000 300.350000 149.500000 301.650000 ;
      RECT 107.500000 300.350000 108.500000 301.650000 ;
      RECT 66.500000 300.350000 99.500000 301.650000 ;
      RECT 57.500000 300.350000 58.500000 301.650000 ;
      RECT 29.500000 300.350000 49.500000 301.650000 ;
      RECT 15.500000 300.350000 16.500000 301.650000 ;
      RECT 0.000000 300.350000 2.500000 303.650000 ;
      RECT 466.500000 299.730000 508.500000 300.350000 ;
      RECT 416.500000 299.730000 458.500000 301.650000 ;
      RECT 1169.500000 299.650000 1186.000000 300.350000 ;
      RECT 1116.500000 299.650000 1156.500000 300.350000 ;
      RECT 1066.500000 299.650000 1108.500000 300.350000 ;
      RECT 1016.500000 299.650000 1058.500000 300.350000 ;
      RECT 966.500000 299.650000 1008.500000 300.350000 ;
      RECT 916.500000 299.650000 958.500000 300.350000 ;
      RECT 866.500000 299.650000 908.500000 300.350000 ;
      RECT 816.500000 299.650000 858.500000 300.350000 ;
      RECT 766.500000 299.650000 808.500000 300.350000 ;
      RECT 716.500000 299.650000 758.500000 300.350000 ;
      RECT 666.500000 299.650000 708.500000 300.350000 ;
      RECT 616.500000 299.650000 658.500000 300.350000 ;
      RECT 566.500000 299.650000 608.500000 300.350000 ;
      RECT 516.500000 299.650000 558.500000 300.350000 ;
      RECT 416.500000 299.650000 508.500000 299.730000 ;
      RECT 366.500000 299.650000 408.500000 300.350000 ;
      RECT 316.500000 299.650000 358.500000 300.350000 ;
      RECT 266.500000 299.650000 308.500000 300.350000 ;
      RECT 216.500000 299.650000 258.500000 300.350000 ;
      RECT 166.500000 299.650000 208.500000 300.350000 ;
      RECT 116.500000 299.650000 158.500000 300.350000 ;
      RECT 66.500000 299.650000 108.500000 300.350000 ;
      RECT 29.500000 299.650000 58.500000 300.350000 ;
      RECT 0.000000 299.650000 16.500000 300.350000 ;
      RECT 1169.500000 298.350000 1170.500000 299.650000 ;
      RECT 1116.500000 298.350000 1149.500000 299.650000 ;
      RECT 1107.500000 298.350000 1108.500000 299.650000 ;
      RECT 1066.500000 298.350000 1099.500000 299.650000 ;
      RECT 1057.500000 298.350000 1058.500000 299.650000 ;
      RECT 1016.500000 298.350000 1049.500000 299.650000 ;
      RECT 1007.500000 298.350000 1008.500000 299.650000 ;
      RECT 966.500000 298.350000 999.500000 299.650000 ;
      RECT 957.500000 298.350000 958.500000 299.650000 ;
      RECT 916.500000 298.350000 949.500000 299.650000 ;
      RECT 907.500000 298.350000 908.500000 299.650000 ;
      RECT 866.500000 298.350000 899.500000 299.650000 ;
      RECT 857.500000 298.350000 858.500000 299.650000 ;
      RECT 816.500000 298.350000 849.500000 299.650000 ;
      RECT 807.500000 298.350000 808.500000 299.650000 ;
      RECT 766.500000 298.350000 799.500000 299.650000 ;
      RECT 757.500000 298.350000 758.500000 299.650000 ;
      RECT 716.500000 298.350000 749.500000 299.650000 ;
      RECT 707.500000 298.350000 708.500000 299.650000 ;
      RECT 666.500000 298.350000 699.500000 299.650000 ;
      RECT 657.500000 298.350000 658.500000 299.650000 ;
      RECT 616.500000 298.350000 649.500000 299.650000 ;
      RECT 607.500000 298.350000 608.500000 299.650000 ;
      RECT 566.500000 298.350000 599.500000 299.650000 ;
      RECT 557.500000 298.350000 558.500000 299.650000 ;
      RECT 516.500000 298.350000 549.500000 299.650000 ;
      RECT 507.500000 298.350000 508.500000 299.650000 ;
      RECT 416.500000 298.350000 449.500000 299.650000 ;
      RECT 407.500000 298.350000 408.500000 299.650000 ;
      RECT 366.500000 298.350000 399.500000 299.650000 ;
      RECT 357.500000 298.350000 358.500000 299.650000 ;
      RECT 316.500000 298.350000 349.500000 299.650000 ;
      RECT 307.500000 298.350000 308.500000 299.650000 ;
      RECT 266.500000 298.350000 299.500000 299.650000 ;
      RECT 257.500000 298.350000 258.500000 299.650000 ;
      RECT 216.500000 298.350000 249.500000 299.650000 ;
      RECT 207.500000 298.350000 208.500000 299.650000 ;
      RECT 166.500000 298.350000 199.500000 299.650000 ;
      RECT 157.500000 298.350000 158.500000 299.650000 ;
      RECT 116.500000 298.350000 149.500000 299.650000 ;
      RECT 107.500000 298.350000 108.500000 299.650000 ;
      RECT 66.500000 298.350000 99.500000 299.650000 ;
      RECT 57.500000 298.350000 58.500000 299.650000 ;
      RECT 29.500000 298.350000 49.500000 299.650000 ;
      RECT 15.500000 298.350000 16.500000 299.650000 ;
      RECT 1157.500000 297.650000 1170.500000 298.350000 ;
      RECT 1107.500000 297.650000 1149.500000 298.350000 ;
      RECT 1057.500000 297.650000 1099.500000 298.350000 ;
      RECT 1007.500000 297.650000 1049.500000 298.350000 ;
      RECT 957.500000 297.650000 999.500000 298.350000 ;
      RECT 907.500000 297.650000 949.500000 298.350000 ;
      RECT 857.500000 297.650000 899.500000 298.350000 ;
      RECT 807.500000 297.650000 849.500000 298.350000 ;
      RECT 757.500000 297.650000 799.500000 298.350000 ;
      RECT 707.500000 297.650000 749.500000 298.350000 ;
      RECT 657.500000 297.650000 699.500000 298.350000 ;
      RECT 607.500000 297.650000 649.500000 298.350000 ;
      RECT 557.500000 297.650000 599.500000 298.350000 ;
      RECT 507.500000 297.650000 549.500000 298.350000 ;
      RECT 457.500000 297.650000 499.500000 299.650000 ;
      RECT 407.500000 297.650000 449.500000 298.350000 ;
      RECT 357.500000 297.650000 399.500000 298.350000 ;
      RECT 307.500000 297.650000 349.500000 298.350000 ;
      RECT 257.500000 297.650000 299.500000 298.350000 ;
      RECT 207.500000 297.650000 249.500000 298.350000 ;
      RECT 157.500000 297.650000 199.500000 298.350000 ;
      RECT 107.500000 297.650000 149.500000 298.350000 ;
      RECT 57.500000 297.650000 99.500000 298.350000 ;
      RECT 15.500000 297.650000 49.500000 298.350000 ;
      RECT 1183.500000 296.350000 1186.000000 299.650000 ;
      RECT 1169.500000 296.350000 1170.500000 297.650000 ;
      RECT 1116.500000 296.350000 1149.500000 297.650000 ;
      RECT 1107.500000 296.350000 1108.500000 297.650000 ;
      RECT 1066.500000 296.350000 1099.500000 297.650000 ;
      RECT 1057.500000 296.350000 1058.500000 297.650000 ;
      RECT 1016.500000 296.350000 1049.500000 297.650000 ;
      RECT 1007.500000 296.350000 1008.500000 297.650000 ;
      RECT 966.500000 296.350000 999.500000 297.650000 ;
      RECT 957.500000 296.350000 958.500000 297.650000 ;
      RECT 916.500000 296.350000 949.500000 297.650000 ;
      RECT 907.500000 296.350000 908.500000 297.650000 ;
      RECT 866.500000 296.350000 899.500000 297.650000 ;
      RECT 857.500000 296.350000 858.500000 297.650000 ;
      RECT 816.500000 296.350000 849.500000 297.650000 ;
      RECT 807.500000 296.350000 808.500000 297.650000 ;
      RECT 766.500000 296.350000 799.500000 297.650000 ;
      RECT 757.500000 296.350000 758.500000 297.650000 ;
      RECT 716.500000 296.350000 749.500000 297.650000 ;
      RECT 707.500000 296.350000 708.500000 297.650000 ;
      RECT 666.500000 296.350000 699.500000 297.650000 ;
      RECT 657.500000 296.350000 658.500000 297.650000 ;
      RECT 616.500000 296.350000 649.500000 297.650000 ;
      RECT 607.500000 296.350000 608.500000 297.650000 ;
      RECT 566.500000 296.350000 599.500000 297.650000 ;
      RECT 557.500000 296.350000 558.500000 297.650000 ;
      RECT 516.500000 296.350000 549.500000 297.650000 ;
      RECT 507.500000 296.350000 508.500000 297.650000 ;
      RECT 466.500000 296.350000 499.500000 297.650000 ;
      RECT 457.500000 296.350000 458.500000 297.650000 ;
      RECT 416.500000 296.350000 449.500000 297.650000 ;
      RECT 407.500000 296.350000 408.500000 297.650000 ;
      RECT 366.500000 296.350000 399.500000 297.650000 ;
      RECT 357.500000 296.350000 358.500000 297.650000 ;
      RECT 316.500000 296.350000 349.500000 297.650000 ;
      RECT 307.500000 296.350000 308.500000 297.650000 ;
      RECT 266.500000 296.350000 299.500000 297.650000 ;
      RECT 257.500000 296.350000 258.500000 297.650000 ;
      RECT 216.500000 296.350000 249.500000 297.650000 ;
      RECT 207.500000 296.350000 208.500000 297.650000 ;
      RECT 166.500000 296.350000 199.500000 297.650000 ;
      RECT 157.500000 296.350000 158.500000 297.650000 ;
      RECT 116.500000 296.350000 149.500000 297.650000 ;
      RECT 107.500000 296.350000 108.500000 297.650000 ;
      RECT 66.500000 296.350000 99.500000 297.650000 ;
      RECT 57.500000 296.350000 58.500000 297.650000 ;
      RECT 29.500000 296.350000 49.500000 297.650000 ;
      RECT 15.500000 296.350000 16.500000 297.650000 ;
      RECT 0.000000 296.350000 2.500000 299.650000 ;
      RECT 1169.500000 295.650000 1186.000000 296.350000 ;
      RECT 1116.500000 295.650000 1156.500000 296.350000 ;
      RECT 1066.500000 295.650000 1108.500000 296.350000 ;
      RECT 1016.500000 295.650000 1058.500000 296.350000 ;
      RECT 966.500000 295.650000 1008.500000 296.350000 ;
      RECT 916.500000 295.650000 958.500000 296.350000 ;
      RECT 866.500000 295.650000 908.500000 296.350000 ;
      RECT 816.500000 295.650000 858.500000 296.350000 ;
      RECT 766.500000 295.650000 808.500000 296.350000 ;
      RECT 716.500000 295.650000 758.500000 296.350000 ;
      RECT 666.500000 295.650000 708.500000 296.350000 ;
      RECT 616.500000 295.650000 658.500000 296.350000 ;
      RECT 566.500000 295.650000 608.500000 296.350000 ;
      RECT 516.500000 295.650000 558.500000 296.350000 ;
      RECT 466.500000 295.650000 508.500000 296.350000 ;
      RECT 416.500000 295.650000 458.500000 296.350000 ;
      RECT 366.500000 295.650000 408.500000 296.350000 ;
      RECT 316.500000 295.650000 358.500000 296.350000 ;
      RECT 266.500000 295.650000 308.500000 296.350000 ;
      RECT 216.500000 295.650000 258.500000 296.350000 ;
      RECT 166.500000 295.650000 208.500000 296.350000 ;
      RECT 116.500000 295.650000 158.500000 296.350000 ;
      RECT 66.500000 295.650000 108.500000 296.350000 ;
      RECT 29.500000 295.650000 58.500000 296.350000 ;
      RECT 0.000000 295.650000 16.500000 296.350000 ;
      RECT 1169.500000 294.350000 1170.500000 295.650000 ;
      RECT 1116.500000 294.350000 1149.500000 295.650000 ;
      RECT 1107.500000 294.350000 1108.500000 295.650000 ;
      RECT 1066.500000 294.350000 1099.500000 295.650000 ;
      RECT 1057.500000 294.350000 1058.500000 295.650000 ;
      RECT 1016.500000 294.350000 1049.500000 295.650000 ;
      RECT 1007.500000 294.350000 1008.500000 295.650000 ;
      RECT 966.500000 294.350000 999.500000 295.650000 ;
      RECT 957.500000 294.350000 958.500000 295.650000 ;
      RECT 916.500000 294.350000 949.500000 295.650000 ;
      RECT 907.500000 294.350000 908.500000 295.650000 ;
      RECT 866.500000 294.350000 899.500000 295.650000 ;
      RECT 857.500000 294.350000 858.500000 295.650000 ;
      RECT 816.500000 294.350000 849.500000 295.650000 ;
      RECT 807.500000 294.350000 808.500000 295.650000 ;
      RECT 766.500000 294.350000 799.500000 295.650000 ;
      RECT 757.500000 294.350000 758.500000 295.650000 ;
      RECT 716.500000 294.350000 749.500000 295.650000 ;
      RECT 707.500000 294.350000 708.500000 295.650000 ;
      RECT 666.500000 294.350000 699.500000 295.650000 ;
      RECT 657.500000 294.350000 658.500000 295.650000 ;
      RECT 616.500000 294.350000 649.500000 295.650000 ;
      RECT 607.500000 294.350000 608.500000 295.650000 ;
      RECT 566.500000 294.350000 599.500000 295.650000 ;
      RECT 557.500000 294.350000 558.500000 295.650000 ;
      RECT 516.500000 294.350000 549.500000 295.650000 ;
      RECT 507.500000 294.350000 508.500000 295.650000 ;
      RECT 466.500000 294.350000 499.500000 295.650000 ;
      RECT 457.500000 294.350000 458.500000 295.650000 ;
      RECT 416.500000 294.350000 449.500000 295.650000 ;
      RECT 407.500000 294.350000 408.500000 295.650000 ;
      RECT 366.500000 294.350000 399.500000 295.650000 ;
      RECT 357.500000 294.350000 358.500000 295.650000 ;
      RECT 316.500000 294.350000 349.500000 295.650000 ;
      RECT 307.500000 294.350000 308.500000 295.650000 ;
      RECT 266.500000 294.350000 299.500000 295.650000 ;
      RECT 257.500000 294.350000 258.500000 295.650000 ;
      RECT 216.500000 294.350000 249.500000 295.650000 ;
      RECT 207.500000 294.350000 208.500000 295.650000 ;
      RECT 166.500000 294.350000 199.500000 295.650000 ;
      RECT 157.500000 294.350000 158.500000 295.650000 ;
      RECT 116.500000 294.350000 149.500000 295.650000 ;
      RECT 107.500000 294.350000 108.500000 295.650000 ;
      RECT 66.500000 294.350000 99.500000 295.650000 ;
      RECT 57.500000 294.350000 58.500000 295.650000 ;
      RECT 29.500000 294.350000 49.500000 295.650000 ;
      RECT 15.500000 294.350000 16.500000 295.650000 ;
      RECT 1157.500000 293.650000 1170.500000 294.350000 ;
      RECT 1107.500000 293.650000 1149.500000 294.350000 ;
      RECT 1057.500000 293.650000 1099.500000 294.350000 ;
      RECT 1007.500000 293.650000 1049.500000 294.350000 ;
      RECT 957.500000 293.650000 999.500000 294.350000 ;
      RECT 907.500000 293.650000 949.500000 294.350000 ;
      RECT 857.500000 293.650000 899.500000 294.350000 ;
      RECT 807.500000 293.650000 849.500000 294.350000 ;
      RECT 757.500000 293.650000 799.500000 294.350000 ;
      RECT 707.500000 293.650000 749.500000 294.350000 ;
      RECT 657.500000 293.650000 699.500000 294.350000 ;
      RECT 607.500000 293.650000 649.500000 294.350000 ;
      RECT 557.500000 293.650000 599.500000 294.350000 ;
      RECT 507.500000 293.650000 549.500000 294.350000 ;
      RECT 457.500000 293.650000 499.500000 294.350000 ;
      RECT 407.500000 293.650000 449.500000 294.350000 ;
      RECT 357.500000 293.650000 399.500000 294.350000 ;
      RECT 307.500000 293.650000 349.500000 294.350000 ;
      RECT 257.500000 293.650000 299.500000 294.350000 ;
      RECT 207.500000 293.650000 249.500000 294.350000 ;
      RECT 157.500000 293.650000 199.500000 294.350000 ;
      RECT 107.500000 293.650000 149.500000 294.350000 ;
      RECT 57.500000 293.650000 99.500000 294.350000 ;
      RECT 15.500000 293.650000 49.500000 294.350000 ;
      RECT 1183.500000 292.350000 1186.000000 295.650000 ;
      RECT 1169.500000 292.350000 1170.500000 293.650000 ;
      RECT 1116.500000 292.350000 1149.500000 293.650000 ;
      RECT 1107.500000 292.350000 1108.500000 293.650000 ;
      RECT 1066.500000 292.350000 1099.500000 293.650000 ;
      RECT 1057.500000 292.350000 1058.500000 293.650000 ;
      RECT 1016.500000 292.350000 1049.500000 293.650000 ;
      RECT 1007.500000 292.350000 1008.500000 293.650000 ;
      RECT 966.500000 292.350000 999.500000 293.650000 ;
      RECT 957.500000 292.350000 958.500000 293.650000 ;
      RECT 916.500000 292.350000 949.500000 293.650000 ;
      RECT 907.500000 292.350000 908.500000 293.650000 ;
      RECT 866.500000 292.350000 899.500000 293.650000 ;
      RECT 857.500000 292.350000 858.500000 293.650000 ;
      RECT 816.500000 292.350000 849.500000 293.650000 ;
      RECT 807.500000 292.350000 808.500000 293.650000 ;
      RECT 766.500000 292.350000 799.500000 293.650000 ;
      RECT 757.500000 292.350000 758.500000 293.650000 ;
      RECT 716.500000 292.350000 749.500000 293.650000 ;
      RECT 707.500000 292.350000 708.500000 293.650000 ;
      RECT 666.500000 292.350000 699.500000 293.650000 ;
      RECT 657.500000 292.350000 658.500000 293.650000 ;
      RECT 616.500000 292.350000 649.500000 293.650000 ;
      RECT 607.500000 292.350000 608.500000 293.650000 ;
      RECT 566.500000 292.350000 599.500000 293.650000 ;
      RECT 557.500000 292.350000 558.500000 293.650000 ;
      RECT 516.500000 292.350000 549.500000 293.650000 ;
      RECT 507.500000 292.350000 508.500000 293.650000 ;
      RECT 466.500000 292.350000 499.500000 293.650000 ;
      RECT 457.500000 292.350000 458.500000 293.650000 ;
      RECT 416.500000 292.350000 449.500000 293.650000 ;
      RECT 407.500000 292.350000 408.500000 293.650000 ;
      RECT 366.500000 292.350000 399.500000 293.650000 ;
      RECT 357.500000 292.350000 358.500000 293.650000 ;
      RECT 316.500000 292.350000 349.500000 293.650000 ;
      RECT 307.500000 292.350000 308.500000 293.650000 ;
      RECT 266.500000 292.350000 299.500000 293.650000 ;
      RECT 257.500000 292.350000 258.500000 293.650000 ;
      RECT 216.500000 292.350000 249.500000 293.650000 ;
      RECT 207.500000 292.350000 208.500000 293.650000 ;
      RECT 166.500000 292.350000 199.500000 293.650000 ;
      RECT 157.500000 292.350000 158.500000 293.650000 ;
      RECT 116.500000 292.350000 149.500000 293.650000 ;
      RECT 107.500000 292.350000 108.500000 293.650000 ;
      RECT 66.500000 292.350000 99.500000 293.650000 ;
      RECT 57.500000 292.350000 58.500000 293.650000 ;
      RECT 29.500000 292.350000 49.500000 293.650000 ;
      RECT 15.500000 292.350000 16.500000 293.650000 ;
      RECT 0.000000 292.350000 2.500000 295.650000 ;
      RECT 1169.500000 291.650000 1186.000000 292.350000 ;
      RECT 1116.500000 291.650000 1156.500000 292.350000 ;
      RECT 1066.500000 291.650000 1108.500000 292.350000 ;
      RECT 1016.500000 291.650000 1058.500000 292.350000 ;
      RECT 966.500000 291.650000 1008.500000 292.350000 ;
      RECT 916.500000 291.650000 958.500000 292.350000 ;
      RECT 866.500000 291.650000 908.500000 292.350000 ;
      RECT 816.500000 291.650000 858.500000 292.350000 ;
      RECT 766.500000 291.650000 808.500000 292.350000 ;
      RECT 716.500000 291.650000 758.500000 292.350000 ;
      RECT 666.500000 291.650000 708.500000 292.350000 ;
      RECT 616.500000 291.650000 658.500000 292.350000 ;
      RECT 566.500000 291.650000 608.500000 292.350000 ;
      RECT 516.500000 291.650000 558.500000 292.350000 ;
      RECT 466.500000 291.650000 508.500000 292.350000 ;
      RECT 416.500000 291.650000 458.500000 292.350000 ;
      RECT 366.500000 291.650000 408.500000 292.350000 ;
      RECT 316.500000 291.650000 358.500000 292.350000 ;
      RECT 266.500000 291.650000 308.500000 292.350000 ;
      RECT 216.500000 291.650000 258.500000 292.350000 ;
      RECT 166.500000 291.650000 208.500000 292.350000 ;
      RECT 116.500000 291.650000 158.500000 292.350000 ;
      RECT 66.500000 291.650000 108.500000 292.350000 ;
      RECT 29.500000 291.650000 58.500000 292.350000 ;
      RECT 0.000000 291.650000 16.500000 292.350000 ;
      RECT 1169.500000 290.350000 1170.500000 291.650000 ;
      RECT 1116.500000 290.350000 1149.500000 291.650000 ;
      RECT 1107.500000 290.350000 1108.500000 291.650000 ;
      RECT 1066.500000 290.350000 1099.500000 291.650000 ;
      RECT 1057.500000 290.350000 1058.500000 291.650000 ;
      RECT 1016.500000 290.350000 1049.500000 291.650000 ;
      RECT 1007.500000 290.350000 1008.500000 291.650000 ;
      RECT 966.500000 290.350000 999.500000 291.650000 ;
      RECT 957.500000 290.350000 958.500000 291.650000 ;
      RECT 916.500000 290.350000 949.500000 291.650000 ;
      RECT 907.500000 290.350000 908.500000 291.650000 ;
      RECT 866.500000 290.350000 899.500000 291.650000 ;
      RECT 857.500000 290.350000 858.500000 291.650000 ;
      RECT 816.500000 290.350000 849.500000 291.650000 ;
      RECT 807.500000 290.350000 808.500000 291.650000 ;
      RECT 766.500000 290.350000 799.500000 291.650000 ;
      RECT 757.500000 290.350000 758.500000 291.650000 ;
      RECT 716.500000 290.350000 749.500000 291.650000 ;
      RECT 707.500000 290.350000 708.500000 291.650000 ;
      RECT 666.500000 290.350000 699.500000 291.650000 ;
      RECT 657.500000 290.350000 658.500000 291.650000 ;
      RECT 616.500000 290.350000 649.500000 291.650000 ;
      RECT 607.500000 290.350000 608.500000 291.650000 ;
      RECT 566.500000 290.350000 599.500000 291.650000 ;
      RECT 557.500000 290.350000 558.500000 291.650000 ;
      RECT 516.500000 290.350000 549.500000 291.650000 ;
      RECT 507.500000 290.350000 508.500000 291.650000 ;
      RECT 466.500000 290.350000 499.500000 291.650000 ;
      RECT 457.500000 290.350000 458.500000 291.650000 ;
      RECT 416.500000 290.350000 449.500000 291.650000 ;
      RECT 407.500000 290.350000 408.500000 291.650000 ;
      RECT 366.500000 290.350000 399.500000 291.650000 ;
      RECT 357.500000 290.350000 358.500000 291.650000 ;
      RECT 316.500000 290.350000 349.500000 291.650000 ;
      RECT 307.500000 290.350000 308.500000 291.650000 ;
      RECT 266.500000 290.350000 299.500000 291.650000 ;
      RECT 257.500000 290.350000 258.500000 291.650000 ;
      RECT 216.500000 290.350000 249.500000 291.650000 ;
      RECT 207.500000 290.350000 208.500000 291.650000 ;
      RECT 166.500000 290.350000 199.500000 291.650000 ;
      RECT 157.500000 290.350000 158.500000 291.650000 ;
      RECT 116.500000 290.350000 149.500000 291.650000 ;
      RECT 107.500000 290.350000 108.500000 291.650000 ;
      RECT 66.500000 290.350000 99.500000 291.650000 ;
      RECT 57.500000 290.350000 58.500000 291.650000 ;
      RECT 29.500000 290.350000 49.500000 291.650000 ;
      RECT 15.500000 290.350000 16.500000 291.650000 ;
      RECT 1157.500000 289.650000 1170.500000 290.350000 ;
      RECT 1107.500000 289.650000 1149.500000 290.350000 ;
      RECT 1057.500000 289.650000 1099.500000 290.350000 ;
      RECT 1007.500000 289.650000 1049.500000 290.350000 ;
      RECT 957.500000 289.650000 999.500000 290.350000 ;
      RECT 907.500000 289.650000 949.500000 290.350000 ;
      RECT 857.500000 289.650000 899.500000 290.350000 ;
      RECT 807.500000 289.650000 849.500000 290.350000 ;
      RECT 757.500000 289.650000 799.500000 290.350000 ;
      RECT 707.500000 289.650000 749.500000 290.350000 ;
      RECT 657.500000 289.650000 699.500000 290.350000 ;
      RECT 607.500000 289.650000 649.500000 290.350000 ;
      RECT 557.500000 289.650000 599.500000 290.350000 ;
      RECT 507.500000 289.650000 549.500000 290.350000 ;
      RECT 457.500000 289.650000 499.500000 290.350000 ;
      RECT 407.500000 289.650000 449.500000 290.350000 ;
      RECT 357.500000 289.650000 399.500000 290.350000 ;
      RECT 307.500000 289.650000 349.500000 290.350000 ;
      RECT 257.500000 289.650000 299.500000 290.350000 ;
      RECT 207.500000 289.650000 249.500000 290.350000 ;
      RECT 157.500000 289.650000 199.500000 290.350000 ;
      RECT 107.500000 289.650000 149.500000 290.350000 ;
      RECT 57.500000 289.650000 99.500000 290.350000 ;
      RECT 15.500000 289.650000 49.500000 290.350000 ;
      RECT 1183.500000 288.350000 1186.000000 291.650000 ;
      RECT 1169.500000 288.350000 1170.500000 289.650000 ;
      RECT 1116.500000 288.350000 1149.500000 289.650000 ;
      RECT 1107.500000 288.350000 1108.500000 289.650000 ;
      RECT 1066.500000 288.350000 1099.500000 289.650000 ;
      RECT 1057.500000 288.350000 1058.500000 289.650000 ;
      RECT 1016.500000 288.350000 1049.500000 289.650000 ;
      RECT 1007.500000 288.350000 1008.500000 289.650000 ;
      RECT 966.500000 288.350000 999.500000 289.650000 ;
      RECT 957.500000 288.350000 958.500000 289.650000 ;
      RECT 916.500000 288.350000 949.500000 289.650000 ;
      RECT 907.500000 288.350000 908.500000 289.650000 ;
      RECT 866.500000 288.350000 899.500000 289.650000 ;
      RECT 857.500000 288.350000 858.500000 289.650000 ;
      RECT 816.500000 288.350000 849.500000 289.650000 ;
      RECT 807.500000 288.350000 808.500000 289.650000 ;
      RECT 766.500000 288.350000 799.500000 289.650000 ;
      RECT 757.500000 288.350000 758.500000 289.650000 ;
      RECT 716.500000 288.350000 749.500000 289.650000 ;
      RECT 707.500000 288.350000 708.500000 289.650000 ;
      RECT 666.500000 288.350000 699.500000 289.650000 ;
      RECT 657.500000 288.350000 658.500000 289.650000 ;
      RECT 616.500000 288.350000 649.500000 289.650000 ;
      RECT 607.500000 288.350000 608.500000 289.650000 ;
      RECT 566.500000 288.350000 599.500000 289.650000 ;
      RECT 557.500000 288.350000 558.500000 289.650000 ;
      RECT 516.500000 288.350000 549.500000 289.650000 ;
      RECT 507.500000 288.350000 508.500000 289.650000 ;
      RECT 466.500000 288.350000 499.500000 289.650000 ;
      RECT 457.500000 288.350000 458.500000 289.650000 ;
      RECT 416.500000 288.350000 449.500000 289.650000 ;
      RECT 407.500000 288.350000 408.500000 289.650000 ;
      RECT 366.500000 288.350000 399.500000 289.650000 ;
      RECT 357.500000 288.350000 358.500000 289.650000 ;
      RECT 316.500000 288.350000 349.500000 289.650000 ;
      RECT 307.500000 288.350000 308.500000 289.650000 ;
      RECT 266.500000 288.350000 299.500000 289.650000 ;
      RECT 257.500000 288.350000 258.500000 289.650000 ;
      RECT 216.500000 288.350000 249.500000 289.650000 ;
      RECT 207.500000 288.350000 208.500000 289.650000 ;
      RECT 166.500000 288.350000 199.500000 289.650000 ;
      RECT 157.500000 288.350000 158.500000 289.650000 ;
      RECT 116.500000 288.350000 149.500000 289.650000 ;
      RECT 107.500000 288.350000 108.500000 289.650000 ;
      RECT 66.500000 288.350000 99.500000 289.650000 ;
      RECT 57.500000 288.350000 58.500000 289.650000 ;
      RECT 29.500000 288.350000 49.500000 289.650000 ;
      RECT 15.500000 288.350000 16.500000 289.650000 ;
      RECT 0.000000 288.350000 2.500000 291.650000 ;
      RECT 1169.500000 287.650000 1186.000000 288.350000 ;
      RECT 1116.500000 287.650000 1156.500000 288.350000 ;
      RECT 1066.500000 287.650000 1108.500000 288.350000 ;
      RECT 1016.500000 287.650000 1058.500000 288.350000 ;
      RECT 966.500000 287.650000 1008.500000 288.350000 ;
      RECT 916.500000 287.650000 958.500000 288.350000 ;
      RECT 866.500000 287.650000 908.500000 288.350000 ;
      RECT 816.500000 287.650000 858.500000 288.350000 ;
      RECT 766.500000 287.650000 808.500000 288.350000 ;
      RECT 716.500000 287.650000 758.500000 288.350000 ;
      RECT 666.500000 287.650000 708.500000 288.350000 ;
      RECT 616.500000 287.650000 658.500000 288.350000 ;
      RECT 566.500000 287.650000 608.500000 288.350000 ;
      RECT 516.500000 287.650000 558.500000 288.350000 ;
      RECT 466.500000 287.650000 508.500000 288.350000 ;
      RECT 416.500000 287.650000 458.500000 288.350000 ;
      RECT 366.500000 287.650000 408.500000 288.350000 ;
      RECT 316.500000 287.650000 358.500000 288.350000 ;
      RECT 266.500000 287.650000 308.500000 288.350000 ;
      RECT 216.500000 287.650000 258.500000 288.350000 ;
      RECT 166.500000 287.650000 208.500000 288.350000 ;
      RECT 116.500000 287.650000 158.500000 288.350000 ;
      RECT 66.500000 287.650000 108.500000 288.350000 ;
      RECT 29.500000 287.650000 58.500000 288.350000 ;
      RECT 0.000000 287.650000 16.500000 288.350000 ;
      RECT 1169.500000 286.350000 1170.500000 287.650000 ;
      RECT 1116.500000 286.350000 1149.500000 287.650000 ;
      RECT 1107.500000 286.350000 1108.500000 287.650000 ;
      RECT 1066.500000 286.350000 1099.500000 287.650000 ;
      RECT 1057.500000 286.350000 1058.500000 287.650000 ;
      RECT 1016.500000 286.350000 1049.500000 287.650000 ;
      RECT 1007.500000 286.350000 1008.500000 287.650000 ;
      RECT 966.500000 286.350000 999.500000 287.650000 ;
      RECT 957.500000 286.350000 958.500000 287.650000 ;
      RECT 916.500000 286.350000 949.500000 287.650000 ;
      RECT 907.500000 286.350000 908.500000 287.650000 ;
      RECT 866.500000 286.350000 899.500000 287.650000 ;
      RECT 857.500000 286.350000 858.500000 287.650000 ;
      RECT 816.500000 286.350000 849.500000 287.650000 ;
      RECT 807.500000 286.350000 808.500000 287.650000 ;
      RECT 766.500000 286.350000 799.500000 287.650000 ;
      RECT 757.500000 286.350000 758.500000 287.650000 ;
      RECT 716.500000 286.350000 749.500000 287.650000 ;
      RECT 707.500000 286.350000 708.500000 287.650000 ;
      RECT 666.500000 286.350000 699.500000 287.650000 ;
      RECT 657.500000 286.350000 658.500000 287.650000 ;
      RECT 616.500000 286.350000 649.500000 287.650000 ;
      RECT 607.500000 286.350000 608.500000 287.650000 ;
      RECT 566.500000 286.350000 599.500000 287.650000 ;
      RECT 557.500000 286.350000 558.500000 287.650000 ;
      RECT 516.500000 286.350000 549.500000 287.650000 ;
      RECT 507.500000 286.350000 508.500000 287.650000 ;
      RECT 466.500000 286.350000 499.500000 287.650000 ;
      RECT 457.500000 286.350000 458.500000 287.650000 ;
      RECT 416.500000 286.350000 449.500000 287.650000 ;
      RECT 407.500000 286.350000 408.500000 287.650000 ;
      RECT 366.500000 286.350000 399.500000 287.650000 ;
      RECT 357.500000 286.350000 358.500000 287.650000 ;
      RECT 316.500000 286.350000 349.500000 287.650000 ;
      RECT 307.500000 286.350000 308.500000 287.650000 ;
      RECT 266.500000 286.350000 299.500000 287.650000 ;
      RECT 257.500000 286.350000 258.500000 287.650000 ;
      RECT 216.500000 286.350000 249.500000 287.650000 ;
      RECT 207.500000 286.350000 208.500000 287.650000 ;
      RECT 166.500000 286.350000 199.500000 287.650000 ;
      RECT 157.500000 286.350000 158.500000 287.650000 ;
      RECT 116.500000 286.350000 149.500000 287.650000 ;
      RECT 107.500000 286.350000 108.500000 287.650000 ;
      RECT 66.500000 286.350000 99.500000 287.650000 ;
      RECT 57.500000 286.350000 58.500000 287.650000 ;
      RECT 29.500000 286.350000 49.500000 287.650000 ;
      RECT 15.500000 286.350000 16.500000 287.650000 ;
      RECT 1157.500000 285.650000 1170.500000 286.350000 ;
      RECT 1107.500000 285.650000 1149.500000 286.350000 ;
      RECT 1057.500000 285.650000 1099.500000 286.350000 ;
      RECT 1007.500000 285.650000 1049.500000 286.350000 ;
      RECT 957.500000 285.650000 999.500000 286.350000 ;
      RECT 907.500000 285.650000 949.500000 286.350000 ;
      RECT 857.500000 285.650000 899.500000 286.350000 ;
      RECT 807.500000 285.650000 849.500000 286.350000 ;
      RECT 757.500000 285.650000 799.500000 286.350000 ;
      RECT 707.500000 285.650000 749.500000 286.350000 ;
      RECT 657.500000 285.650000 699.500000 286.350000 ;
      RECT 607.500000 285.650000 649.500000 286.350000 ;
      RECT 557.500000 285.650000 599.500000 286.350000 ;
      RECT 507.500000 285.650000 549.500000 286.350000 ;
      RECT 457.500000 285.650000 499.500000 286.350000 ;
      RECT 407.500000 285.650000 449.500000 286.350000 ;
      RECT 357.500000 285.650000 399.500000 286.350000 ;
      RECT 307.500000 285.650000 349.500000 286.350000 ;
      RECT 257.500000 285.650000 299.500000 286.350000 ;
      RECT 207.500000 285.650000 249.500000 286.350000 ;
      RECT 157.500000 285.650000 199.500000 286.350000 ;
      RECT 107.500000 285.650000 149.500000 286.350000 ;
      RECT 57.500000 285.650000 99.500000 286.350000 ;
      RECT 15.500000 285.650000 49.500000 286.350000 ;
      RECT 1183.500000 284.350000 1186.000000 287.650000 ;
      RECT 1169.500000 284.350000 1170.500000 285.650000 ;
      RECT 1116.500000 284.350000 1149.500000 285.650000 ;
      RECT 1107.500000 284.350000 1108.500000 285.650000 ;
      RECT 1066.500000 284.350000 1099.500000 285.650000 ;
      RECT 1057.500000 284.350000 1058.500000 285.650000 ;
      RECT 1016.500000 284.350000 1049.500000 285.650000 ;
      RECT 1007.500000 284.350000 1008.500000 285.650000 ;
      RECT 966.500000 284.350000 999.500000 285.650000 ;
      RECT 957.500000 284.350000 958.500000 285.650000 ;
      RECT 916.500000 284.350000 949.500000 285.650000 ;
      RECT 907.500000 284.350000 908.500000 285.650000 ;
      RECT 866.500000 284.350000 899.500000 285.650000 ;
      RECT 857.500000 284.350000 858.500000 285.650000 ;
      RECT 816.500000 284.350000 849.500000 285.650000 ;
      RECT 807.500000 284.350000 808.500000 285.650000 ;
      RECT 766.500000 284.350000 799.500000 285.650000 ;
      RECT 757.500000 284.350000 758.500000 285.650000 ;
      RECT 716.500000 284.350000 749.500000 285.650000 ;
      RECT 707.500000 284.350000 708.500000 285.650000 ;
      RECT 666.500000 284.350000 699.500000 285.650000 ;
      RECT 657.500000 284.350000 658.500000 285.650000 ;
      RECT 616.500000 284.350000 649.500000 285.650000 ;
      RECT 607.500000 284.350000 608.500000 285.650000 ;
      RECT 566.500000 284.350000 599.500000 285.650000 ;
      RECT 557.500000 284.350000 558.500000 285.650000 ;
      RECT 516.500000 284.350000 549.500000 285.650000 ;
      RECT 507.500000 284.350000 508.500000 285.650000 ;
      RECT 466.500000 284.350000 499.500000 285.650000 ;
      RECT 457.500000 284.350000 458.500000 285.650000 ;
      RECT 416.500000 284.350000 449.500000 285.650000 ;
      RECT 407.500000 284.350000 408.500000 285.650000 ;
      RECT 366.500000 284.350000 399.500000 285.650000 ;
      RECT 357.500000 284.350000 358.500000 285.650000 ;
      RECT 316.500000 284.350000 349.500000 285.650000 ;
      RECT 307.500000 284.350000 308.500000 285.650000 ;
      RECT 266.500000 284.350000 299.500000 285.650000 ;
      RECT 257.500000 284.350000 258.500000 285.650000 ;
      RECT 216.500000 284.350000 249.500000 285.650000 ;
      RECT 207.500000 284.350000 208.500000 285.650000 ;
      RECT 166.500000 284.350000 199.500000 285.650000 ;
      RECT 157.500000 284.350000 158.500000 285.650000 ;
      RECT 116.500000 284.350000 149.500000 285.650000 ;
      RECT 107.500000 284.350000 108.500000 285.650000 ;
      RECT 66.500000 284.350000 99.500000 285.650000 ;
      RECT 57.500000 284.350000 58.500000 285.650000 ;
      RECT 29.500000 284.350000 49.500000 285.650000 ;
      RECT 15.500000 284.350000 16.500000 285.650000 ;
      RECT 0.000000 284.350000 2.500000 287.650000 ;
      RECT 1169.500000 283.650000 1186.000000 284.350000 ;
      RECT 1116.500000 283.650000 1156.500000 284.350000 ;
      RECT 1066.500000 283.650000 1108.500000 284.350000 ;
      RECT 1016.500000 283.650000 1058.500000 284.350000 ;
      RECT 966.500000 283.650000 1008.500000 284.350000 ;
      RECT 916.500000 283.650000 958.500000 284.350000 ;
      RECT 866.500000 283.650000 908.500000 284.350000 ;
      RECT 816.500000 283.650000 858.500000 284.350000 ;
      RECT 766.500000 283.650000 808.500000 284.350000 ;
      RECT 716.500000 283.650000 758.500000 284.350000 ;
      RECT 666.500000 283.650000 708.500000 284.350000 ;
      RECT 616.500000 283.650000 658.500000 284.350000 ;
      RECT 566.500000 283.650000 608.500000 284.350000 ;
      RECT 516.500000 283.650000 558.500000 284.350000 ;
      RECT 466.500000 283.650000 508.500000 284.350000 ;
      RECT 416.500000 283.650000 458.500000 284.350000 ;
      RECT 366.500000 283.650000 408.500000 284.350000 ;
      RECT 316.500000 283.650000 358.500000 284.350000 ;
      RECT 266.500000 283.650000 308.500000 284.350000 ;
      RECT 216.500000 283.650000 258.500000 284.350000 ;
      RECT 166.500000 283.650000 208.500000 284.350000 ;
      RECT 116.500000 283.650000 158.500000 284.350000 ;
      RECT 66.500000 283.650000 108.500000 284.350000 ;
      RECT 29.500000 283.650000 58.500000 284.350000 ;
      RECT 0.000000 283.650000 16.500000 284.350000 ;
      RECT 1169.500000 282.350000 1170.500000 283.650000 ;
      RECT 1116.500000 282.350000 1149.500000 283.650000 ;
      RECT 1107.500000 282.350000 1108.500000 283.650000 ;
      RECT 1066.500000 282.350000 1099.500000 283.650000 ;
      RECT 1057.500000 282.350000 1058.500000 283.650000 ;
      RECT 1016.500000 282.350000 1049.500000 283.650000 ;
      RECT 1007.500000 282.350000 1008.500000 283.650000 ;
      RECT 966.500000 282.350000 999.500000 283.650000 ;
      RECT 957.500000 282.350000 958.500000 283.650000 ;
      RECT 916.500000 282.350000 949.500000 283.650000 ;
      RECT 907.500000 282.350000 908.500000 283.650000 ;
      RECT 866.500000 282.350000 899.500000 283.650000 ;
      RECT 857.500000 282.350000 858.500000 283.650000 ;
      RECT 816.500000 282.350000 849.500000 283.650000 ;
      RECT 807.500000 282.350000 808.500000 283.650000 ;
      RECT 766.500000 282.350000 799.500000 283.650000 ;
      RECT 757.500000 282.350000 758.500000 283.650000 ;
      RECT 716.500000 282.350000 749.500000 283.650000 ;
      RECT 707.500000 282.350000 708.500000 283.650000 ;
      RECT 666.500000 282.350000 699.500000 283.650000 ;
      RECT 657.500000 282.350000 658.500000 283.650000 ;
      RECT 616.500000 282.350000 649.500000 283.650000 ;
      RECT 607.500000 282.350000 608.500000 283.650000 ;
      RECT 566.500000 282.350000 599.500000 283.650000 ;
      RECT 557.500000 282.350000 558.500000 283.650000 ;
      RECT 516.500000 282.350000 549.500000 283.650000 ;
      RECT 507.500000 282.350000 508.500000 283.650000 ;
      RECT 466.500000 282.350000 499.500000 283.650000 ;
      RECT 457.500000 282.350000 458.500000 283.650000 ;
      RECT 416.500000 282.350000 449.500000 283.650000 ;
      RECT 407.500000 282.350000 408.500000 283.650000 ;
      RECT 366.500000 282.350000 399.500000 283.650000 ;
      RECT 357.500000 282.350000 358.500000 283.650000 ;
      RECT 316.500000 282.350000 349.500000 283.650000 ;
      RECT 307.500000 282.350000 308.500000 283.650000 ;
      RECT 266.500000 282.350000 299.500000 283.650000 ;
      RECT 257.500000 282.350000 258.500000 283.650000 ;
      RECT 216.500000 282.350000 249.500000 283.650000 ;
      RECT 207.500000 282.350000 208.500000 283.650000 ;
      RECT 166.500000 282.350000 199.500000 283.650000 ;
      RECT 157.500000 282.350000 158.500000 283.650000 ;
      RECT 116.500000 282.350000 149.500000 283.650000 ;
      RECT 107.500000 282.350000 108.500000 283.650000 ;
      RECT 66.500000 282.350000 99.500000 283.650000 ;
      RECT 57.500000 282.350000 58.500000 283.650000 ;
      RECT 29.500000 282.350000 49.500000 283.650000 ;
      RECT 15.500000 282.350000 16.500000 283.650000 ;
      RECT 1157.500000 281.650000 1170.500000 282.350000 ;
      RECT 1107.500000 281.650000 1149.500000 282.350000 ;
      RECT 1057.500000 281.650000 1099.500000 282.350000 ;
      RECT 1007.500000 281.650000 1049.500000 282.350000 ;
      RECT 957.500000 281.650000 999.500000 282.350000 ;
      RECT 907.500000 281.650000 949.500000 282.350000 ;
      RECT 857.500000 281.650000 899.500000 282.350000 ;
      RECT 807.500000 281.650000 849.500000 282.350000 ;
      RECT 757.500000 281.650000 799.500000 282.350000 ;
      RECT 707.500000 281.650000 749.500000 282.350000 ;
      RECT 657.500000 281.650000 699.500000 282.350000 ;
      RECT 607.500000 281.650000 649.500000 282.350000 ;
      RECT 557.500000 281.650000 599.500000 282.350000 ;
      RECT 507.500000 281.650000 549.500000 282.350000 ;
      RECT 457.500000 281.650000 499.500000 282.350000 ;
      RECT 407.500000 281.650000 449.500000 282.350000 ;
      RECT 357.500000 281.650000 399.500000 282.350000 ;
      RECT 307.500000 281.650000 349.500000 282.350000 ;
      RECT 257.500000 281.650000 299.500000 282.350000 ;
      RECT 207.500000 281.650000 249.500000 282.350000 ;
      RECT 157.500000 281.650000 199.500000 282.350000 ;
      RECT 107.500000 281.650000 149.500000 282.350000 ;
      RECT 57.500000 281.650000 99.500000 282.350000 ;
      RECT 15.500000 281.650000 49.500000 282.350000 ;
      RECT 1183.500000 280.350000 1186.000000 283.650000 ;
      RECT 1169.500000 280.350000 1170.500000 281.650000 ;
      RECT 1116.500000 280.350000 1149.500000 281.650000 ;
      RECT 1107.500000 280.350000 1108.500000 281.650000 ;
      RECT 1066.500000 280.350000 1099.500000 281.650000 ;
      RECT 1057.500000 280.350000 1058.500000 281.650000 ;
      RECT 1016.500000 280.350000 1049.500000 281.650000 ;
      RECT 1007.500000 280.350000 1008.500000 281.650000 ;
      RECT 966.500000 280.350000 999.500000 281.650000 ;
      RECT 957.500000 280.350000 958.500000 281.650000 ;
      RECT 916.500000 280.350000 949.500000 281.650000 ;
      RECT 907.500000 280.350000 908.500000 281.650000 ;
      RECT 866.500000 280.350000 899.500000 281.650000 ;
      RECT 857.500000 280.350000 858.500000 281.650000 ;
      RECT 816.500000 280.350000 849.500000 281.650000 ;
      RECT 807.500000 280.350000 808.500000 281.650000 ;
      RECT 766.500000 280.350000 799.500000 281.650000 ;
      RECT 757.500000 280.350000 758.500000 281.650000 ;
      RECT 716.500000 280.350000 749.500000 281.650000 ;
      RECT 707.500000 280.350000 708.500000 281.650000 ;
      RECT 666.500000 280.350000 699.500000 281.650000 ;
      RECT 657.500000 280.350000 658.500000 281.650000 ;
      RECT 616.500000 280.350000 649.500000 281.650000 ;
      RECT 607.500000 280.350000 608.500000 281.650000 ;
      RECT 566.500000 280.350000 599.500000 281.650000 ;
      RECT 557.500000 280.350000 558.500000 281.650000 ;
      RECT 516.500000 280.350000 549.500000 281.650000 ;
      RECT 507.500000 280.350000 508.500000 281.650000 ;
      RECT 466.500000 280.350000 499.500000 281.650000 ;
      RECT 457.500000 280.350000 458.500000 281.650000 ;
      RECT 416.500000 280.350000 449.500000 281.650000 ;
      RECT 407.500000 280.350000 408.500000 281.650000 ;
      RECT 366.500000 280.350000 399.500000 281.650000 ;
      RECT 357.500000 280.350000 358.500000 281.650000 ;
      RECT 316.500000 280.350000 349.500000 281.650000 ;
      RECT 307.500000 280.350000 308.500000 281.650000 ;
      RECT 266.500000 280.350000 299.500000 281.650000 ;
      RECT 257.500000 280.350000 258.500000 281.650000 ;
      RECT 216.500000 280.350000 249.500000 281.650000 ;
      RECT 207.500000 280.350000 208.500000 281.650000 ;
      RECT 166.500000 280.350000 199.500000 281.650000 ;
      RECT 157.500000 280.350000 158.500000 281.650000 ;
      RECT 116.500000 280.350000 149.500000 281.650000 ;
      RECT 107.500000 280.350000 108.500000 281.650000 ;
      RECT 66.500000 280.350000 99.500000 281.650000 ;
      RECT 57.500000 280.350000 58.500000 281.650000 ;
      RECT 29.500000 280.350000 49.500000 281.650000 ;
      RECT 15.500000 280.350000 16.500000 281.650000 ;
      RECT 0.000000 280.350000 2.500000 283.650000 ;
      RECT 1169.500000 279.650000 1186.000000 280.350000 ;
      RECT 1116.500000 279.650000 1156.500000 280.350000 ;
      RECT 1066.500000 279.650000 1108.500000 280.350000 ;
      RECT 1016.500000 279.650000 1058.500000 280.350000 ;
      RECT 966.500000 279.650000 1008.500000 280.350000 ;
      RECT 916.500000 279.650000 958.500000 280.350000 ;
      RECT 866.500000 279.650000 908.500000 280.350000 ;
      RECT 816.500000 279.650000 858.500000 280.350000 ;
      RECT 766.500000 279.650000 808.500000 280.350000 ;
      RECT 716.500000 279.650000 758.500000 280.350000 ;
      RECT 666.500000 279.650000 708.500000 280.350000 ;
      RECT 616.500000 279.650000 658.500000 280.350000 ;
      RECT 566.500000 279.650000 608.500000 280.350000 ;
      RECT 516.500000 279.650000 558.500000 280.350000 ;
      RECT 466.500000 279.650000 508.500000 280.350000 ;
      RECT 416.500000 279.650000 458.500000 280.350000 ;
      RECT 366.500000 279.650000 408.500000 280.350000 ;
      RECT 316.500000 279.650000 358.500000 280.350000 ;
      RECT 266.500000 279.650000 308.500000 280.350000 ;
      RECT 216.500000 279.650000 258.500000 280.350000 ;
      RECT 166.500000 279.650000 208.500000 280.350000 ;
      RECT 116.500000 279.650000 158.500000 280.350000 ;
      RECT 66.500000 279.650000 108.500000 280.350000 ;
      RECT 29.500000 279.650000 58.500000 280.350000 ;
      RECT 0.000000 279.650000 16.500000 280.350000 ;
      RECT 1169.500000 278.350000 1170.500000 279.650000 ;
      RECT 1116.500000 278.350000 1149.500000 279.650000 ;
      RECT 1107.500000 278.350000 1108.500000 279.650000 ;
      RECT 1066.500000 278.350000 1099.500000 279.650000 ;
      RECT 1057.500000 278.350000 1058.500000 279.650000 ;
      RECT 1016.500000 278.350000 1049.500000 279.650000 ;
      RECT 1007.500000 278.350000 1008.500000 279.650000 ;
      RECT 966.500000 278.350000 999.500000 279.650000 ;
      RECT 957.500000 278.350000 958.500000 279.650000 ;
      RECT 916.500000 278.350000 949.500000 279.650000 ;
      RECT 907.500000 278.350000 908.500000 279.650000 ;
      RECT 866.500000 278.350000 899.500000 279.650000 ;
      RECT 857.500000 278.350000 858.500000 279.650000 ;
      RECT 816.500000 278.350000 849.500000 279.650000 ;
      RECT 807.500000 278.350000 808.500000 279.650000 ;
      RECT 766.500000 278.350000 799.500000 279.650000 ;
      RECT 757.500000 278.350000 758.500000 279.650000 ;
      RECT 716.500000 278.350000 749.500000 279.650000 ;
      RECT 707.500000 278.350000 708.500000 279.650000 ;
      RECT 666.500000 278.350000 699.500000 279.650000 ;
      RECT 657.500000 278.350000 658.500000 279.650000 ;
      RECT 616.500000 278.350000 649.500000 279.650000 ;
      RECT 607.500000 278.350000 608.500000 279.650000 ;
      RECT 566.500000 278.350000 599.500000 279.650000 ;
      RECT 557.500000 278.350000 558.500000 279.650000 ;
      RECT 516.500000 278.350000 549.500000 279.650000 ;
      RECT 507.500000 278.350000 508.500000 279.650000 ;
      RECT 466.500000 278.350000 499.500000 279.650000 ;
      RECT 457.500000 278.350000 458.500000 279.650000 ;
      RECT 416.500000 278.350000 449.500000 279.650000 ;
      RECT 407.500000 278.350000 408.500000 279.650000 ;
      RECT 366.500000 278.350000 399.500000 279.650000 ;
      RECT 357.500000 278.350000 358.500000 279.650000 ;
      RECT 316.500000 278.350000 349.500000 279.650000 ;
      RECT 307.500000 278.350000 308.500000 279.650000 ;
      RECT 266.500000 278.350000 299.500000 279.650000 ;
      RECT 257.500000 278.350000 258.500000 279.650000 ;
      RECT 216.500000 278.350000 249.500000 279.650000 ;
      RECT 207.500000 278.350000 208.500000 279.650000 ;
      RECT 166.500000 278.350000 199.500000 279.650000 ;
      RECT 157.500000 278.350000 158.500000 279.650000 ;
      RECT 116.500000 278.350000 149.500000 279.650000 ;
      RECT 107.500000 278.350000 108.500000 279.650000 ;
      RECT 66.500000 278.350000 99.500000 279.650000 ;
      RECT 57.500000 278.350000 58.500000 279.650000 ;
      RECT 29.500000 278.350000 49.500000 279.650000 ;
      RECT 15.500000 278.350000 16.500000 279.650000 ;
      RECT 1157.500000 277.650000 1170.500000 278.350000 ;
      RECT 1107.500000 277.650000 1149.500000 278.350000 ;
      RECT 1057.500000 277.650000 1099.500000 278.350000 ;
      RECT 1007.500000 277.650000 1049.500000 278.350000 ;
      RECT 957.500000 277.650000 999.500000 278.350000 ;
      RECT 907.500000 277.650000 949.500000 278.350000 ;
      RECT 857.500000 277.650000 899.500000 278.350000 ;
      RECT 807.500000 277.650000 849.500000 278.350000 ;
      RECT 757.500000 277.650000 799.500000 278.350000 ;
      RECT 707.500000 277.650000 749.500000 278.350000 ;
      RECT 657.500000 277.650000 699.500000 278.350000 ;
      RECT 607.500000 277.650000 649.500000 278.350000 ;
      RECT 557.500000 277.650000 599.500000 278.350000 ;
      RECT 507.500000 277.650000 549.500000 278.350000 ;
      RECT 457.500000 277.650000 499.500000 278.350000 ;
      RECT 407.500000 277.650000 449.500000 278.350000 ;
      RECT 357.500000 277.650000 399.500000 278.350000 ;
      RECT 307.500000 277.650000 349.500000 278.350000 ;
      RECT 257.500000 277.650000 299.500000 278.350000 ;
      RECT 207.500000 277.650000 249.500000 278.350000 ;
      RECT 157.500000 277.650000 199.500000 278.350000 ;
      RECT 107.500000 277.650000 149.500000 278.350000 ;
      RECT 57.500000 277.650000 99.500000 278.350000 ;
      RECT 15.500000 277.650000 49.500000 278.350000 ;
      RECT 1183.500000 276.350000 1186.000000 279.650000 ;
      RECT 1169.500000 276.350000 1170.500000 277.650000 ;
      RECT 1116.500000 276.350000 1149.500000 277.650000 ;
      RECT 1107.500000 276.350000 1108.500000 277.650000 ;
      RECT 1066.500000 276.350000 1099.500000 277.650000 ;
      RECT 1057.500000 276.350000 1058.500000 277.650000 ;
      RECT 1016.500000 276.350000 1049.500000 277.650000 ;
      RECT 1007.500000 276.350000 1008.500000 277.650000 ;
      RECT 966.500000 276.350000 999.500000 277.650000 ;
      RECT 957.500000 276.350000 958.500000 277.650000 ;
      RECT 916.500000 276.350000 949.500000 277.650000 ;
      RECT 907.500000 276.350000 908.500000 277.650000 ;
      RECT 866.500000 276.350000 899.500000 277.650000 ;
      RECT 857.500000 276.350000 858.500000 277.650000 ;
      RECT 816.500000 276.350000 849.500000 277.650000 ;
      RECT 807.500000 276.350000 808.500000 277.650000 ;
      RECT 766.500000 276.350000 799.500000 277.650000 ;
      RECT 757.500000 276.350000 758.500000 277.650000 ;
      RECT 716.500000 276.350000 749.500000 277.650000 ;
      RECT 707.500000 276.350000 708.500000 277.650000 ;
      RECT 666.500000 276.350000 699.500000 277.650000 ;
      RECT 657.500000 276.350000 658.500000 277.650000 ;
      RECT 616.500000 276.350000 649.500000 277.650000 ;
      RECT 607.500000 276.350000 608.500000 277.650000 ;
      RECT 566.500000 276.350000 599.500000 277.650000 ;
      RECT 557.500000 276.350000 558.500000 277.650000 ;
      RECT 516.500000 276.350000 549.500000 277.650000 ;
      RECT 507.500000 276.350000 508.500000 277.650000 ;
      RECT 466.500000 276.350000 499.500000 277.650000 ;
      RECT 457.500000 276.350000 458.500000 277.650000 ;
      RECT 416.500000 276.350000 449.500000 277.650000 ;
      RECT 407.500000 276.350000 408.500000 277.650000 ;
      RECT 366.500000 276.350000 399.500000 277.650000 ;
      RECT 357.500000 276.350000 358.500000 277.650000 ;
      RECT 316.500000 276.350000 349.500000 277.650000 ;
      RECT 307.500000 276.350000 308.500000 277.650000 ;
      RECT 266.500000 276.350000 299.500000 277.650000 ;
      RECT 257.500000 276.350000 258.500000 277.650000 ;
      RECT 216.500000 276.350000 249.500000 277.650000 ;
      RECT 207.500000 276.350000 208.500000 277.650000 ;
      RECT 166.500000 276.350000 199.500000 277.650000 ;
      RECT 157.500000 276.350000 158.500000 277.650000 ;
      RECT 116.500000 276.350000 149.500000 277.650000 ;
      RECT 107.500000 276.350000 108.500000 277.650000 ;
      RECT 66.500000 276.350000 99.500000 277.650000 ;
      RECT 57.500000 276.350000 58.500000 277.650000 ;
      RECT 29.500000 276.350000 49.500000 277.650000 ;
      RECT 15.500000 276.350000 16.500000 277.650000 ;
      RECT 0.000000 276.350000 2.500000 279.650000 ;
      RECT 1169.500000 275.650000 1186.000000 276.350000 ;
      RECT 1116.500000 275.650000 1156.500000 276.350000 ;
      RECT 1066.500000 275.650000 1108.500000 276.350000 ;
      RECT 1016.500000 275.650000 1058.500000 276.350000 ;
      RECT 966.500000 275.650000 1008.500000 276.350000 ;
      RECT 916.500000 275.650000 958.500000 276.350000 ;
      RECT 866.500000 275.650000 908.500000 276.350000 ;
      RECT 816.500000 275.650000 858.500000 276.350000 ;
      RECT 766.500000 275.650000 808.500000 276.350000 ;
      RECT 716.500000 275.650000 758.500000 276.350000 ;
      RECT 666.500000 275.650000 708.500000 276.350000 ;
      RECT 616.500000 275.650000 658.500000 276.350000 ;
      RECT 566.500000 275.650000 608.500000 276.350000 ;
      RECT 516.500000 275.650000 558.500000 276.350000 ;
      RECT 466.500000 275.650000 508.500000 276.350000 ;
      RECT 416.500000 275.650000 458.500000 276.350000 ;
      RECT 366.500000 275.650000 408.500000 276.350000 ;
      RECT 316.500000 275.650000 358.500000 276.350000 ;
      RECT 266.500000 275.650000 308.500000 276.350000 ;
      RECT 216.500000 275.650000 258.500000 276.350000 ;
      RECT 166.500000 275.650000 208.500000 276.350000 ;
      RECT 116.500000 275.650000 158.500000 276.350000 ;
      RECT 66.500000 275.650000 108.500000 276.350000 ;
      RECT 29.500000 275.650000 58.500000 276.350000 ;
      RECT 0.000000 275.650000 16.500000 276.350000 ;
      RECT 1169.500000 274.350000 1170.500000 275.650000 ;
      RECT 1116.500000 274.350000 1149.500000 275.650000 ;
      RECT 1107.500000 274.350000 1108.500000 275.650000 ;
      RECT 1066.500000 274.350000 1099.500000 275.650000 ;
      RECT 1057.500000 274.350000 1058.500000 275.650000 ;
      RECT 1016.500000 274.350000 1049.500000 275.650000 ;
      RECT 1007.500000 274.350000 1008.500000 275.650000 ;
      RECT 966.500000 274.350000 999.500000 275.650000 ;
      RECT 957.500000 274.350000 958.500000 275.650000 ;
      RECT 916.500000 274.350000 949.500000 275.650000 ;
      RECT 907.500000 274.350000 908.500000 275.650000 ;
      RECT 866.500000 274.350000 899.500000 275.650000 ;
      RECT 857.500000 274.350000 858.500000 275.650000 ;
      RECT 816.500000 274.350000 849.500000 275.650000 ;
      RECT 807.500000 274.350000 808.500000 275.650000 ;
      RECT 766.500000 274.350000 799.500000 275.650000 ;
      RECT 757.500000 274.350000 758.500000 275.650000 ;
      RECT 716.500000 274.350000 749.500000 275.650000 ;
      RECT 707.500000 274.350000 708.500000 275.650000 ;
      RECT 666.500000 274.350000 699.500000 275.650000 ;
      RECT 657.500000 274.350000 658.500000 275.650000 ;
      RECT 616.500000 274.350000 649.500000 275.650000 ;
      RECT 607.500000 274.350000 608.500000 275.650000 ;
      RECT 566.500000 274.350000 599.500000 275.650000 ;
      RECT 557.500000 274.350000 558.500000 275.650000 ;
      RECT 516.500000 274.350000 549.500000 275.650000 ;
      RECT 507.500000 274.350000 508.500000 275.650000 ;
      RECT 466.500000 274.350000 499.500000 275.650000 ;
      RECT 457.500000 274.350000 458.500000 275.650000 ;
      RECT 416.500000 274.350000 449.500000 275.650000 ;
      RECT 407.500000 274.350000 408.500000 275.650000 ;
      RECT 366.500000 274.350000 399.500000 275.650000 ;
      RECT 357.500000 274.350000 358.500000 275.650000 ;
      RECT 316.500000 274.350000 349.500000 275.650000 ;
      RECT 307.500000 274.350000 308.500000 275.650000 ;
      RECT 266.500000 274.350000 299.500000 275.650000 ;
      RECT 257.500000 274.350000 258.500000 275.650000 ;
      RECT 216.500000 274.350000 249.500000 275.650000 ;
      RECT 207.500000 274.350000 208.500000 275.650000 ;
      RECT 166.500000 274.350000 199.500000 275.650000 ;
      RECT 157.500000 274.350000 158.500000 275.650000 ;
      RECT 116.500000 274.350000 149.500000 275.650000 ;
      RECT 107.500000 274.350000 108.500000 275.650000 ;
      RECT 66.500000 274.350000 99.500000 275.650000 ;
      RECT 57.500000 274.350000 58.500000 275.650000 ;
      RECT 29.500000 274.350000 49.500000 275.650000 ;
      RECT 15.500000 274.350000 16.500000 275.650000 ;
      RECT 1157.500000 273.650000 1170.500000 274.350000 ;
      RECT 1107.500000 273.650000 1149.500000 274.350000 ;
      RECT 1057.500000 273.650000 1099.500000 274.350000 ;
      RECT 1007.500000 273.650000 1049.500000 274.350000 ;
      RECT 957.500000 273.650000 999.500000 274.350000 ;
      RECT 907.500000 273.650000 949.500000 274.350000 ;
      RECT 857.500000 273.650000 899.500000 274.350000 ;
      RECT 807.500000 273.650000 849.500000 274.350000 ;
      RECT 757.500000 273.650000 799.500000 274.350000 ;
      RECT 707.500000 273.650000 749.500000 274.350000 ;
      RECT 657.500000 273.650000 699.500000 274.350000 ;
      RECT 607.500000 273.650000 649.500000 274.350000 ;
      RECT 557.500000 273.650000 599.500000 274.350000 ;
      RECT 507.500000 273.650000 549.500000 274.350000 ;
      RECT 457.500000 273.650000 499.500000 274.350000 ;
      RECT 407.500000 273.650000 449.500000 274.350000 ;
      RECT 357.500000 273.650000 399.500000 274.350000 ;
      RECT 307.500000 273.650000 349.500000 274.350000 ;
      RECT 257.500000 273.650000 299.500000 274.350000 ;
      RECT 207.500000 273.650000 249.500000 274.350000 ;
      RECT 157.500000 273.650000 199.500000 274.350000 ;
      RECT 107.500000 273.650000 149.500000 274.350000 ;
      RECT 57.500000 273.650000 99.500000 274.350000 ;
      RECT 15.500000 273.650000 49.500000 274.350000 ;
      RECT 1183.500000 272.350000 1186.000000 275.650000 ;
      RECT 1169.500000 272.350000 1170.500000 273.650000 ;
      RECT 1116.500000 272.350000 1149.500000 273.650000 ;
      RECT 1107.500000 272.350000 1108.500000 273.650000 ;
      RECT 1066.500000 272.350000 1099.500000 273.650000 ;
      RECT 1057.500000 272.350000 1058.500000 273.650000 ;
      RECT 1016.500000 272.350000 1049.500000 273.650000 ;
      RECT 1007.500000 272.350000 1008.500000 273.650000 ;
      RECT 966.500000 272.350000 999.500000 273.650000 ;
      RECT 957.500000 272.350000 958.500000 273.650000 ;
      RECT 916.500000 272.350000 949.500000 273.650000 ;
      RECT 907.500000 272.350000 908.500000 273.650000 ;
      RECT 866.500000 272.350000 899.500000 273.650000 ;
      RECT 857.500000 272.350000 858.500000 273.650000 ;
      RECT 816.500000 272.350000 849.500000 273.650000 ;
      RECT 807.500000 272.350000 808.500000 273.650000 ;
      RECT 766.500000 272.350000 799.500000 273.650000 ;
      RECT 757.500000 272.350000 758.500000 273.650000 ;
      RECT 716.500000 272.350000 749.500000 273.650000 ;
      RECT 707.500000 272.350000 708.500000 273.650000 ;
      RECT 666.500000 272.350000 699.500000 273.650000 ;
      RECT 657.500000 272.350000 658.500000 273.650000 ;
      RECT 616.500000 272.350000 649.500000 273.650000 ;
      RECT 607.500000 272.350000 608.500000 273.650000 ;
      RECT 566.500000 272.350000 599.500000 273.650000 ;
      RECT 557.500000 272.350000 558.500000 273.650000 ;
      RECT 516.500000 272.350000 549.500000 273.650000 ;
      RECT 507.500000 272.350000 508.500000 273.650000 ;
      RECT 466.500000 272.350000 499.500000 273.650000 ;
      RECT 457.500000 272.350000 458.500000 273.650000 ;
      RECT 416.500000 272.350000 449.500000 273.650000 ;
      RECT 407.500000 272.350000 408.500000 273.650000 ;
      RECT 366.500000 272.350000 399.500000 273.650000 ;
      RECT 357.500000 272.350000 358.500000 273.650000 ;
      RECT 316.500000 272.350000 349.500000 273.650000 ;
      RECT 307.500000 272.350000 308.500000 273.650000 ;
      RECT 266.500000 272.350000 299.500000 273.650000 ;
      RECT 257.500000 272.350000 258.500000 273.650000 ;
      RECT 216.500000 272.350000 249.500000 273.650000 ;
      RECT 207.500000 272.350000 208.500000 273.650000 ;
      RECT 166.500000 272.350000 199.500000 273.650000 ;
      RECT 157.500000 272.350000 158.500000 273.650000 ;
      RECT 116.500000 272.350000 149.500000 273.650000 ;
      RECT 107.500000 272.350000 108.500000 273.650000 ;
      RECT 66.500000 272.350000 99.500000 273.650000 ;
      RECT 57.500000 272.350000 58.500000 273.650000 ;
      RECT 29.500000 272.350000 49.500000 273.650000 ;
      RECT 15.500000 272.350000 16.500000 273.650000 ;
      RECT 0.000000 272.350000 2.500000 275.650000 ;
      RECT 1169.500000 271.650000 1186.000000 272.350000 ;
      RECT 1116.500000 271.650000 1156.500000 272.350000 ;
      RECT 1066.500000 271.650000 1108.500000 272.350000 ;
      RECT 1016.500000 271.650000 1058.500000 272.350000 ;
      RECT 966.500000 271.650000 1008.500000 272.350000 ;
      RECT 916.500000 271.650000 958.500000 272.350000 ;
      RECT 866.500000 271.650000 908.500000 272.350000 ;
      RECT 816.500000 271.650000 858.500000 272.350000 ;
      RECT 766.500000 271.650000 808.500000 272.350000 ;
      RECT 716.500000 271.650000 758.500000 272.350000 ;
      RECT 666.500000 271.650000 708.500000 272.350000 ;
      RECT 616.500000 271.650000 658.500000 272.350000 ;
      RECT 566.500000 271.650000 608.500000 272.350000 ;
      RECT 516.500000 271.650000 558.500000 272.350000 ;
      RECT 466.500000 271.650000 508.500000 272.350000 ;
      RECT 416.500000 271.650000 458.500000 272.350000 ;
      RECT 366.500000 271.650000 408.500000 272.350000 ;
      RECT 316.500000 271.650000 358.500000 272.350000 ;
      RECT 266.500000 271.650000 308.500000 272.350000 ;
      RECT 216.500000 271.650000 258.500000 272.350000 ;
      RECT 166.500000 271.650000 208.500000 272.350000 ;
      RECT 116.500000 271.650000 158.500000 272.350000 ;
      RECT 66.500000 271.650000 108.500000 272.350000 ;
      RECT 29.500000 271.650000 58.500000 272.350000 ;
      RECT 0.000000 271.650000 16.500000 272.350000 ;
      RECT 1169.500000 270.350000 1170.500000 271.650000 ;
      RECT 1116.500000 270.350000 1149.500000 271.650000 ;
      RECT 1107.500000 270.350000 1108.500000 271.650000 ;
      RECT 1066.500000 270.350000 1099.500000 271.650000 ;
      RECT 1057.500000 270.350000 1058.500000 271.650000 ;
      RECT 1016.500000 270.350000 1049.500000 271.650000 ;
      RECT 1007.500000 270.350000 1008.500000 271.650000 ;
      RECT 966.500000 270.350000 999.500000 271.650000 ;
      RECT 957.500000 270.350000 958.500000 271.650000 ;
      RECT 916.500000 270.350000 949.500000 271.650000 ;
      RECT 907.500000 270.350000 908.500000 271.650000 ;
      RECT 866.500000 270.350000 899.500000 271.650000 ;
      RECT 857.500000 270.350000 858.500000 271.650000 ;
      RECT 816.500000 270.350000 849.500000 271.650000 ;
      RECT 807.500000 270.350000 808.500000 271.650000 ;
      RECT 766.500000 270.350000 799.500000 271.650000 ;
      RECT 757.500000 270.350000 758.500000 271.650000 ;
      RECT 716.500000 270.350000 749.500000 271.650000 ;
      RECT 707.500000 270.350000 708.500000 271.650000 ;
      RECT 666.500000 270.350000 699.500000 271.650000 ;
      RECT 657.500000 270.350000 658.500000 271.650000 ;
      RECT 616.500000 270.350000 649.500000 271.650000 ;
      RECT 607.500000 270.350000 608.500000 271.650000 ;
      RECT 566.500000 270.350000 599.500000 271.650000 ;
      RECT 557.500000 270.350000 558.500000 271.650000 ;
      RECT 516.500000 270.350000 549.500000 271.650000 ;
      RECT 507.500000 270.350000 508.500000 271.650000 ;
      RECT 466.500000 270.350000 499.500000 271.650000 ;
      RECT 457.500000 270.350000 458.500000 271.650000 ;
      RECT 416.500000 270.350000 449.500000 271.650000 ;
      RECT 407.500000 270.350000 408.500000 271.650000 ;
      RECT 366.500000 270.350000 399.500000 271.650000 ;
      RECT 357.500000 270.350000 358.500000 271.650000 ;
      RECT 316.500000 270.350000 349.500000 271.650000 ;
      RECT 307.500000 270.350000 308.500000 271.650000 ;
      RECT 266.500000 270.350000 299.500000 271.650000 ;
      RECT 257.500000 270.350000 258.500000 271.650000 ;
      RECT 216.500000 270.350000 249.500000 271.650000 ;
      RECT 207.500000 270.350000 208.500000 271.650000 ;
      RECT 166.500000 270.350000 199.500000 271.650000 ;
      RECT 157.500000 270.350000 158.500000 271.650000 ;
      RECT 116.500000 270.350000 149.500000 271.650000 ;
      RECT 107.500000 270.350000 108.500000 271.650000 ;
      RECT 66.500000 270.350000 99.500000 271.650000 ;
      RECT 57.500000 270.350000 58.500000 271.650000 ;
      RECT 29.500000 270.350000 49.500000 271.650000 ;
      RECT 15.500000 270.350000 16.500000 271.650000 ;
      RECT 1157.500000 269.650000 1170.500000 270.350000 ;
      RECT 1107.500000 269.650000 1149.500000 270.350000 ;
      RECT 1057.500000 269.650000 1099.500000 270.350000 ;
      RECT 1007.500000 269.650000 1049.500000 270.350000 ;
      RECT 957.500000 269.650000 999.500000 270.350000 ;
      RECT 907.500000 269.650000 949.500000 270.350000 ;
      RECT 857.500000 269.650000 899.500000 270.350000 ;
      RECT 807.500000 269.650000 849.500000 270.350000 ;
      RECT 757.500000 269.650000 799.500000 270.350000 ;
      RECT 707.500000 269.650000 749.500000 270.350000 ;
      RECT 657.500000 269.650000 699.500000 270.350000 ;
      RECT 607.500000 269.650000 649.500000 270.350000 ;
      RECT 557.500000 269.650000 599.500000 270.350000 ;
      RECT 507.500000 269.650000 549.500000 270.350000 ;
      RECT 457.500000 269.650000 499.500000 270.350000 ;
      RECT 407.500000 269.650000 449.500000 270.350000 ;
      RECT 357.500000 269.650000 399.500000 270.350000 ;
      RECT 307.500000 269.650000 349.500000 270.350000 ;
      RECT 257.500000 269.650000 299.500000 270.350000 ;
      RECT 207.500000 269.650000 249.500000 270.350000 ;
      RECT 157.500000 269.650000 199.500000 270.350000 ;
      RECT 107.500000 269.650000 149.500000 270.350000 ;
      RECT 57.500000 269.650000 99.500000 270.350000 ;
      RECT 15.500000 269.650000 49.500000 270.350000 ;
      RECT 1183.500000 268.350000 1186.000000 271.650000 ;
      RECT 1169.500000 268.350000 1170.500000 269.650000 ;
      RECT 1116.500000 268.350000 1149.500000 269.650000 ;
      RECT 1107.500000 268.350000 1108.500000 269.650000 ;
      RECT 1066.500000 268.350000 1099.500000 269.650000 ;
      RECT 1057.500000 268.350000 1058.500000 269.650000 ;
      RECT 1016.500000 268.350000 1049.500000 269.650000 ;
      RECT 1007.500000 268.350000 1008.500000 269.650000 ;
      RECT 966.500000 268.350000 999.500000 269.650000 ;
      RECT 957.500000 268.350000 958.500000 269.650000 ;
      RECT 916.500000 268.350000 949.500000 269.650000 ;
      RECT 907.500000 268.350000 908.500000 269.650000 ;
      RECT 866.500000 268.350000 899.500000 269.650000 ;
      RECT 857.500000 268.350000 858.500000 269.650000 ;
      RECT 816.500000 268.350000 849.500000 269.650000 ;
      RECT 807.500000 268.350000 808.500000 269.650000 ;
      RECT 766.500000 268.350000 799.500000 269.650000 ;
      RECT 757.500000 268.350000 758.500000 269.650000 ;
      RECT 716.500000 268.350000 749.500000 269.650000 ;
      RECT 707.500000 268.350000 708.500000 269.650000 ;
      RECT 666.500000 268.350000 699.500000 269.650000 ;
      RECT 657.500000 268.350000 658.500000 269.650000 ;
      RECT 616.500000 268.350000 649.500000 269.650000 ;
      RECT 607.500000 268.350000 608.500000 269.650000 ;
      RECT 566.500000 268.350000 599.500000 269.650000 ;
      RECT 557.500000 268.350000 558.500000 269.650000 ;
      RECT 516.500000 268.350000 549.500000 269.650000 ;
      RECT 507.500000 268.350000 508.500000 269.650000 ;
      RECT 466.500000 268.350000 499.500000 269.650000 ;
      RECT 457.500000 268.350000 458.500000 269.650000 ;
      RECT 416.500000 268.350000 449.500000 269.650000 ;
      RECT 407.500000 268.350000 408.500000 269.650000 ;
      RECT 366.500000 268.350000 399.500000 269.650000 ;
      RECT 357.500000 268.350000 358.500000 269.650000 ;
      RECT 316.500000 268.350000 349.500000 269.650000 ;
      RECT 307.500000 268.350000 308.500000 269.650000 ;
      RECT 266.500000 268.350000 299.500000 269.650000 ;
      RECT 257.500000 268.350000 258.500000 269.650000 ;
      RECT 216.500000 268.350000 249.500000 269.650000 ;
      RECT 207.500000 268.350000 208.500000 269.650000 ;
      RECT 166.500000 268.350000 199.500000 269.650000 ;
      RECT 157.500000 268.350000 158.500000 269.650000 ;
      RECT 116.500000 268.350000 149.500000 269.650000 ;
      RECT 107.500000 268.350000 108.500000 269.650000 ;
      RECT 66.500000 268.350000 99.500000 269.650000 ;
      RECT 57.500000 268.350000 58.500000 269.650000 ;
      RECT 29.500000 268.350000 49.500000 269.650000 ;
      RECT 15.500000 268.350000 16.500000 269.650000 ;
      RECT 0.000000 268.350000 2.500000 271.650000 ;
      RECT 1169.500000 267.650000 1186.000000 268.350000 ;
      RECT 1116.500000 267.650000 1156.500000 268.350000 ;
      RECT 1066.500000 267.650000 1108.500000 268.350000 ;
      RECT 1016.500000 267.650000 1058.500000 268.350000 ;
      RECT 966.500000 267.650000 1008.500000 268.350000 ;
      RECT 916.500000 267.650000 958.500000 268.350000 ;
      RECT 866.500000 267.650000 908.500000 268.350000 ;
      RECT 816.500000 267.650000 858.500000 268.350000 ;
      RECT 766.500000 267.650000 808.500000 268.350000 ;
      RECT 716.500000 267.650000 758.500000 268.350000 ;
      RECT 666.500000 267.650000 708.500000 268.350000 ;
      RECT 616.500000 267.650000 658.500000 268.350000 ;
      RECT 566.500000 267.650000 608.500000 268.350000 ;
      RECT 516.500000 267.650000 558.500000 268.350000 ;
      RECT 466.500000 267.650000 508.500000 268.350000 ;
      RECT 416.500000 267.650000 458.500000 268.350000 ;
      RECT 366.500000 267.650000 408.500000 268.350000 ;
      RECT 316.500000 267.650000 358.500000 268.350000 ;
      RECT 266.500000 267.650000 308.500000 268.350000 ;
      RECT 216.500000 267.650000 258.500000 268.350000 ;
      RECT 166.500000 267.650000 208.500000 268.350000 ;
      RECT 116.500000 267.650000 158.500000 268.350000 ;
      RECT 66.500000 267.650000 108.500000 268.350000 ;
      RECT 29.500000 267.650000 58.500000 268.350000 ;
      RECT 0.000000 267.650000 16.500000 268.350000 ;
      RECT 1169.500000 266.350000 1170.500000 267.650000 ;
      RECT 1116.500000 266.350000 1149.500000 267.650000 ;
      RECT 1107.500000 266.350000 1108.500000 267.650000 ;
      RECT 1066.500000 266.350000 1099.500000 267.650000 ;
      RECT 1057.500000 266.350000 1058.500000 267.650000 ;
      RECT 1016.500000 266.350000 1049.500000 267.650000 ;
      RECT 1007.500000 266.350000 1008.500000 267.650000 ;
      RECT 966.500000 266.350000 999.500000 267.650000 ;
      RECT 957.500000 266.350000 958.500000 267.650000 ;
      RECT 916.500000 266.350000 949.500000 267.650000 ;
      RECT 907.500000 266.350000 908.500000 267.650000 ;
      RECT 866.500000 266.350000 899.500000 267.650000 ;
      RECT 857.500000 266.350000 858.500000 267.650000 ;
      RECT 816.500000 266.350000 849.500000 267.650000 ;
      RECT 807.500000 266.350000 808.500000 267.650000 ;
      RECT 766.500000 266.350000 799.500000 267.650000 ;
      RECT 757.500000 266.350000 758.500000 267.650000 ;
      RECT 716.500000 266.350000 749.500000 267.650000 ;
      RECT 707.500000 266.350000 708.500000 267.650000 ;
      RECT 666.500000 266.350000 699.500000 267.650000 ;
      RECT 657.500000 266.350000 658.500000 267.650000 ;
      RECT 616.500000 266.350000 649.500000 267.650000 ;
      RECT 607.500000 266.350000 608.500000 267.650000 ;
      RECT 566.500000 266.350000 599.500000 267.650000 ;
      RECT 557.500000 266.350000 558.500000 267.650000 ;
      RECT 516.500000 266.350000 549.500000 267.650000 ;
      RECT 507.500000 266.350000 508.500000 267.650000 ;
      RECT 466.500000 266.350000 499.500000 267.650000 ;
      RECT 457.500000 266.350000 458.500000 267.650000 ;
      RECT 416.500000 266.350000 449.500000 267.650000 ;
      RECT 407.500000 266.350000 408.500000 267.650000 ;
      RECT 366.500000 266.350000 399.500000 267.650000 ;
      RECT 357.500000 266.350000 358.500000 267.650000 ;
      RECT 316.500000 266.350000 349.500000 267.650000 ;
      RECT 307.500000 266.350000 308.500000 267.650000 ;
      RECT 266.500000 266.350000 299.500000 267.650000 ;
      RECT 257.500000 266.350000 258.500000 267.650000 ;
      RECT 216.500000 266.350000 249.500000 267.650000 ;
      RECT 207.500000 266.350000 208.500000 267.650000 ;
      RECT 166.500000 266.350000 199.500000 267.650000 ;
      RECT 157.500000 266.350000 158.500000 267.650000 ;
      RECT 116.500000 266.350000 149.500000 267.650000 ;
      RECT 107.500000 266.350000 108.500000 267.650000 ;
      RECT 66.500000 266.350000 99.500000 267.650000 ;
      RECT 57.500000 266.350000 58.500000 267.650000 ;
      RECT 29.500000 266.350000 49.500000 267.650000 ;
      RECT 15.500000 266.350000 16.500000 267.650000 ;
      RECT 1157.500000 265.650000 1170.500000 266.350000 ;
      RECT 1107.500000 265.650000 1149.500000 266.350000 ;
      RECT 1057.500000 265.650000 1099.500000 266.350000 ;
      RECT 1007.500000 265.650000 1049.500000 266.350000 ;
      RECT 957.500000 265.650000 999.500000 266.350000 ;
      RECT 907.500000 265.650000 949.500000 266.350000 ;
      RECT 857.500000 265.650000 899.500000 266.350000 ;
      RECT 807.500000 265.650000 849.500000 266.350000 ;
      RECT 757.500000 265.650000 799.500000 266.350000 ;
      RECT 707.500000 265.650000 749.500000 266.350000 ;
      RECT 657.500000 265.650000 699.500000 266.350000 ;
      RECT 607.500000 265.650000 649.500000 266.350000 ;
      RECT 557.500000 265.650000 599.500000 266.350000 ;
      RECT 507.500000 265.650000 549.500000 266.350000 ;
      RECT 457.500000 265.650000 499.500000 266.350000 ;
      RECT 407.500000 265.650000 449.500000 266.350000 ;
      RECT 357.500000 265.650000 399.500000 266.350000 ;
      RECT 307.500000 265.650000 349.500000 266.350000 ;
      RECT 257.500000 265.650000 299.500000 266.350000 ;
      RECT 207.500000 265.650000 249.500000 266.350000 ;
      RECT 157.500000 265.650000 199.500000 266.350000 ;
      RECT 107.500000 265.650000 149.500000 266.350000 ;
      RECT 57.500000 265.650000 99.500000 266.350000 ;
      RECT 15.500000 265.650000 49.500000 266.350000 ;
      RECT 1183.500000 264.350000 1186.000000 267.650000 ;
      RECT 1169.500000 264.350000 1170.500000 265.650000 ;
      RECT 1116.500000 264.350000 1149.500000 265.650000 ;
      RECT 1107.500000 264.350000 1108.500000 265.650000 ;
      RECT 1066.500000 264.350000 1099.500000 265.650000 ;
      RECT 1057.500000 264.350000 1058.500000 265.650000 ;
      RECT 1016.500000 264.350000 1049.500000 265.650000 ;
      RECT 1007.500000 264.350000 1008.500000 265.650000 ;
      RECT 966.500000 264.350000 999.500000 265.650000 ;
      RECT 957.500000 264.350000 958.500000 265.650000 ;
      RECT 916.500000 264.350000 949.500000 265.650000 ;
      RECT 907.500000 264.350000 908.500000 265.650000 ;
      RECT 866.500000 264.350000 899.500000 265.650000 ;
      RECT 857.500000 264.350000 858.500000 265.650000 ;
      RECT 816.500000 264.350000 849.500000 265.650000 ;
      RECT 807.500000 264.350000 808.500000 265.650000 ;
      RECT 766.500000 264.350000 799.500000 265.650000 ;
      RECT 757.500000 264.350000 758.500000 265.650000 ;
      RECT 716.500000 264.350000 749.500000 265.650000 ;
      RECT 707.500000 264.350000 708.500000 265.650000 ;
      RECT 666.500000 264.350000 699.500000 265.650000 ;
      RECT 657.500000 264.350000 658.500000 265.650000 ;
      RECT 616.500000 264.350000 649.500000 265.650000 ;
      RECT 607.500000 264.350000 608.500000 265.650000 ;
      RECT 566.500000 264.350000 599.500000 265.650000 ;
      RECT 557.500000 264.350000 558.500000 265.650000 ;
      RECT 516.500000 264.350000 549.500000 265.650000 ;
      RECT 507.500000 264.350000 508.500000 265.650000 ;
      RECT 466.500000 264.350000 499.500000 265.650000 ;
      RECT 457.500000 264.350000 458.500000 265.650000 ;
      RECT 416.500000 264.350000 449.500000 265.650000 ;
      RECT 407.500000 264.350000 408.500000 265.650000 ;
      RECT 366.500000 264.350000 399.500000 265.650000 ;
      RECT 357.500000 264.350000 358.500000 265.650000 ;
      RECT 316.500000 264.350000 349.500000 265.650000 ;
      RECT 307.500000 264.350000 308.500000 265.650000 ;
      RECT 266.500000 264.350000 299.500000 265.650000 ;
      RECT 257.500000 264.350000 258.500000 265.650000 ;
      RECT 216.500000 264.350000 249.500000 265.650000 ;
      RECT 207.500000 264.350000 208.500000 265.650000 ;
      RECT 166.500000 264.350000 199.500000 265.650000 ;
      RECT 157.500000 264.350000 158.500000 265.650000 ;
      RECT 116.500000 264.350000 149.500000 265.650000 ;
      RECT 107.500000 264.350000 108.500000 265.650000 ;
      RECT 66.500000 264.350000 99.500000 265.650000 ;
      RECT 57.500000 264.350000 58.500000 265.650000 ;
      RECT 29.500000 264.350000 49.500000 265.650000 ;
      RECT 15.500000 264.350000 16.500000 265.650000 ;
      RECT 0.000000 264.350000 2.500000 267.650000 ;
      RECT 1169.500000 263.650000 1186.000000 264.350000 ;
      RECT 1116.500000 263.650000 1156.500000 264.350000 ;
      RECT 1066.500000 263.650000 1108.500000 264.350000 ;
      RECT 1016.500000 263.650000 1058.500000 264.350000 ;
      RECT 966.500000 263.650000 1008.500000 264.350000 ;
      RECT 916.500000 263.650000 958.500000 264.350000 ;
      RECT 866.500000 263.650000 908.500000 264.350000 ;
      RECT 816.500000 263.650000 858.500000 264.350000 ;
      RECT 766.500000 263.650000 808.500000 264.350000 ;
      RECT 716.500000 263.650000 758.500000 264.350000 ;
      RECT 666.500000 263.650000 708.500000 264.350000 ;
      RECT 616.500000 263.650000 658.500000 264.350000 ;
      RECT 566.500000 263.650000 608.500000 264.350000 ;
      RECT 516.500000 263.650000 558.500000 264.350000 ;
      RECT 466.500000 263.650000 508.500000 264.350000 ;
      RECT 416.500000 263.650000 458.500000 264.350000 ;
      RECT 366.500000 263.650000 408.500000 264.350000 ;
      RECT 316.500000 263.650000 358.500000 264.350000 ;
      RECT 266.500000 263.650000 308.500000 264.350000 ;
      RECT 216.500000 263.650000 258.500000 264.350000 ;
      RECT 166.500000 263.650000 208.500000 264.350000 ;
      RECT 116.500000 263.650000 158.500000 264.350000 ;
      RECT 66.500000 263.650000 108.500000 264.350000 ;
      RECT 29.500000 263.650000 58.500000 264.350000 ;
      RECT 0.000000 263.650000 16.500000 264.350000 ;
      RECT 1169.500000 262.350000 1170.500000 263.650000 ;
      RECT 1116.500000 262.350000 1149.500000 263.650000 ;
      RECT 1107.500000 262.350000 1108.500000 263.650000 ;
      RECT 1066.500000 262.350000 1099.500000 263.650000 ;
      RECT 1057.500000 262.350000 1058.500000 263.650000 ;
      RECT 1016.500000 262.350000 1049.500000 263.650000 ;
      RECT 1007.500000 262.350000 1008.500000 263.650000 ;
      RECT 966.500000 262.350000 999.500000 263.650000 ;
      RECT 957.500000 262.350000 958.500000 263.650000 ;
      RECT 916.500000 262.350000 949.500000 263.650000 ;
      RECT 907.500000 262.350000 908.500000 263.650000 ;
      RECT 866.500000 262.350000 899.500000 263.650000 ;
      RECT 857.500000 262.350000 858.500000 263.650000 ;
      RECT 816.500000 262.350000 849.500000 263.650000 ;
      RECT 807.500000 262.350000 808.500000 263.650000 ;
      RECT 766.500000 262.350000 799.500000 263.650000 ;
      RECT 757.500000 262.350000 758.500000 263.650000 ;
      RECT 716.500000 262.350000 749.500000 263.650000 ;
      RECT 707.500000 262.350000 708.500000 263.650000 ;
      RECT 666.500000 262.350000 699.500000 263.650000 ;
      RECT 657.500000 262.350000 658.500000 263.650000 ;
      RECT 616.500000 262.350000 649.500000 263.650000 ;
      RECT 607.500000 262.350000 608.500000 263.650000 ;
      RECT 566.500000 262.350000 599.500000 263.650000 ;
      RECT 557.500000 262.350000 558.500000 263.650000 ;
      RECT 516.500000 262.350000 549.500000 263.650000 ;
      RECT 507.500000 262.350000 508.500000 263.650000 ;
      RECT 466.500000 262.350000 499.500000 263.650000 ;
      RECT 457.500000 262.350000 458.500000 263.650000 ;
      RECT 416.500000 262.350000 449.500000 263.650000 ;
      RECT 407.500000 262.350000 408.500000 263.650000 ;
      RECT 366.500000 262.350000 399.500000 263.650000 ;
      RECT 357.500000 262.350000 358.500000 263.650000 ;
      RECT 316.500000 262.350000 349.500000 263.650000 ;
      RECT 307.500000 262.350000 308.500000 263.650000 ;
      RECT 266.500000 262.350000 299.500000 263.650000 ;
      RECT 257.500000 262.350000 258.500000 263.650000 ;
      RECT 216.500000 262.350000 249.500000 263.650000 ;
      RECT 207.500000 262.350000 208.500000 263.650000 ;
      RECT 166.500000 262.350000 199.500000 263.650000 ;
      RECT 157.500000 262.350000 158.500000 263.650000 ;
      RECT 116.500000 262.350000 149.500000 263.650000 ;
      RECT 107.500000 262.350000 108.500000 263.650000 ;
      RECT 66.500000 262.350000 99.500000 263.650000 ;
      RECT 57.500000 262.350000 58.500000 263.650000 ;
      RECT 29.500000 262.350000 49.500000 263.650000 ;
      RECT 15.500000 262.350000 16.500000 263.650000 ;
      RECT 1157.500000 261.650000 1170.500000 262.350000 ;
      RECT 1107.500000 261.650000 1149.500000 262.350000 ;
      RECT 1057.500000 261.650000 1099.500000 262.350000 ;
      RECT 1007.500000 261.650000 1049.500000 262.350000 ;
      RECT 957.500000 261.650000 999.500000 262.350000 ;
      RECT 907.500000 261.650000 949.500000 262.350000 ;
      RECT 857.500000 261.650000 899.500000 262.350000 ;
      RECT 807.500000 261.650000 849.500000 262.350000 ;
      RECT 757.500000 261.650000 799.500000 262.350000 ;
      RECT 707.500000 261.650000 749.500000 262.350000 ;
      RECT 657.500000 261.650000 699.500000 262.350000 ;
      RECT 607.500000 261.650000 649.500000 262.350000 ;
      RECT 557.500000 261.650000 599.500000 262.350000 ;
      RECT 507.500000 261.650000 549.500000 262.350000 ;
      RECT 457.500000 261.650000 499.500000 262.350000 ;
      RECT 407.500000 261.650000 449.500000 262.350000 ;
      RECT 357.500000 261.650000 399.500000 262.350000 ;
      RECT 307.500000 261.650000 349.500000 262.350000 ;
      RECT 257.500000 261.650000 299.500000 262.350000 ;
      RECT 207.500000 261.650000 249.500000 262.350000 ;
      RECT 157.500000 261.650000 199.500000 262.350000 ;
      RECT 107.500000 261.650000 149.500000 262.350000 ;
      RECT 57.500000 261.650000 99.500000 262.350000 ;
      RECT 15.500000 261.650000 49.500000 262.350000 ;
      RECT 1183.500000 260.350000 1186.000000 263.650000 ;
      RECT 1169.500000 260.350000 1170.500000 261.650000 ;
      RECT 1116.500000 260.350000 1149.500000 261.650000 ;
      RECT 1107.500000 260.350000 1108.500000 261.650000 ;
      RECT 1066.500000 260.350000 1099.500000 261.650000 ;
      RECT 1057.500000 260.350000 1058.500000 261.650000 ;
      RECT 1016.500000 260.350000 1049.500000 261.650000 ;
      RECT 1007.500000 260.350000 1008.500000 261.650000 ;
      RECT 966.500000 260.350000 999.500000 261.650000 ;
      RECT 957.500000 260.350000 958.500000 261.650000 ;
      RECT 916.500000 260.350000 949.500000 261.650000 ;
      RECT 907.500000 260.350000 908.500000 261.650000 ;
      RECT 866.500000 260.350000 899.500000 261.650000 ;
      RECT 857.500000 260.350000 858.500000 261.650000 ;
      RECT 816.500000 260.350000 849.500000 261.650000 ;
      RECT 807.500000 260.350000 808.500000 261.650000 ;
      RECT 766.500000 260.350000 799.500000 261.650000 ;
      RECT 757.500000 260.350000 758.500000 261.650000 ;
      RECT 716.500000 260.350000 749.500000 261.650000 ;
      RECT 707.500000 260.350000 708.500000 261.650000 ;
      RECT 666.500000 260.350000 699.500000 261.650000 ;
      RECT 657.500000 260.350000 658.500000 261.650000 ;
      RECT 616.500000 260.350000 649.500000 261.650000 ;
      RECT 607.500000 260.350000 608.500000 261.650000 ;
      RECT 566.500000 260.350000 599.500000 261.650000 ;
      RECT 557.500000 260.350000 558.500000 261.650000 ;
      RECT 516.500000 260.350000 549.500000 261.650000 ;
      RECT 507.500000 260.350000 508.500000 261.650000 ;
      RECT 466.500000 260.350000 499.500000 261.650000 ;
      RECT 457.500000 260.350000 458.500000 261.650000 ;
      RECT 416.500000 260.350000 449.500000 261.650000 ;
      RECT 407.500000 260.350000 408.500000 261.650000 ;
      RECT 366.500000 260.350000 399.500000 261.650000 ;
      RECT 357.500000 260.350000 358.500000 261.650000 ;
      RECT 316.500000 260.350000 349.500000 261.650000 ;
      RECT 307.500000 260.350000 308.500000 261.650000 ;
      RECT 266.500000 260.350000 299.500000 261.650000 ;
      RECT 257.500000 260.350000 258.500000 261.650000 ;
      RECT 216.500000 260.350000 249.500000 261.650000 ;
      RECT 207.500000 260.350000 208.500000 261.650000 ;
      RECT 166.500000 260.350000 199.500000 261.650000 ;
      RECT 157.500000 260.350000 158.500000 261.650000 ;
      RECT 116.500000 260.350000 149.500000 261.650000 ;
      RECT 107.500000 260.350000 108.500000 261.650000 ;
      RECT 66.500000 260.350000 99.500000 261.650000 ;
      RECT 57.500000 260.350000 58.500000 261.650000 ;
      RECT 29.500000 260.350000 49.500000 261.650000 ;
      RECT 15.500000 260.350000 16.500000 261.650000 ;
      RECT 0.000000 260.350000 2.500000 263.650000 ;
      RECT 1169.500000 259.650000 1186.000000 260.350000 ;
      RECT 1116.500000 259.650000 1156.500000 260.350000 ;
      RECT 1169.500000 258.350000 1170.500000 259.650000 ;
      RECT 1116.500000 258.350000 1149.500000 259.650000 ;
      RECT 1066.500000 258.350000 1108.500000 260.350000 ;
      RECT 1016.500000 258.350000 1058.500000 260.350000 ;
      RECT 966.500000 258.350000 1008.500000 260.350000 ;
      RECT 916.500000 258.350000 958.500000 260.350000 ;
      RECT 866.500000 258.350000 908.500000 260.350000 ;
      RECT 816.500000 258.350000 858.500000 260.350000 ;
      RECT 766.500000 258.350000 808.500000 260.350000 ;
      RECT 716.500000 258.350000 758.500000 260.350000 ;
      RECT 666.500000 258.350000 708.500000 260.350000 ;
      RECT 616.500000 258.350000 658.500000 260.350000 ;
      RECT 566.500000 258.350000 608.500000 260.350000 ;
      RECT 516.500000 258.350000 558.500000 260.350000 ;
      RECT 466.500000 258.350000 508.500000 260.350000 ;
      RECT 416.500000 258.350000 458.500000 260.350000 ;
      RECT 366.500000 258.350000 408.500000 260.350000 ;
      RECT 316.500000 258.350000 358.500000 260.350000 ;
      RECT 266.500000 258.350000 308.500000 260.350000 ;
      RECT 216.500000 258.350000 258.500000 260.350000 ;
      RECT 166.500000 258.350000 208.500000 260.350000 ;
      RECT 116.500000 258.350000 158.500000 260.350000 ;
      RECT 66.500000 258.350000 108.500000 260.350000 ;
      RECT 29.500000 258.350000 58.500000 260.350000 ;
      RECT 0.000000 258.350000 16.500000 260.350000 ;
      RECT 1157.500000 257.650000 1170.500000 258.350000 ;
      RECT 1183.500000 256.350000 1186.000000 259.650000 ;
      RECT 1169.500000 256.350000 1170.500000 257.650000 ;
      RECT 0.000000 256.350000 1149.500000 258.350000 ;
      RECT 1169.500000 255.650000 1186.000000 256.350000 ;
      RECT 1169.500000 254.350000 1170.500000 255.650000 ;
      RECT 0.000000 254.350000 1156.500000 256.350000 ;
      RECT 0.000000 253.650000 1170.500000 254.350000 ;
      RECT 1183.500000 252.350000 1186.000000 255.650000 ;
      RECT 1169.500000 252.350000 1170.500000 253.650000 ;
      RECT 1169.500000 251.650000 1186.000000 252.350000 ;
      RECT 1169.500000 250.350000 1170.500000 251.650000 ;
      RECT 0.000000 250.350000 1156.500000 253.650000 ;
      RECT 0.000000 249.650000 1170.500000 250.350000 ;
      RECT 1183.500000 248.350000 1186.000000 251.650000 ;
      RECT 1169.500000 248.350000 1170.500000 249.650000 ;
      RECT 1169.500000 247.650000 1186.000000 248.350000 ;
      RECT 1169.500000 246.350000 1170.500000 247.650000 ;
      RECT 0.000000 246.350000 1156.500000 249.650000 ;
      RECT 0.000000 245.650000 1170.500000 246.350000 ;
      RECT 1183.500000 244.350000 1186.000000 247.650000 ;
      RECT 1169.500000 244.350000 1170.500000 245.650000 ;
      RECT 1169.500000 243.650000 1186.000000 244.350000 ;
      RECT 1169.500000 242.350000 1170.500000 243.650000 ;
      RECT 0.000000 242.350000 1156.500000 245.650000 ;
      RECT 0.000000 241.650000 1170.500000 242.350000 ;
      RECT 1183.500000 240.350000 1186.000000 243.650000 ;
      RECT 1169.500000 240.350000 1170.500000 241.650000 ;
      RECT 1169.500000 239.650000 1186.000000 240.350000 ;
      RECT 1169.500000 238.350000 1170.500000 239.650000 ;
      RECT 0.000000 238.350000 1156.500000 241.650000 ;
      RECT 0.000000 237.650000 1170.500000 238.350000 ;
      RECT 1183.500000 236.350000 1186.000000 239.650000 ;
      RECT 1169.500000 236.350000 1170.500000 237.650000 ;
      RECT 1169.500000 235.650000 1186.000000 236.350000 ;
      RECT 1169.500000 234.350000 1170.500000 235.650000 ;
      RECT 0.000000 234.350000 1156.500000 237.650000 ;
      RECT 0.000000 233.650000 1170.500000 234.350000 ;
      RECT 1183.500000 232.350000 1186.000000 235.650000 ;
      RECT 1169.500000 232.350000 1170.500000 233.650000 ;
      RECT 1169.500000 231.650000 1186.000000 232.350000 ;
      RECT 1169.500000 230.350000 1170.500000 231.650000 ;
      RECT 0.000000 230.350000 1156.500000 233.650000 ;
      RECT 0.000000 229.650000 1170.500000 230.350000 ;
      RECT 1183.500000 228.350000 1186.000000 231.650000 ;
      RECT 1169.500000 228.350000 1170.500000 229.650000 ;
      RECT 1169.500000 227.650000 1186.000000 228.350000 ;
      RECT 1169.500000 226.350000 1170.500000 227.650000 ;
      RECT 0.000000 226.350000 1156.500000 229.650000 ;
      RECT 0.000000 225.650000 1170.500000 226.350000 ;
      RECT 1183.500000 224.350000 1186.000000 227.650000 ;
      RECT 1169.500000 224.350000 1170.500000 225.650000 ;
      RECT 1169.500000 223.650000 1186.000000 224.350000 ;
      RECT 1169.500000 222.350000 1170.500000 223.650000 ;
      RECT 0.000000 222.350000 1156.500000 225.650000 ;
      RECT 0.000000 221.650000 1170.500000 222.350000 ;
      RECT 1183.500000 220.350000 1186.000000 223.650000 ;
      RECT 1169.500000 220.350000 1170.500000 221.650000 ;
      RECT 1169.500000 219.650000 1186.000000 220.350000 ;
      RECT 1169.500000 218.350000 1170.500000 219.650000 ;
      RECT 0.000000 218.350000 1156.500000 221.650000 ;
      RECT 0.000000 217.650000 1170.500000 218.350000 ;
      RECT 1183.500000 216.350000 1186.000000 219.650000 ;
      RECT 1169.500000 216.350000 1170.500000 217.650000 ;
      RECT 1169.500000 215.650000 1186.000000 216.350000 ;
      RECT 1169.500000 214.350000 1170.500000 215.650000 ;
      RECT 0.000000 214.350000 1156.500000 217.650000 ;
      RECT 0.000000 213.650000 1170.500000 214.350000 ;
      RECT 1183.500000 212.350000 1186.000000 215.650000 ;
      RECT 1169.500000 212.350000 1170.500000 213.650000 ;
      RECT 1169.500000 211.650000 1186.000000 212.350000 ;
      RECT 1169.500000 210.350000 1170.500000 211.650000 ;
      RECT 0.000000 210.350000 1156.500000 213.650000 ;
      RECT 0.000000 209.650000 1170.500000 210.350000 ;
      RECT 1183.500000 208.350000 1186.000000 211.650000 ;
      RECT 1169.500000 208.350000 1170.500000 209.650000 ;
      RECT 1169.500000 207.650000 1186.000000 208.350000 ;
      RECT 1169.500000 206.350000 1170.500000 207.650000 ;
      RECT 0.000000 206.350000 1156.500000 209.650000 ;
      RECT 0.000000 205.650000 1170.500000 206.350000 ;
      RECT 1183.500000 204.350000 1186.000000 207.650000 ;
      RECT 1169.500000 204.350000 1170.500000 205.650000 ;
      RECT 1169.500000 203.650000 1186.000000 204.350000 ;
      RECT 1169.500000 202.350000 1170.500000 203.650000 ;
      RECT 0.000000 202.350000 1156.500000 205.650000 ;
      RECT 0.000000 201.650000 1170.500000 202.350000 ;
      RECT 1183.500000 200.350000 1186.000000 203.650000 ;
      RECT 1169.500000 200.350000 1170.500000 201.650000 ;
      RECT 1169.500000 199.650000 1186.000000 200.350000 ;
      RECT 1169.500000 198.350000 1170.500000 199.650000 ;
      RECT 0.000000 198.350000 1156.500000 201.650000 ;
      RECT 0.000000 197.650000 1170.500000 198.350000 ;
      RECT 1183.500000 196.350000 1186.000000 199.650000 ;
      RECT 1169.500000 196.350000 1170.500000 197.650000 ;
      RECT 1169.500000 195.650000 1186.000000 196.350000 ;
      RECT 1169.500000 194.350000 1170.500000 195.650000 ;
      RECT 0.000000 194.350000 1156.500000 197.650000 ;
      RECT 0.000000 193.650000 1170.500000 194.350000 ;
      RECT 1183.500000 192.350000 1186.000000 195.650000 ;
      RECT 1169.500000 192.350000 1170.500000 193.650000 ;
      RECT 1169.500000 191.650000 1186.000000 192.350000 ;
      RECT 1169.500000 190.350000 1170.500000 191.650000 ;
      RECT 0.000000 190.350000 1156.500000 193.650000 ;
      RECT 0.000000 189.650000 1170.500000 190.350000 ;
      RECT 1183.500000 188.350000 1186.000000 191.650000 ;
      RECT 1169.500000 188.350000 1170.500000 189.650000 ;
      RECT 1169.500000 187.650000 1186.000000 188.350000 ;
      RECT 1169.500000 186.350000 1170.500000 187.650000 ;
      RECT 0.000000 186.350000 1156.500000 189.650000 ;
      RECT 0.000000 185.650000 1170.500000 186.350000 ;
      RECT 1183.500000 184.350000 1186.000000 187.650000 ;
      RECT 1169.500000 184.350000 1170.500000 185.650000 ;
      RECT 1169.500000 183.650000 1186.000000 184.350000 ;
      RECT 1169.500000 182.350000 1170.500000 183.650000 ;
      RECT 0.000000 182.350000 1156.500000 185.650000 ;
      RECT 0.000000 181.650000 1170.500000 182.350000 ;
      RECT 1183.500000 180.350000 1186.000000 183.650000 ;
      RECT 1169.500000 180.350000 1170.500000 181.650000 ;
      RECT 1169.500000 179.650000 1186.000000 180.350000 ;
      RECT 1169.500000 178.350000 1170.500000 179.650000 ;
      RECT 0.000000 178.350000 1156.500000 181.650000 ;
      RECT 0.000000 177.650000 1170.500000 178.350000 ;
      RECT 1183.500000 176.350000 1186.000000 179.650000 ;
      RECT 1169.500000 176.350000 1170.500000 177.650000 ;
      RECT 1169.500000 175.650000 1186.000000 176.350000 ;
      RECT 1169.500000 174.350000 1170.500000 175.650000 ;
      RECT 0.000000 174.350000 1156.500000 177.650000 ;
      RECT 0.000000 173.650000 1170.500000 174.350000 ;
      RECT 1183.500000 172.350000 1186.000000 175.650000 ;
      RECT 1169.500000 172.350000 1170.500000 173.650000 ;
      RECT 1169.500000 171.650000 1186.000000 172.350000 ;
      RECT 1169.500000 170.350000 1170.500000 171.650000 ;
      RECT 0.000000 170.350000 1156.500000 173.650000 ;
      RECT 0.000000 169.650000 1170.500000 170.350000 ;
      RECT 1183.500000 168.350000 1186.000000 171.650000 ;
      RECT 1169.500000 168.350000 1170.500000 169.650000 ;
      RECT 1169.500000 167.650000 1186.000000 168.350000 ;
      RECT 1169.500000 166.350000 1170.500000 167.650000 ;
      RECT 0.000000 166.350000 1156.500000 169.650000 ;
      RECT 0.000000 165.650000 1170.500000 166.350000 ;
      RECT 1183.500000 164.350000 1186.000000 167.650000 ;
      RECT 1169.500000 164.350000 1170.500000 165.650000 ;
      RECT 1169.500000 163.650000 1186.000000 164.350000 ;
      RECT 1169.500000 162.350000 1170.500000 163.650000 ;
      RECT 0.000000 162.350000 1156.500000 165.650000 ;
      RECT 0.000000 161.650000 1170.500000 162.350000 ;
      RECT 1183.500000 160.350000 1186.000000 163.650000 ;
      RECT 1169.500000 160.350000 1170.500000 161.650000 ;
      RECT 1169.500000 159.650000 1186.000000 160.350000 ;
      RECT 1169.500000 158.350000 1170.500000 159.650000 ;
      RECT 0.000000 158.350000 1156.500000 161.650000 ;
      RECT 0.000000 157.650000 1170.500000 158.350000 ;
      RECT 1183.500000 156.350000 1186.000000 159.650000 ;
      RECT 1169.500000 156.350000 1170.500000 157.650000 ;
      RECT 1169.500000 155.650000 1186.000000 156.350000 ;
      RECT 1169.500000 154.350000 1170.500000 155.650000 ;
      RECT 0.000000 154.350000 1156.500000 157.650000 ;
      RECT 0.000000 153.650000 1170.500000 154.350000 ;
      RECT 1183.500000 152.350000 1186.000000 155.650000 ;
      RECT 1169.500000 152.350000 1170.500000 153.650000 ;
      RECT 1169.500000 151.650000 1186.000000 152.350000 ;
      RECT 1169.500000 150.350000 1170.500000 151.650000 ;
      RECT 0.000000 150.350000 1156.500000 153.650000 ;
      RECT 0.000000 149.650000 1170.500000 150.350000 ;
      RECT 1183.500000 148.350000 1186.000000 151.650000 ;
      RECT 1169.500000 148.350000 1170.500000 149.650000 ;
      RECT 1169.500000 147.650000 1186.000000 148.350000 ;
      RECT 1169.500000 146.350000 1170.500000 147.650000 ;
      RECT 0.000000 146.350000 1156.500000 149.650000 ;
      RECT 0.000000 145.650000 1170.500000 146.350000 ;
      RECT 1183.500000 144.350000 1186.000000 147.650000 ;
      RECT 1169.500000 144.350000 1170.500000 145.650000 ;
      RECT 1169.500000 143.650000 1186.000000 144.350000 ;
      RECT 1169.500000 142.350000 1170.500000 143.650000 ;
      RECT 0.000000 142.350000 1156.500000 145.650000 ;
      RECT 0.000000 141.650000 1170.500000 142.350000 ;
      RECT 1183.500000 140.350000 1186.000000 143.650000 ;
      RECT 1169.500000 140.350000 1170.500000 141.650000 ;
      RECT 1169.500000 139.650000 1186.000000 140.350000 ;
      RECT 1169.500000 138.350000 1170.500000 139.650000 ;
      RECT 0.000000 138.350000 1156.500000 141.650000 ;
      RECT 0.000000 137.650000 1170.500000 138.350000 ;
      RECT 1183.500000 136.350000 1186.000000 139.650000 ;
      RECT 1169.500000 136.350000 1170.500000 137.650000 ;
      RECT 1169.500000 135.650000 1186.000000 136.350000 ;
      RECT 0.000000 135.650000 1156.500000 137.650000 ;
      RECT 1169.500000 134.350000 1170.500000 135.650000 ;
      RECT 1157.500000 133.650000 1170.500000 134.350000 ;
      RECT 1183.500000 132.350000 1186.000000 135.650000 ;
      RECT 1169.500000 132.350000 1170.500000 133.650000 ;
      RECT 0.000000 132.350000 1149.500000 135.650000 ;
      RECT 1169.500000 131.650000 1186.000000 132.350000 ;
      RECT 1169.500000 130.350000 1170.500000 131.650000 ;
      RECT 0.000000 130.350000 1156.500000 132.350000 ;
      RECT 0.000000 129.650000 1170.500000 130.350000 ;
      RECT 1183.500000 128.350000 1186.000000 131.650000 ;
      RECT 1169.500000 128.350000 1170.500000 129.650000 ;
      RECT 1169.500000 127.650000 1186.000000 128.350000 ;
      RECT 1169.500000 126.350000 1170.500000 127.650000 ;
      RECT 0.000000 126.350000 1156.500000 129.650000 ;
      RECT 0.000000 125.650000 1170.500000 126.350000 ;
      RECT 1183.500000 124.350000 1186.000000 127.650000 ;
      RECT 1169.500000 124.350000 1170.500000 125.650000 ;
      RECT 1169.500000 123.650000 1186.000000 124.350000 ;
      RECT 1169.500000 122.350000 1170.500000 123.650000 ;
      RECT 0.000000 122.350000 1156.500000 125.650000 ;
      RECT 0.000000 121.650000 1170.500000 122.350000 ;
      RECT 1183.500000 120.350000 1186.000000 123.650000 ;
      RECT 1169.500000 120.350000 1170.500000 121.650000 ;
      RECT 1169.500000 119.650000 1186.000000 120.350000 ;
      RECT 1169.500000 118.350000 1170.500000 119.650000 ;
      RECT 0.000000 118.350000 1156.500000 121.650000 ;
      RECT 0.000000 117.650000 1170.500000 118.350000 ;
      RECT 1183.500000 116.350000 1186.000000 119.650000 ;
      RECT 1169.500000 116.350000 1170.500000 117.650000 ;
      RECT 1169.500000 115.650000 1186.000000 116.350000 ;
      RECT 1169.500000 114.350000 1170.500000 115.650000 ;
      RECT 0.000000 114.350000 1156.500000 117.650000 ;
      RECT 0.000000 113.650000 1170.500000 114.350000 ;
      RECT 1183.500000 112.350000 1186.000000 115.650000 ;
      RECT 1169.500000 112.350000 1170.500000 113.650000 ;
      RECT 1169.500000 111.650000 1186.000000 112.350000 ;
      RECT 1169.500000 110.350000 1170.500000 111.650000 ;
      RECT 0.000000 110.350000 1156.500000 113.650000 ;
      RECT 0.000000 109.650000 1170.500000 110.350000 ;
      RECT 1183.500000 108.350000 1186.000000 111.650000 ;
      RECT 1169.500000 108.350000 1170.500000 109.650000 ;
      RECT 1169.500000 107.650000 1186.000000 108.350000 ;
      RECT 1169.500000 106.350000 1170.500000 107.650000 ;
      RECT 0.000000 106.350000 1156.500000 109.650000 ;
      RECT 0.000000 105.650000 1170.500000 106.350000 ;
      RECT 1183.500000 104.350000 1186.000000 107.650000 ;
      RECT 1169.500000 104.350000 1170.500000 105.650000 ;
      RECT 1169.500000 103.650000 1186.000000 104.350000 ;
      RECT 1169.500000 102.350000 1170.500000 103.650000 ;
      RECT 0.000000 102.350000 1156.500000 105.650000 ;
      RECT 0.000000 101.650000 1170.500000 102.350000 ;
      RECT 1183.500000 100.350000 1186.000000 103.650000 ;
      RECT 1169.500000 100.350000 1170.500000 101.650000 ;
      RECT 1169.500000 99.650000 1186.000000 100.350000 ;
      RECT 1169.500000 98.350000 1170.500000 99.650000 ;
      RECT 0.000000 98.350000 1156.500000 101.650000 ;
      RECT 0.000000 97.650000 1170.500000 98.350000 ;
      RECT 1183.500000 96.350000 1186.000000 99.650000 ;
      RECT 1169.500000 96.350000 1170.500000 97.650000 ;
      RECT 1169.500000 95.650000 1186.000000 96.350000 ;
      RECT 1169.500000 94.350000 1170.500000 95.650000 ;
      RECT 0.000000 94.350000 1156.500000 97.650000 ;
      RECT 0.000000 93.650000 1170.500000 94.350000 ;
      RECT 1183.500000 92.350000 1186.000000 95.650000 ;
      RECT 1169.500000 92.350000 1170.500000 93.650000 ;
      RECT 1169.500000 91.650000 1186.000000 92.350000 ;
      RECT 1169.500000 90.350000 1170.500000 91.650000 ;
      RECT 0.000000 90.350000 1156.500000 93.650000 ;
      RECT 0.000000 89.650000 1170.500000 90.350000 ;
      RECT 1183.500000 88.350000 1186.000000 91.650000 ;
      RECT 1169.500000 88.350000 1170.500000 89.650000 ;
      RECT 1169.500000 87.650000 1186.000000 88.350000 ;
      RECT 1169.500000 86.350000 1170.500000 87.650000 ;
      RECT 0.000000 86.350000 1156.500000 89.650000 ;
      RECT 0.000000 85.650000 1170.500000 86.350000 ;
      RECT 1183.500000 84.350000 1186.000000 87.650000 ;
      RECT 1169.500000 84.350000 1170.500000 85.650000 ;
      RECT 1169.500000 83.650000 1186.000000 84.350000 ;
      RECT 1169.500000 82.350000 1170.500000 83.650000 ;
      RECT 0.000000 82.350000 1156.500000 85.650000 ;
      RECT 0.000000 81.650000 1170.500000 82.350000 ;
      RECT 1183.500000 80.350000 1186.000000 83.650000 ;
      RECT 1169.500000 80.350000 1170.500000 81.650000 ;
      RECT 1169.500000 79.650000 1186.000000 80.350000 ;
      RECT 1169.500000 78.350000 1170.500000 79.650000 ;
      RECT 0.000000 78.350000 1156.500000 81.650000 ;
      RECT 0.000000 77.650000 1170.500000 78.350000 ;
      RECT 1183.500000 76.350000 1186.000000 79.650000 ;
      RECT 1169.500000 76.350000 1170.500000 77.650000 ;
      RECT 1169.500000 75.650000 1186.000000 76.350000 ;
      RECT 1169.500000 74.350000 1170.500000 75.650000 ;
      RECT 0.000000 74.350000 1156.500000 77.650000 ;
      RECT 0.000000 73.650000 1170.500000 74.350000 ;
      RECT 1183.500000 72.350000 1186.000000 75.650000 ;
      RECT 1169.500000 72.350000 1170.500000 73.650000 ;
      RECT 1169.500000 71.650000 1186.000000 72.350000 ;
      RECT 1169.500000 70.350000 1170.500000 71.650000 ;
      RECT 0.000000 70.350000 1156.500000 73.650000 ;
      RECT 0.000000 69.650000 1170.500000 70.350000 ;
      RECT 1183.500000 68.350000 1186.000000 71.650000 ;
      RECT 1169.500000 68.350000 1170.500000 69.650000 ;
      RECT 1169.500000 67.650000 1186.000000 68.350000 ;
      RECT 1169.500000 66.350000 1170.500000 67.650000 ;
      RECT 0.000000 66.350000 1156.500000 69.650000 ;
      RECT 0.000000 65.650000 1170.500000 66.350000 ;
      RECT 1183.500000 64.350000 1186.000000 67.650000 ;
      RECT 1169.500000 64.350000 1170.500000 65.650000 ;
      RECT 1169.500000 63.650000 1186.000000 64.350000 ;
      RECT 1169.500000 62.350000 1170.500000 63.650000 ;
      RECT 0.000000 62.350000 1156.500000 65.650000 ;
      RECT 0.000000 61.650000 1170.500000 62.350000 ;
      RECT 1183.500000 60.350000 1186.000000 63.650000 ;
      RECT 1169.500000 60.350000 1170.500000 61.650000 ;
      RECT 1169.500000 59.650000 1186.000000 60.350000 ;
      RECT 1169.500000 58.350000 1170.500000 59.650000 ;
      RECT 0.000000 58.350000 1156.500000 61.650000 ;
      RECT 0.000000 57.650000 1170.500000 58.350000 ;
      RECT 1183.500000 56.350000 1186.000000 59.650000 ;
      RECT 1169.500000 56.350000 1170.500000 57.650000 ;
      RECT 1169.500000 55.650000 1186.000000 56.350000 ;
      RECT 1169.500000 54.350000 1170.500000 55.650000 ;
      RECT 0.000000 54.350000 1156.500000 57.650000 ;
      RECT 0.000000 53.650000 1170.500000 54.350000 ;
      RECT 1183.500000 52.350000 1186.000000 55.650000 ;
      RECT 1169.500000 52.350000 1170.500000 53.650000 ;
      RECT 1169.500000 51.650000 1186.000000 52.350000 ;
      RECT 1169.500000 50.350000 1170.500000 51.650000 ;
      RECT 0.000000 50.350000 1156.500000 53.650000 ;
      RECT 0.000000 49.650000 1170.500000 50.350000 ;
      RECT 1183.500000 48.350000 1186.000000 51.650000 ;
      RECT 1169.500000 48.350000 1170.500000 49.650000 ;
      RECT 1169.500000 47.650000 1186.000000 48.350000 ;
      RECT 1169.500000 46.350000 1170.500000 47.650000 ;
      RECT 0.000000 46.350000 1156.500000 49.650000 ;
      RECT 0.000000 45.650000 1170.500000 46.350000 ;
      RECT 1183.500000 44.350000 1186.000000 47.650000 ;
      RECT 1169.500000 44.350000 1170.500000 45.650000 ;
      RECT 1169.500000 43.650000 1186.000000 44.350000 ;
      RECT 1169.500000 42.350000 1170.500000 43.650000 ;
      RECT 0.000000 42.350000 1156.500000 45.650000 ;
      RECT 0.000000 41.650000 1170.500000 42.350000 ;
      RECT 1183.500000 40.350000 1186.000000 43.650000 ;
      RECT 1169.500000 40.350000 1170.500000 41.650000 ;
      RECT 1169.500000 39.650000 1186.000000 40.350000 ;
      RECT 1169.500000 38.350000 1170.500000 39.650000 ;
      RECT 0.000000 38.350000 1156.500000 41.650000 ;
      RECT 0.000000 37.650000 1170.500000 38.350000 ;
      RECT 1183.500000 36.350000 1186.000000 39.650000 ;
      RECT 1169.500000 36.350000 1170.500000 37.650000 ;
      RECT 1169.500000 35.650000 1186.000000 36.350000 ;
      RECT 1169.500000 34.350000 1170.500000 35.650000 ;
      RECT 0.000000 34.350000 1156.500000 37.650000 ;
      RECT 0.000000 33.650000 1170.500000 34.350000 ;
      RECT 1183.500000 32.350000 1186.000000 35.650000 ;
      RECT 1169.500000 32.350000 1170.500000 33.650000 ;
      RECT 1169.500000 31.650000 1186.000000 32.350000 ;
      RECT 1169.500000 30.350000 1170.500000 31.650000 ;
      RECT 0.000000 30.350000 1156.500000 33.650000 ;
      RECT 0.000000 29.650000 1170.500000 30.350000 ;
      RECT 1183.500000 28.350000 1186.000000 31.650000 ;
      RECT 1169.500000 28.350000 1170.500000 29.650000 ;
      RECT 1169.500000 27.650000 1186.000000 28.350000 ;
      RECT 1169.500000 26.350000 1170.500000 27.650000 ;
      RECT 0.000000 26.350000 1156.500000 29.650000 ;
      RECT 0.000000 25.650000 1170.500000 26.350000 ;
      RECT 1183.500000 24.350000 1186.000000 27.650000 ;
      RECT 1169.500000 24.350000 1170.500000 25.650000 ;
      RECT 1169.500000 23.650000 1186.000000 24.350000 ;
      RECT 1169.500000 22.350000 1170.500000 23.650000 ;
      RECT 0.000000 22.350000 1156.500000 25.650000 ;
      RECT 0.000000 21.650000 1170.500000 22.350000 ;
      RECT 1183.500000 20.350000 1186.000000 23.650000 ;
      RECT 1169.500000 20.350000 1170.500000 21.650000 ;
      RECT 1169.500000 19.650000 1186.000000 20.350000 ;
      RECT 1169.500000 18.350000 1170.500000 19.650000 ;
      RECT 0.000000 18.350000 1156.500000 21.650000 ;
      RECT 0.000000 17.650000 1170.500000 18.350000 ;
      RECT 1183.500000 16.350000 1186.000000 19.650000 ;
      RECT 1166.500000 16.350000 1170.500000 17.650000 ;
      RECT 1166.500000 15.650000 1186.000000 16.350000 ;
      RECT 1166.500000 14.350000 1170.500000 15.650000 ;
      RECT 0.000000 14.350000 1158.500000 17.650000 ;
      RECT 0.000000 13.650000 1170.500000 14.350000 ;
      RECT 1183.500000 12.350000 1186.000000 15.650000 ;
      RECT 1166.500000 12.350000 1170.500000 13.650000 ;
      RECT 1166.500000 11.650000 1186.000000 12.350000 ;
      RECT 1166.500000 10.350000 1170.500000 11.650000 ;
      RECT 0.000000 10.350000 1158.500000 13.650000 ;
      RECT 0.000000 9.650000 1170.500000 10.350000 ;
      RECT 1183.500000 8.350000 1186.000000 11.650000 ;
      RECT 1166.500000 8.350000 1170.500000 9.650000 ;
      RECT 1166.500000 7.650000 1186.000000 8.350000 ;
      RECT 1116.500000 7.650000 1158.500000 9.650000 ;
      RECT 1066.500000 7.650000 1108.500000 9.650000 ;
      RECT 1016.500000 7.650000 1058.500000 9.650000 ;
      RECT 966.500000 7.650000 1008.500000 9.650000 ;
      RECT 916.500000 7.650000 958.500000 9.650000 ;
      RECT 866.500000 7.650000 908.500000 9.650000 ;
      RECT 816.500000 7.650000 858.500000 9.650000 ;
      RECT 766.500000 7.650000 808.500000 9.650000 ;
      RECT 716.500000 7.650000 758.500000 9.650000 ;
      RECT 666.500000 7.650000 708.500000 9.650000 ;
      RECT 616.500000 7.650000 658.500000 9.650000 ;
      RECT 566.500000 7.650000 608.500000 9.650000 ;
      RECT 516.500000 7.650000 558.500000 9.650000 ;
      RECT 466.500000 7.650000 508.500000 9.650000 ;
      RECT 416.500000 7.650000 458.500000 9.650000 ;
      RECT 366.500000 7.650000 408.500000 9.650000 ;
      RECT 316.500000 7.650000 358.500000 9.650000 ;
      RECT 266.500000 7.650000 308.500000 9.650000 ;
      RECT 216.500000 7.650000 258.500000 9.650000 ;
      RECT 166.500000 7.650000 208.500000 9.650000 ;
      RECT 116.500000 7.650000 158.500000 9.650000 ;
      RECT 66.500000 7.650000 108.500000 9.650000 ;
      RECT 0.000000 7.650000 58.500000 9.650000 ;
      RECT 1166.500000 6.350000 1170.500000 7.650000 ;
      RECT 1157.500000 6.350000 1158.500000 7.650000 ;
      RECT 1116.500000 6.350000 1149.500000 7.650000 ;
      RECT 1107.500000 6.350000 1108.500000 7.650000 ;
      RECT 1066.500000 6.350000 1099.500000 7.650000 ;
      RECT 1057.500000 6.350000 1058.500000 7.650000 ;
      RECT 1016.500000 6.350000 1049.500000 7.650000 ;
      RECT 1007.500000 6.350000 1008.500000 7.650000 ;
      RECT 966.500000 6.350000 999.500000 7.650000 ;
      RECT 957.500000 6.350000 958.500000 7.650000 ;
      RECT 916.500000 6.350000 949.500000 7.650000 ;
      RECT 907.500000 6.350000 908.500000 7.650000 ;
      RECT 866.500000 6.350000 899.500000 7.650000 ;
      RECT 857.500000 6.350000 858.500000 7.650000 ;
      RECT 816.500000 6.350000 849.500000 7.650000 ;
      RECT 807.500000 6.350000 808.500000 7.650000 ;
      RECT 766.500000 6.350000 799.500000 7.650000 ;
      RECT 757.500000 6.350000 758.500000 7.650000 ;
      RECT 716.500000 6.350000 749.500000 7.650000 ;
      RECT 707.500000 6.350000 708.500000 7.650000 ;
      RECT 666.500000 6.350000 699.500000 7.650000 ;
      RECT 657.500000 6.350000 658.500000 7.650000 ;
      RECT 616.500000 6.350000 649.500000 7.650000 ;
      RECT 607.500000 6.350000 608.500000 7.650000 ;
      RECT 566.500000 6.350000 599.500000 7.650000 ;
      RECT 557.500000 6.350000 558.500000 7.650000 ;
      RECT 516.500000 6.350000 549.500000 7.650000 ;
      RECT 507.500000 6.350000 508.500000 7.650000 ;
      RECT 466.500000 6.350000 499.500000 7.650000 ;
      RECT 457.500000 6.350000 458.500000 7.650000 ;
      RECT 416.500000 6.350000 449.500000 7.650000 ;
      RECT 407.500000 6.350000 408.500000 7.650000 ;
      RECT 366.500000 6.350000 399.500000 7.650000 ;
      RECT 357.500000 6.350000 358.500000 7.650000 ;
      RECT 316.500000 6.350000 349.500000 7.650000 ;
      RECT 307.500000 6.350000 308.500000 7.650000 ;
      RECT 266.500000 6.350000 299.500000 7.650000 ;
      RECT 257.500000 6.350000 258.500000 7.650000 ;
      RECT 216.500000 6.350000 249.500000 7.650000 ;
      RECT 207.500000 6.350000 208.500000 7.650000 ;
      RECT 166.500000 6.350000 199.500000 7.650000 ;
      RECT 157.500000 6.350000 158.500000 7.650000 ;
      RECT 116.500000 6.350000 149.500000 7.650000 ;
      RECT 107.500000 6.350000 108.500000 7.650000 ;
      RECT 66.500000 6.350000 99.500000 7.650000 ;
      RECT 57.500000 6.350000 58.500000 7.650000 ;
      RECT 1157.500000 5.650000 1170.500000 6.350000 ;
      RECT 1107.500000 5.650000 1149.500000 6.350000 ;
      RECT 1057.500000 5.650000 1099.500000 6.350000 ;
      RECT 1007.500000 5.650000 1049.500000 6.350000 ;
      RECT 957.500000 5.650000 999.500000 6.350000 ;
      RECT 907.500000 5.650000 949.500000 6.350000 ;
      RECT 857.500000 5.650000 899.500000 6.350000 ;
      RECT 807.500000 5.650000 849.500000 6.350000 ;
      RECT 757.500000 5.650000 799.500000 6.350000 ;
      RECT 707.500000 5.650000 749.500000 6.350000 ;
      RECT 657.500000 5.650000 699.500000 6.350000 ;
      RECT 607.500000 5.650000 649.500000 6.350000 ;
      RECT 557.500000 5.650000 599.500000 6.350000 ;
      RECT 507.500000 5.650000 549.500000 6.350000 ;
      RECT 457.500000 5.650000 499.500000 6.350000 ;
      RECT 407.500000 5.650000 449.500000 6.350000 ;
      RECT 357.500000 5.650000 399.500000 6.350000 ;
      RECT 307.500000 5.650000 349.500000 6.350000 ;
      RECT 257.500000 5.650000 299.500000 6.350000 ;
      RECT 207.500000 5.650000 249.500000 6.350000 ;
      RECT 157.500000 5.650000 199.500000 6.350000 ;
      RECT 107.500000 5.650000 149.500000 6.350000 ;
      RECT 57.500000 5.650000 99.500000 6.350000 ;
      RECT 1183.500000 4.350000 1186.000000 7.650000 ;
      RECT 1166.500000 4.350000 1170.500000 5.650000 ;
      RECT 1157.500000 4.350000 1158.500000 5.650000 ;
      RECT 1116.500000 4.350000 1149.500000 5.650000 ;
      RECT 1107.500000 4.350000 1108.500000 5.650000 ;
      RECT 1066.500000 4.350000 1099.500000 5.650000 ;
      RECT 1057.500000 4.350000 1058.500000 5.650000 ;
      RECT 1016.500000 4.350000 1049.500000 5.650000 ;
      RECT 1007.500000 4.350000 1008.500000 5.650000 ;
      RECT 966.500000 4.350000 999.500000 5.650000 ;
      RECT 957.500000 4.350000 958.500000 5.650000 ;
      RECT 916.500000 4.350000 949.500000 5.650000 ;
      RECT 907.500000 4.350000 908.500000 5.650000 ;
      RECT 866.500000 4.350000 899.500000 5.650000 ;
      RECT 857.500000 4.350000 858.500000 5.650000 ;
      RECT 816.500000 4.350000 849.500000 5.650000 ;
      RECT 807.500000 4.350000 808.500000 5.650000 ;
      RECT 766.500000 4.350000 799.500000 5.650000 ;
      RECT 757.500000 4.350000 758.500000 5.650000 ;
      RECT 716.500000 4.350000 749.500000 5.650000 ;
      RECT 707.500000 4.350000 708.500000 5.650000 ;
      RECT 666.500000 4.350000 699.500000 5.650000 ;
      RECT 657.500000 4.350000 658.500000 5.650000 ;
      RECT 616.500000 4.350000 649.500000 5.650000 ;
      RECT 607.500000 4.350000 608.500000 5.650000 ;
      RECT 566.500000 4.350000 599.500000 5.650000 ;
      RECT 557.500000 4.350000 558.500000 5.650000 ;
      RECT 516.500000 4.350000 549.500000 5.650000 ;
      RECT 507.500000 4.350000 508.500000 5.650000 ;
      RECT 466.500000 4.350000 499.500000 5.650000 ;
      RECT 457.500000 4.350000 458.500000 5.650000 ;
      RECT 416.500000 4.350000 449.500000 5.650000 ;
      RECT 407.500000 4.350000 408.500000 5.650000 ;
      RECT 366.500000 4.350000 399.500000 5.650000 ;
      RECT 357.500000 4.350000 358.500000 5.650000 ;
      RECT 316.500000 4.350000 349.500000 5.650000 ;
      RECT 307.500000 4.350000 308.500000 5.650000 ;
      RECT 266.500000 4.350000 299.500000 5.650000 ;
      RECT 257.500000 4.350000 258.500000 5.650000 ;
      RECT 216.500000 4.350000 249.500000 5.650000 ;
      RECT 207.500000 4.350000 208.500000 5.650000 ;
      RECT 166.500000 4.350000 199.500000 5.650000 ;
      RECT 157.500000 4.350000 158.500000 5.650000 ;
      RECT 116.500000 4.350000 149.500000 5.650000 ;
      RECT 107.500000 4.350000 108.500000 5.650000 ;
      RECT 66.500000 4.350000 99.500000 5.650000 ;
      RECT 57.500000 4.350000 58.500000 5.650000 ;
      RECT 15.500000 4.350000 49.500000 7.650000 ;
      RECT 0.000000 4.350000 2.500000 7.650000 ;
      RECT 1116.500000 3.650000 1158.500000 4.350000 ;
      RECT 1066.500000 3.650000 1108.500000 4.350000 ;
      RECT 1016.500000 3.650000 1058.500000 4.350000 ;
      RECT 966.500000 3.650000 1008.500000 4.350000 ;
      RECT 916.500000 3.650000 958.500000 4.350000 ;
      RECT 866.500000 3.650000 908.500000 4.350000 ;
      RECT 816.500000 3.650000 858.500000 4.350000 ;
      RECT 766.500000 3.650000 808.500000 4.350000 ;
      RECT 716.500000 3.650000 758.500000 4.350000 ;
      RECT 666.500000 3.650000 708.500000 4.350000 ;
      RECT 616.500000 3.650000 658.500000 4.350000 ;
      RECT 566.500000 3.650000 608.500000 4.350000 ;
      RECT 516.500000 3.650000 558.500000 4.350000 ;
      RECT 466.500000 3.650000 508.500000 4.350000 ;
      RECT 416.500000 3.650000 458.500000 4.350000 ;
      RECT 366.500000 3.650000 408.500000 4.350000 ;
      RECT 316.500000 3.650000 358.500000 4.350000 ;
      RECT 266.500000 3.650000 308.500000 4.350000 ;
      RECT 216.500000 3.650000 258.500000 4.350000 ;
      RECT 166.500000 3.650000 208.500000 4.350000 ;
      RECT 116.500000 3.650000 158.500000 4.350000 ;
      RECT 66.500000 3.650000 108.500000 4.350000 ;
      RECT 0.000000 3.650000 58.500000 4.350000 ;
      RECT 1166.500000 2.350000 1186.000000 4.350000 ;
      RECT 1157.500000 2.350000 1158.500000 3.650000 ;
      RECT 1116.500000 2.350000 1149.500000 3.650000 ;
      RECT 1107.500000 2.350000 1108.500000 3.650000 ;
      RECT 1066.500000 2.350000 1099.500000 3.650000 ;
      RECT 1057.500000 2.350000 1058.500000 3.650000 ;
      RECT 1016.500000 2.350000 1049.500000 3.650000 ;
      RECT 1007.500000 2.350000 1008.500000 3.650000 ;
      RECT 966.500000 2.350000 999.500000 3.650000 ;
      RECT 957.500000 2.350000 958.500000 3.650000 ;
      RECT 916.500000 2.350000 949.500000 3.650000 ;
      RECT 907.500000 2.350000 908.500000 3.650000 ;
      RECT 866.500000 2.350000 899.500000 3.650000 ;
      RECT 857.500000 2.350000 858.500000 3.650000 ;
      RECT 816.500000 2.350000 849.500000 3.650000 ;
      RECT 807.500000 2.350000 808.500000 3.650000 ;
      RECT 766.500000 2.350000 799.500000 3.650000 ;
      RECT 757.500000 2.350000 758.500000 3.650000 ;
      RECT 716.500000 2.350000 749.500000 3.650000 ;
      RECT 707.500000 2.350000 708.500000 3.650000 ;
      RECT 666.500000 2.350000 699.500000 3.650000 ;
      RECT 657.500000 2.350000 658.500000 3.650000 ;
      RECT 616.500000 2.350000 649.500000 3.650000 ;
      RECT 607.500000 2.350000 608.500000 3.650000 ;
      RECT 566.500000 2.350000 599.500000 3.650000 ;
      RECT 557.500000 2.350000 558.500000 3.650000 ;
      RECT 516.500000 2.350000 549.500000 3.650000 ;
      RECT 507.500000 2.350000 508.500000 3.650000 ;
      RECT 466.500000 2.350000 499.500000 3.650000 ;
      RECT 457.500000 2.350000 458.500000 3.650000 ;
      RECT 416.500000 2.350000 449.500000 3.650000 ;
      RECT 407.500000 2.350000 408.500000 3.650000 ;
      RECT 366.500000 2.350000 399.500000 3.650000 ;
      RECT 357.500000 2.350000 358.500000 3.650000 ;
      RECT 316.500000 2.350000 349.500000 3.650000 ;
      RECT 307.500000 2.350000 308.500000 3.650000 ;
      RECT 266.500000 2.350000 299.500000 3.650000 ;
      RECT 257.500000 2.350000 258.500000 3.650000 ;
      RECT 216.500000 2.350000 249.500000 3.650000 ;
      RECT 207.500000 2.350000 208.500000 3.650000 ;
      RECT 166.500000 2.350000 199.500000 3.650000 ;
      RECT 157.500000 2.350000 158.500000 3.650000 ;
      RECT 116.500000 2.350000 149.500000 3.650000 ;
      RECT 107.500000 2.350000 108.500000 3.650000 ;
      RECT 66.500000 2.350000 99.500000 3.650000 ;
      RECT 57.500000 2.350000 58.500000 3.650000 ;
      RECT 1157.500000 0.350000 1186.000000 2.350000 ;
      RECT 1107.500000 0.350000 1149.500000 2.350000 ;
      RECT 1057.500000 0.350000 1099.500000 2.350000 ;
      RECT 1007.500000 0.350000 1049.500000 2.350000 ;
      RECT 957.500000 0.350000 999.500000 2.350000 ;
      RECT 907.500000 0.350000 949.500000 2.350000 ;
      RECT 857.500000 0.350000 899.500000 2.350000 ;
      RECT 807.500000 0.350000 849.500000 2.350000 ;
      RECT 757.500000 0.350000 799.500000 2.350000 ;
      RECT 707.500000 0.350000 749.500000 2.350000 ;
      RECT 657.500000 0.350000 699.500000 2.350000 ;
      RECT 607.500000 0.350000 649.500000 2.350000 ;
      RECT 557.500000 0.350000 599.500000 2.350000 ;
      RECT 507.500000 0.350000 549.500000 2.350000 ;
      RECT 457.500000 0.350000 499.500000 2.350000 ;
      RECT 407.500000 0.350000 449.500000 2.350000 ;
      RECT 357.500000 0.350000 399.500000 2.350000 ;
      RECT 307.500000 0.350000 349.500000 2.350000 ;
      RECT 257.500000 0.350000 299.500000 2.350000 ;
      RECT 207.500000 0.350000 249.500000 2.350000 ;
      RECT 157.500000 0.350000 199.500000 2.350000 ;
      RECT 107.500000 0.350000 149.500000 2.350000 ;
      RECT 57.500000 0.350000 99.500000 2.350000 ;
      RECT 0.000000 0.350000 49.500000 3.650000 ;
      RECT 0.000000 0.000000 1186.000000 0.350000 ;
  END
END MCU

END LIBRARY
