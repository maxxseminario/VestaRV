##
## LEF for PtnCells ;
## created by Innovus v20.12-s088_1 on Sat Nov 22 14:45:59 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO MCU
  CLASS BLOCK ;
  SIZE 1186.000000 BY 686.000000 ;
  FOREIGN MCU 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN resetn_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9625 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.235 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.658 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9392 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 24.822 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 109.261 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6  ;
    ANTENNAMAXAREACAR 947.445 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 4175.42 LAYER M6  ;
    ANTENNAMAXCUTCAR 3.32103 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 131.365000 0.000000 131.465000 0.520000 ;
    END
  END resetn_in
  PIN resetn_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.301 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3684 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 111.130000 0.000000 111.230000 0.520000 ;
    END
  END resetn_out
  PIN resetn_dir
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.3585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6654 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 121.725000 0.000000 121.825000 0.520000 ;
    END
  END resetn_dir
  PIN resetn_ren
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.7635 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4474 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 125.685000 0.000000 125.785000 0.520000 ;
    END
  END resetn_ren
  PIN prt1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.7525 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.711 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 5.302 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3728 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0447 LAYER M3  ;
    ANTENNAMAXAREACAR 138.548 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 604.264 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.894855 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 45.565000 1186.000000 45.665000 ;
    END
  END prt1_in[7]
  PIN prt1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.5745 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.3718 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 6.958 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.6592 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M3  ;
    ANTENNAMAXAREACAR 38.0959 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 167.594 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.209644 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 133.565000 1186.000000 133.665000 ;
    END
  END prt1_in[6]
  PIN prt1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7925 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.887 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 14.322 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.0608 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M3  ;
    ANTENNAMAXAREACAR 115.252 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 503.994 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.314465 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 221.565000 1186.000000 221.665000 ;
    END
  END prt1_in[5]
  PIN prt1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6125 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.695 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 14.402 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.4128 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 6.982 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 30.7648 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M5  ;
    ANTENNAMAXAREACAR 62.1745 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 274.23 LAYER M5  ;
    ANTENNAMAXCUTCAR 0.628931 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 309.565000 1186.000000 309.665000 ;
    END
  END prt1_in[4]
  PIN prt1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.282 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5862 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 7.76 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.712 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 LAYER M4  ;
    ANTENNAMAXAREACAR 47.6053 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 62.8176 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.786164 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 397.565000 1186.000000 397.665000 ;
    END
  END prt1_in[3]
  PIN prt1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0935 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.0554 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 9.322 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.0608 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 13.902 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 61.2128 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M5  ;
    ANTENNAMAXAREACAR 395.441 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 1741.66 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.01511 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 485.565000 1186.000000 485.665000 ;
    END
  END prt1_in[2]
  PIN prt1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0135 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.3034 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 8.802 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.7728 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0671 LAYER M3  ;
    ANTENNAMAXAREACAR 154.676 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 673.103 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.596125 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 573.565000 1186.000000 573.665000 ;
    END
  END prt1_in[1]
  PIN prt1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.1195 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 97.3258 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 7.058 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.0992 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0595 LAYER M3  ;
    ANTENNAMAXAREACAR 129.861 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 568.531 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.672269 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 661.565000 1186.000000 661.665000 ;
    END
  END prt1_in[0]
  PIN prt1_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.496 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.7824 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 25.330000 1186.000000 25.430000 ;
    END
  END prt1_out[7]
  PIN prt1_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.426 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7184 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 113.330000 1186.000000 113.430000 ;
    END
  END prt1_out[6]
  PIN prt1_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 11.643 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.3172 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 201.330000 1186.000000 201.430000 ;
    END
  END prt1_out[5]
  PIN prt1_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 289.330000 1186.000000 289.430000 ;
    END
  END prt1_out[4]
  PIN prt1_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.41 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.848 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 377.330000 1186.000000 377.430000 ;
    END
  END prt1_out[3]
  PIN prt1_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 465.330000 1186.000000 465.430000 ;
    END
  END prt1_out[2]
  PIN prt1_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 553.330000 1186.000000 553.430000 ;
    END
  END prt1_out[1]
  PIN prt1_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 6.45 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.424 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 641.330000 1186.000000 641.430000 ;
    END
  END prt1_out[0]
  PIN prt1_dir[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 35.925000 1186.000000 36.025000 ;
    END
  END prt1_dir[7]
  PIN prt1_dir[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.446 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8064 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 123.925000 1186.000000 124.025000 ;
    END
  END prt1_dir[6]
  PIN prt1_dir[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 211.925000 1186.000000 212.025000 ;
    END
  END prt1_dir[5]
  PIN prt1_dir[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 299.925000 1186.000000 300.025000 ;
    END
  END prt1_dir[4]
  PIN prt1_dir[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 387.925000 1186.000000 388.025000 ;
    END
  END prt1_dir[3]
  PIN prt1_dir[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 475.925000 1186.000000 476.025000 ;
    END
  END prt1_dir[2]
  PIN prt1_dir[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 12.9945 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.2638 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 563.925000 1186.000000 564.025000 ;
    END
  END prt1_dir[1]
  PIN prt1_dir[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 5.1535 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.7194 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 651.925000 1186.000000 652.025000 ;
    END
  END prt1_dir[0]
  PIN prt1_ren[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 39.885000 1186.000000 39.985000 ;
    END
  END prt1_ren[7]
  PIN prt1_ren[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5302 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.326 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4784 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 127.885000 1186.000000 127.985000 ;
    END
  END prt1_ren[6]
  PIN prt1_ren[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0805 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3542 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.326 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2784 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 215.885000 1186.000000 215.985000 ;
    END
  END prt1_ren[5]
  PIN prt1_ren[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 303.885000 1186.000000 303.985000 ;
    END
  END prt1_ren[4]
  PIN prt1_ren[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9075 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.993 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 4.242 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7088 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 391.885000 1186.000000 391.985000 ;
    END
  END prt1_ren[3]
  PIN prt1_ren[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5455 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 3.708 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4032 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 479.885000 1186.000000 479.985000 ;
    END
  END prt1_ren[2]
  PIN prt1_ren[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 567.885000 1186.000000 567.985000 ;
    END
  END prt1_ren[1]
  PIN prt1_ren[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 655.885000 1186.000000 655.985000 ;
    END
  END prt1_ren[0]
  PIN prt2_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5545 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4838 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2214 LAYER M2  ;
    ANTENNAMAXAREACAR 2.82385 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 12.2674 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.0903342 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 302.965000 0.000000 303.065000 0.520000 ;
    END
  END prt2_in[7]
  PIN prt2_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3175 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.441 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2  ;
    ANTENNAMAXAREACAR 7.41509 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 30.5173 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 388.765000 0.000000 388.865000 0.520000 ;
    END
  END prt2_in[6]
  PIN prt2_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4125 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.815 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3408 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3  ;
    ANTENNAMAXAREACAR 36.2639 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 159.377 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 474.565000 0.000000 474.665000 0.520000 ;
    END
  END prt2_in[5]
  PIN prt2_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3175 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.441 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2  ;
    ANTENNAMAXAREACAR 29.6974 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 122.813 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 560.365000 0.000000 560.465000 0.520000 ;
    END
  END prt2_in[4]
  PIN prt2_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.344 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4378 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 2.564 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9964 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 2.64 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.08 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6996 LAYER M4  ;
    ANTENNAMAXAREACAR 4.58433 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 6.73871 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.0857633 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 646.165000 0.000000 646.265000 0.520000 ;
    END
  END prt2_in[3]
  PIN prt2_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3125 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.375 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2  ;
    ANTENNAMAXAREACAR 3.41352 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 14.1494 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 731.965000 0.000000 732.065000 0.520000 ;
    END
  END prt2_in[2]
  PIN prt2_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.691 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 15.998 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.4352 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 LAYER M3  ;
    ANTENNAMAXAREACAR 156.76 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 683.874 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.37037 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 817.765000 0.000000 817.865000 0.520000 ;
    END
  END prt2_in[1]
  PIN prt2_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1755 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7722 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 29.522 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.941 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3  ;
    ANTENNAMAXAREACAR 336.377 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1479.88 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 903.565000 0.000000 903.665000 0.520000 ;
    END
  END prt2_in[0]
  PIN prt2_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.701 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1284 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 282.730000 0.000000 282.830000 0.520000 ;
    END
  END prt2_out[7]
  PIN prt2_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.691 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 5.422 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.9008 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 368.530000 0.000000 368.630000 0.520000 ;
    END
  END prt2_out[6]
  PIN prt2_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 11.138 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.0512 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 454.330000 0.000000 454.430000 0.520000 ;
    END
  END prt2_out[5]
  PIN prt2_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.721 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 540.130000 0.000000 540.230000 0.520000 ;
    END
  END prt2_out[4]
  PIN prt2_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.717 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1988 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 625.930000 0.000000 626.030000 0.520000 ;
    END
  END prt2_out[3]
  PIN prt2_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.759 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4276 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 711.730000 0.000000 711.830000 0.520000 ;
    END
  END prt2_out[2]
  PIN prt2_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.649 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8996 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 797.530000 0.000000 797.630000 0.520000 ;
    END
  END prt2_out[1]
  PIN prt2_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.512 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 883.330000 0.000000 883.430000 0.520000 ;
    END
  END prt2_out[0]
  PIN prt2_dir[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3165 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3926 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.306 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.9904 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 293.325000 0.000000 293.425000 0.520000 ;
    END
  END prt2_dir[7]
  PIN prt2_dir[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5165 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2726 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 8.102 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.6928 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 379.125000 0.000000 379.225000 0.520000 ;
    END
  END prt2_dir[6]
  PIN prt2_dir[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.7195 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2538 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 464.925000 0.000000 465.025000 0.520000 ;
    END
  END prt2_dir[5]
  PIN prt2_dir[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.411 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8084 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.922 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5008 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 550.725000 0.000000 550.825000 0.520000 ;
    END
  END prt2_dir[4]
  PIN prt2_dir[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.6965 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1086 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 636.525000 0.000000 636.625000 0.520000 ;
    END
  END prt2_dir[3]
  PIN prt2_dir[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.3115 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3706 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 722.325000 0.000000 722.425000 0.520000 ;
    END
  END prt2_dir[2]
  PIN prt2_dir[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.3205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4102 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 808.125000 0.000000 808.225000 0.520000 ;
    END
  END prt2_dir[1]
  PIN prt2_dir[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.691 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 3.402 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0128 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 893.925000 0.000000 894.025000 0.520000 ;
    END
  END prt2_dir[0]
  PIN prt2_ren[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4405 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9382 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.306 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.9904 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 297.285000 0.000000 297.385000 0.520000 ;
    END
  END prt2_ren[7]
  PIN prt2_ren[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6405 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8182 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 7.586 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.4224 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 383.085000 0.000000 383.185000 0.520000 ;
    END
  END prt2_ren[6]
  PIN prt2_ren[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5005 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2022 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 10.642 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.8688 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 468.885000 0.000000 468.985000 0.520000 ;
    END
  END prt2_ren[5]
  PIN prt2_ren[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1035 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4554 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.782 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8848 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 554.685000 0.000000 554.785000 0.520000 ;
    END
  END prt2_ren[4]
  PIN prt2_ren[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.5125 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.299 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 640.485000 0.000000 640.585000 0.520000 ;
    END
  END prt2_ren[3]
  PIN prt2_ren[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.6855 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0602 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 726.285000 0.000000 726.385000 0.520000 ;
    END
  END prt2_ren[2]
  PIN prt2_ren[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9414 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 812.085000 0.000000 812.185000 0.520000 ;
    END
  END prt2_ren[1]
  PIN prt2_ren[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4475 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.969 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 7.606 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.5104 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 897.885000 0.000000 897.985000 0.520000 ;
    END
  END prt2_ren[0]
  PIN prt3_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3285 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.9334 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2  ;
    ANTENNAMAXAREACAR 604.142 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 2660.01 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.369004 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 641.335000 0.520000 641.435000 ;
    END
  END prt3_in[7]
  PIN prt3_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1085 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.3654 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2  ;
    ANTENNAMAXAREACAR 267.399 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 1176.52 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.738007 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 553.335000 0.520000 553.435000 ;
    END
  END prt3_in[6]
  PIN prt3_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9725 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.679 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 17.068 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.1872 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 2.942 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9888 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4  ;
    ANTENNAMAXAREACAR 46.3931 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 195.149 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 465.335000 0.520000 465.435000 ;
    END
  END prt3_in[5]
  PIN prt3_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6125 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.695 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 10.802 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.5728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 6.406 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 28.2304 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M5  ;
    ANTENNAMAXAREACAR 68.5185 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 302.549 LAYER M5  ;
    ANTENNAMAXCUTCAR 0.780649 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 377.335000 0.520000 377.435000 ;
    END
  END prt3_in[4]
  PIN prt3_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2135 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3834 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 10.242 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1088 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 543.312 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 2392.36 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 289.335000 0.520000 289.435000 ;
    END
  END prt3_in[3]
  PIN prt3_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.2135 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.5834 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 14.306 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.9904 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 552.177 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 2422.64 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 201.335000 0.520000 201.435000 ;
    END
  END prt3_in[2]
  PIN prt3_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.3605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.2302 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2  ;
    ANTENNAMAXAREACAR 718.173 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 3158.84 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.738007 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 113.335000 0.520000 113.435000 ;
    END
  END prt3_in[1]
  PIN prt3_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1325 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.383 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 9.518 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.9232 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3  ;
    ANTENNAMAXAREACAR 294.334 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1280.41 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 25.335000 0.520000 25.435000 ;
    END
  END prt3_in[0]
  PIN prt3_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.156 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.6864 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.778 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4672 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 661.570000 0.520000 661.670000 ;
    END
  END prt3_out[7]
  PIN prt3_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 6.463 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.5252 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 573.570000 0.520000 573.670000 ;
    END
  END prt3_out[6]
  PIN prt3_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.316 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 15.978 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3472 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 485.570000 0.520000 485.670000 ;
    END
  END prt3_out[5]
  PIN prt3_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.782 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.0848 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 397.570000 0.520000 397.670000 ;
    END
  END prt3_out[4]
  PIN prt3_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.542 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.0288 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 309.570000 0.520000 309.670000 ;
    END
  END prt3_out[3]
  PIN prt3_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.952 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.1888 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 5.506 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.2704 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 221.570000 0.520000 221.670000 ;
    END
  END prt3_out[2]
  PIN prt3_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 13.355 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.85 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 133.570000 0.520000 133.670000 ;
    END
  END prt3_out[1]
  PIN prt3_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.901 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2084 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 45.570000 0.520000 45.670000 ;
    END
  END prt3_out[0]
  PIN prt3_dir[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 13.8795 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.1578 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 650.975000 0.520000 651.075000 ;
    END
  END prt3_dir[7]
  PIN prt3_dir[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.8595 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.4698 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 562.975000 0.520000 563.075000 ;
    END
  END prt3_dir[6]
  PIN prt3_dir[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 7.0995 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.3258 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 474.975000 0.520000 475.075000 ;
    END
  END prt3_dir[5]
  PIN prt3_dir[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2365 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0406 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.778 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.0672 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 386.975000 0.520000 387.075000 ;
    END
  END prt3_dir[4]
  PIN prt3_dir[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1315 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.606 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.3104 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 298.975000 0.520000 299.075000 ;
    END
  END prt3_dir[3]
  PIN prt3_dir[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 14.4545 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.6878 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 210.975000 0.520000 211.075000 ;
    END
  END prt3_dir[2]
  PIN prt3_dir[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 13.9565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.5406 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 122.975000 0.520000 123.075000 ;
    END
  END prt3_dir[1]
  PIN prt3_dir[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 2.9915 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2506 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 34.975000 0.520000 35.075000 ;
    END
  END prt3_dir[0]
  PIN prt3_ren[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 13.9235 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.3514 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 647.015000 0.520000 647.115000 ;
    END
  END prt3_ren[7]
  PIN prt3_ren[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1185 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.5654 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.058 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0992 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 559.015000 0.520000 559.115000 ;
    END
  END prt3_ren[6]
  PIN prt3_ren[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 6.582 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.0048 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 471.015000 0.520000 471.115000 ;
    END
  END prt3_ren[5]
  PIN prt3_ren[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4405 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9382 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.84 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.384 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0582 LAYER M3  ;
    ANTENNAMAXAREACAR 257.015 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1131.59 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.343643 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 383.015000 0.520000 383.115000 ;
    END
  END prt3_ren[4]
  PIN prt3_ren[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2875 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.665 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 5.662 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9568 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 295.015000 0.520000 295.115000 ;
    END
  END prt3_ren[3]
  PIN prt3_ren[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 6.3085 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.8894 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 207.015000 0.520000 207.115000 ;
    END
  END prt3_ren[2]
  PIN prt3_ren[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 14.3105 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.0542 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 119.015000 0.520000 119.115000 ;
    END
  END prt3_ren[1]
  PIN prt3_ren[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 2.7035 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9834 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 31.015000 0.520000 31.115000 ;
    END
  END prt3_ren[0]
  PIN prt4_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9385 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1294 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 24.786 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.102 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 953.358 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 4183.32 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 646.165000 685.480000 646.265000 686.000000 ;
    END
  END prt4_in[7]
  PIN prt4_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6755 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3722 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 18.618 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.9632 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 3.982 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5648 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M6  ;
    ANTENNAMAXAREACAR 82.445 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 364.755 LAYER M6  ;
    ANTENNAMAXCUTCAR 2.01137 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 560.365000 685.480000 560.465000 686.000000 ;
    END
  END prt4_in[6]
  PIN prt4_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9385 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5294 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 8.932 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.3888 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 4.156 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.3744 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4  ;
    ANTENNAMAXAREACAR 99.0087 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 439.603 LAYER M4  ;
    ANTENNAMAXCUTCAR 2.43902 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 474.565000 685.480000 474.665000 686.000000 ;
    END
  END prt4_in[5]
  PIN prt4_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3185 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8014 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.702 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5328 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 7.262 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 31.9968 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M6  ;
    ANTENNAMAXAREACAR 85.6804 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 366.922 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.66205 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 388.765000 685.480000 388.865000 686.000000 ;
    END
  END prt4_in[4]
  PIN prt4_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 14.036 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.6156 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 1.84 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 LAYER M4  ;
    ANTENNAMAXAREACAR 9.25236 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 13.0747 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.235849 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 302.965000 685.480000 303.065000 686.000000 ;
    END
  END prt4_in[3]
  PIN prt4_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8325 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.663 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 11.986 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.7824 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 8.062 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.5168 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M4  ;
    ANTENNAMAXAREACAR 257.184 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 1134.36 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.44092 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 217.165000 685.480000 217.265000 686.000000 ;
    END
  END prt4_in[2]
  PIN prt4_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.174 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1914 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.244 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4444 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.164 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3564 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.164 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3564 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 69.44 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 76.736 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M6  ;
    ANTENNAMAXAREACAR 587.083 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 655.811 LAYER M6  ;
    ANTENNAMAXCUTCAR 0.707547 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 131.365000 685.480000 131.465000 686.000000 ;
    END
  END prt4_in[1]
  PIN prt4_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1905 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.0822 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2  ;
    ANTENNAMAXAREACAR 240.504 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 1056.8 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 45.565000 685.480000 45.665000 686.000000 ;
    END
  END prt4_in[0]
  PIN prt4_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.14 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4134 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 66.752 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.6032 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 625.930000 685.480000 626.030000 686.000000 ;
    END
  END prt4_out[7]
  PIN prt4_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.572 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0886 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 36.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.656 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 540.130000 685.480000 540.230000 686.000000 ;
    END
  END prt4_out[6]
  PIN prt4_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.172 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 12.162 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5542 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 454.330000 685.480000 454.430000 686.000000 ;
    END
  END prt4_out[5]
  PIN prt4_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.446 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4906 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 5.2 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.072 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 368.530000 685.480000 368.630000 686.000000 ;
    END
  END prt4_out[4]
  PIN prt4_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.939 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1316 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.968 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 5.922 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.1008 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 282.730000 685.480000 282.830000 686.000000 ;
    END
  END prt4_out[3]
  PIN prt4_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.619 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7236 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.266 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.8144 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 196.930000 685.480000 197.030000 686.000000 ;
    END
  END prt4_out[2]
  PIN prt4_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.742 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 73.7088 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 111.130000 685.480000 111.230000 686.000000 ;
    END
  END prt4_out[1]
  PIN prt4_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 25.330000 685.480000 25.430000 686.000000 ;
    END
  END prt4_out[0]
  PIN prt4_dir[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.3015 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3706 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 636.525000 685.480000 636.625000 686.000000 ;
    END
  END prt4_dir[7]
  PIN prt4_dir[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.3165 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4366 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 550.725000 685.480000 550.825000 686.000000 ;
    END
  END prt4_dir[6]
  PIN prt4_dir[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 5.7785 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.5134 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 464.925000 685.480000 465.025000 686.000000 ;
    END
  END prt4_dir[5]
  PIN prt4_dir[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.2545 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1198 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 379.125000 685.480000 379.225000 686.000000 ;
    END
  END prt4_dir[4]
  PIN prt4_dir[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.851 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7444 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.968 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 4.978 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.9472 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 293.325000 685.480000 293.425000 686.000000 ;
    END
  END prt4_dir[3]
  PIN prt4_dir[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.691 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 13.722 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.4208 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 207.525000 685.480000 207.625000 686.000000 ;
    END
  END prt4_dir[2]
  PIN prt4_dir[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.722 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 73.6208 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 121.725000 685.480000 121.825000 686.000000 ;
    END
  END prt4_dir[1]
  PIN prt4_dir[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.386 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 72.1424 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 35.925000 685.480000 36.025000 686.000000 ;
    END
  END prt4_dir[0]
  PIN prt4_ren[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.4965 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2286 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 640.485000 685.480000 640.585000 686.000000 ;
    END
  END prt4_ren[7]
  PIN prt4_ren[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.3475 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.017 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 554.685000 685.480000 554.785000 686.000000 ;
    END
  END prt4_ren[6]
  PIN prt4_ren[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5305 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7342 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 7.862 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.6368 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 468.885000 685.480000 468.985000 686.000000 ;
    END
  END prt4_ren[5]
  PIN prt4_ren[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 2.5585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3014 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 383.085000 685.480000 383.185000 686.000000 ;
    END
  END prt4_ren[4]
  PIN prt4_ren[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7635 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3594 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 4.142 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2688 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 297.285000 685.480000 297.385000 686.000000 ;
    END
  END prt4_ren[3]
  PIN prt4_ren[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9035 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9754 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 12.822 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.4608 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 211.485000 685.480000 211.585000 686.000000 ;
    END
  END prt4_ren[2]
  PIN prt4_ren[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9035 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9754 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.086 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8224 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 15.802 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 69.5728 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 125.685000 685.480000 125.785000 686.000000 ;
    END
  END prt4_ren[1]
  PIN prt4_ren[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.842 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7488 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 39.885000 685.480000 39.985000 686.000000 ;
    END
  END prt4_ren[0]
  PIN use_dac_glb_bias
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1505 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6622 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.986 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3824 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.158 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7392 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.826 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8784 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 10.696 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 47.1504 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 614.515000 389.000000 614.615000 ;
    END
  END use_dac_glb_bias
  PIN en_bias_buf
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.081 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 613.970000 389.000000 614.070000 ;
    END
  END en_bias_buf
  PIN en_bias_gen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.041 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1804 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 612.880000 389.000000 612.980000 ;
    END
  END en_bias_gen
  PIN BIAS_ADJ[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.051 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2244 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.186 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4624 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 10.738 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 47.2912 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 609.610000 389.000000 609.710000 ;
    END
  END BIAS_ADJ[5]
  PIN BIAS_ADJ[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0965 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4246 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.786 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5024 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.886 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9424 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.858 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 43.4192 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 610.155000 389.000000 610.255000 ;
    END
  END BIAS_ADJ[4]
  PIN BIAS_ADJ[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.476 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1824 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 610.700000 389.000000 610.800000 ;
    END
  END BIAS_ADJ[3]
  PIN BIAS_ADJ[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6855 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0602 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 611.245000 389.000000 611.345000 ;
    END
  END BIAS_ADJ[2]
  PIN BIAS_ADJ[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.358 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.178 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.326 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 19.0784 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 10.978 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 48.3472 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 611.790000 389.000000 611.890000 ;
    END
  END BIAS_ADJ[1]
  PIN BIAS_ADJ[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.518 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3232 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 1.002 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4528 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 11.758 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 51.7792 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 612.335000 389.000000 612.435000 ;
    END
  END BIAS_ADJ[0]
  PIN BIAS_DBP[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.142 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2688 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 10.36 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 45.672 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 601.980000 389.000000 602.080000 ;
    END
  END BIAS_DBP[13]
  PIN BIAS_DBP[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.818 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0432 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 2.406 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6304 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.878 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 43.5072 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 602.525000 389.000000 602.625000 ;
    END
  END BIAS_DBP[12]
  PIN BIAS_DBP[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.118 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.726 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4384 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.558 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 42.0992 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 603.070000 389.000000 603.170000 ;
    END
  END BIAS_DBP[11]
  PIN BIAS_DBP[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.2125 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.979 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 603.615000 389.000000 603.715000 ;
    END
  END BIAS_DBP[10]
  PIN BIAS_DBP[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.726 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4384 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 8.598 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 37.8752 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 604.160000 389.000000 604.260000 ;
    END
  END BIAS_DBP[9]
  PIN BIAS_DBP[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0185 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0814 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.318 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4432 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 604.705000 389.000000 604.805000 ;
    END
  END BIAS_DBP[8]
  PIN BIAS_DBP[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.402 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.826 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8784 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 11.102 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 48.8928 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 605.250000 389.000000 605.350000 ;
    END
  END BIAS_DBP[7]
  PIN BIAS_DBP[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.986 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3824 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.442 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1888 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 10.338 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 45.5312 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 605.795000 389.000000 605.895000 ;
    END
  END BIAS_DBP[6]
  PIN BIAS_DBP[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.302 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9152 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.306 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5904 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 11.202 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 49.3328 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 606.340000 389.000000 606.440000 ;
    END
  END BIAS_DBP[5]
  PIN BIAS_DBP[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.802 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.218 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6032 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.638 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 42.4512 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 606.885000 389.000000 606.985000 ;
    END
  END BIAS_DBP[4]
  PIN BIAS_DBP[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.069 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3036 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.686 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0624 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.302 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 11.002 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 48.4528 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 607.430000 389.000000 607.530000 ;
    END
  END BIAS_DBP[3]
  PIN BIAS_DBP[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.546 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 20.0464 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 11.378 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 50.1072 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 607.975000 389.000000 608.075000 ;
    END
  END BIAS_DBP[2]
  PIN BIAS_DBP[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 2.018 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9232 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 0.106 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 608.520000 389.000000 608.620000 ;
    END
  END BIAS_DBP[1]
  PIN BIAS_DBP[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0275 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.165 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 609.065000 389.000000 609.165000 ;
    END
  END BIAS_DBP[0]
  PIN BIAS_DBN[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 5.993 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.4132 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 579.090000 389.000000 579.190000 ;
    END
  END BIAS_DBN[13]
  PIN BIAS_DBN[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0255 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1122 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.482 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5648 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.922 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1008 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.226 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 7.138 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 31.4512 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 579.635000 389.000000 579.735000 ;
    END
  END BIAS_DBN[12]
  PIN BIAS_DBN[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 580.180000 389.000000 580.280000 ;
    END
  END BIAS_DBN[11]
  PIN BIAS_DBN[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 580.725000 389.000000 580.825000 ;
    END
  END BIAS_DBN[10]
  PIN BIAS_DBN[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.491 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2044 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 581.270000 389.000000 581.370000 ;
    END
  END BIAS_DBN[9]
  PIN BIAS_DBN[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 581.815000 389.000000 581.915000 ;
    END
  END BIAS_DBN[8]
  PIN BIAS_DBN[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.442 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.826 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9224 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.968 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 8.626 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 38.0864 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 582.360000 389.000000 582.460000 ;
    END
  END BIAS_DBN[7]
  PIN BIAS_DBN[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9315 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1426 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.226 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4384 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 2.698 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9152 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 582.905000 389.000000 583.005000 ;
    END
  END BIAS_DBN[6]
  PIN BIAS_DBN[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 5.158 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.7392 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 3.738 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4912 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 583.450000 389.000000 583.550000 ;
    END
  END BIAS_DBN[5]
  PIN BIAS_DBN[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0295 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1298 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.666 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3744 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 2.118 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3632 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 6.438 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 28.3712 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 583.995000 389.000000 584.095000 ;
    END
  END BIAS_DBN[4]
  PIN BIAS_DBN[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.211 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.1724 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 584.540000 389.000000 584.640000 ;
    END
  END BIAS_DBN[3]
  PIN BIAS_DBN[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.418 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8832 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 1.182 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2448 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 585.085000 389.000000 585.185000 ;
    END
  END BIAS_DBN[2]
  PIN BIAS_DBN[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.748 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7792 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 4.362 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2368 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 3.518 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5232 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 585.630000 389.000000 585.730000 ;
    END
  END BIAS_DBN[1]
  PIN BIAS_DBN[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0795 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3498 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 4.346 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.1664 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 6.518 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.7232 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.968 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 3.438 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1712 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 586.175000 389.000000 586.275000 ;
    END
  END BIAS_DBN[0]
  PIN BIAS_DBPC[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.194 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8536 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.582 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6048 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 594.350000 389.000000 594.450000 ;
    END
  END BIAS_DBPC[13]
  PIN BIAS_DBPC[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.4715 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1626 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 594.895000 389.000000 594.995000 ;
    END
  END BIAS_DBPC[12]
  PIN BIAS_DBPC[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0624 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 595.440000 389.000000 595.540000 ;
    END
  END BIAS_DBPC[11]
  PIN BIAS_DBPC[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.1555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7282 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 595.985000 389.000000 596.085000 ;
    END
  END BIAS_DBPC[10]
  PIN BIAS_DBPC[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.032 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1408 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.762 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3968 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 596.530000 389.000000 596.630000 ;
    END
  END BIAS_DBPC[9]
  PIN BIAS_DBPC[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.246 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.146 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2864 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 10.138 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 44.6512 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 597.075000 389.000000 597.175000 ;
    END
  END BIAS_DBPC[8]
  PIN BIAS_DBPC[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6336 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.906 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0304 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 597.620000 389.000000 597.720000 ;
    END
  END BIAS_DBPC[7]
  PIN BIAS_DBPC[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.5395 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4618 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 598.165000 389.000000 598.265000 ;
    END
  END BIAS_DBPC[6]
  PIN BIAS_DBPC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.742 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3088 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 598.710000 389.000000 598.810000 ;
    END
  END BIAS_DBPC[5]
  PIN BIAS_DBPC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.258 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 599.255000 389.000000 599.355000 ;
    END
  END BIAS_DBPC[4]
  PIN BIAS_DBPC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.019 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0836 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 599.800000 389.000000 599.900000 ;
    END
  END BIAS_DBPC[3]
  PIN BIAS_DBPC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 600.345000 389.000000 600.445000 ;
    END
  END BIAS_DBPC[2]
  PIN BIAS_DBPC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 7.978 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.1472 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 600.890000 389.000000 600.990000 ;
    END
  END BIAS_DBPC[1]
  PIN BIAS_DBPC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.2875 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.309 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 601.435000 389.000000 601.535000 ;
    END
  END BIAS_DBPC[0]
  PIN BIAS_DBNC[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 5.378 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.7072 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 586.720000 389.000000 586.820000 ;
    END
  END BIAS_DBNC[13]
  PIN BIAS_DBNC[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 8.138 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.8512 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 587.265000 389.000000 587.365000 ;
    END
  END BIAS_DBNC[12]
  PIN BIAS_DBNC[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 6.643 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.3172 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 587.810000 389.000000 587.910000 ;
    END
  END BIAS_DBNC[11]
  PIN BIAS_DBNC[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.438 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3712 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 7.238 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.8912 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 588.355000 389.000000 588.455000 ;
    END
  END BIAS_DBNC[10]
  PIN BIAS_DBNC[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.274 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2496 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 588.900000 389.000000 589.000000 ;
    END
  END BIAS_DBNC[9]
  PIN BIAS_DBNC[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.616 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7984 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 589.445000 389.000000 589.545000 ;
    END
  END BIAS_DBNC[8]
  PIN BIAS_DBNC[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.482 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5648 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.418 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8832 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.792 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.084 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 40.0576 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6  ;
    ANTENNAMAXAREACAR 440.871 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1946.74 LAYER M6  ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 589.990000 389.000000 590.090000 ;
    END
  END BIAS_DBNC[7]
  PIN BIAS_DBNC[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.894 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4656 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 4.838 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3312 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M4  ;
    ANTENNAMAXAREACAR 139.622 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 616.778 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.02881 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 590.535000 389.000000 590.635000 ;
    END
  END BIAS_DBNC[6]
  PIN BIAS_DBNC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.506 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6704 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.118 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 2.842 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5488 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 10.542 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 46.4288 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 591.080000 389.000000 591.180000 ;
    END
  END BIAS_DBNC[5]
  PIN BIAS_DBNC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0695 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3058 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 9.302 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.9728 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 591.625000 389.000000 591.725000 ;
    END
  END BIAS_DBNC[4]
  PIN BIAS_DBNC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.258 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.838 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9312 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.968 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.678 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 42.6272 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 592.170000 389.000000 592.270000 ;
    END
  END BIAS_DBNC[3]
  PIN BIAS_DBNC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.982 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3648 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.526 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5584 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.102 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 40.0928 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M6  ;
    ANTENNAMAXAREACAR 298.459 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1317.47 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 592.715000 389.000000 592.815000 ;
    END
  END BIAS_DBNC[2]
  PIN BIAS_DBNC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.09 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.44 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 593.260000 389.000000 593.360000 ;
    END
  END BIAS_DBNC[1]
  PIN BIAS_DBNC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0195 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.162 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1568 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.498 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4352 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 10.904 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 48.0656 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6  ;
    ANTENNAMAXAREACAR 196.443 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 863.625 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.2987 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 388.480000 593.805000 389.000000 593.905000 ;
    END
  END BIAS_DBNC[0]
  PIN BIAS_TC_POT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.1395 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6578 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.266 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2144 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 0.258 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5  ;
    ANTENNAMAXAREACAR 28.097 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 125.974 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1052.065000 445.480000 1052.165000 446.000000 ;
    END
  END BIAS_TC_POT[5]
  PIN BIAS_TC_POT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.663 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9172 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1052.610000 445.480000 1052.710000 446.000000 ;
    END
  END BIAS_TC_POT[4]
  PIN BIAS_TC_POT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.434 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3536 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4  ;
    ANTENNAMAXAREACAR 25.5934 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 114.323 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1053.155000 445.480000 1053.255000 446.000000 ;
    END
  END BIAS_TC_POT[3]
  PIN BIAS_TC_POT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.482 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6528 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2  ;
    ANTENNAMAXAREACAR 41.6701 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 186.59 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.273224 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 1053.700000 445.480000 1053.800000 446.000000 ;
    END
  END BIAS_TC_POT[2]
  PIN BIAS_TC_POT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3265 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4366 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.358 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.458 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1054.245000 445.480000 1054.345000 446.000000 ;
    END
  END BIAS_TC_POT[1]
  PIN BIAS_TC_POT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.142 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.346 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5  ;
    ANTENNAMAXAREACAR 19.7926 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 89.4343 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1054.790000 445.480000 1054.890000 446.000000 ;
    END
  END BIAS_TC_POT[0]
  PIN BIAS_LC_POT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.9385 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1294 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1055.335000 445.480000 1055.435000 446.000000 ;
    END
  END BIAS_LC_POT[5]
  PIN BIAS_LC_POT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.079 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3916 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.832 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1488 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M4  ;
    ANTENNAMAXAREACAR 62.7254 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 278.497 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.36612 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1055.880000 445.480000 1055.980000 446.000000 ;
    END
  END BIAS_LC_POT[4]
  PIN BIAS_LC_POT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.522 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3408 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1056.425000 445.480000 1056.525000 446.000000 ;
    END
  END BIAS_LC_POT[3]
  PIN BIAS_LC_POT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3608 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.302 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7728 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M4  ;
    ANTENNAMAXAREACAR 78.8456 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 348.224 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.0929 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1056.970000 445.480000 1057.070000 446.000000 ;
    END
  END BIAS_LC_POT[2]
  PIN BIAS_LC_POT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6662 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.332 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9488 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3  ;
    ANTENNAMAXAREACAR 30.5263 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 133.583 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1057.515000 445.480000 1057.615000 446.000000 ;
    END
  END BIAS_LC_POT[1]
  PIN BIAS_LC_POT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.848 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7312 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.874 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8896 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 15.5303 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 68.1501 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1058.060000 445.480000 1058.160000 446.000000 ;
    END
  END BIAS_LC_POT[0]
  PIN BIAS_TIA_G_POT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.094 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4136 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 5.862 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.8368 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1059.150000 445.480000 1059.250000 446.000000 ;
    END
  END BIAS_TIA_G_POT[16]
  PIN BIAS_TIA_G_POT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.551 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4244 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 5.458 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 24.0592 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1043.345000 445.480000 1043.445000 446.000000 ;
    END
  END BIAS_TIA_G_POT[15]
  PIN BIAS_TIA_G_POT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.487 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2308 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1043.890000 445.480000 1043.990000 446.000000 ;
    END
  END BIAS_TIA_G_POT[14]
  PIN BIAS_TIA_G_POT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 4.882 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.5248 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1044.435000 445.480000 1044.535000 446.000000 ;
    END
  END BIAS_TIA_G_POT[13]
  PIN BIAS_TIA_G_POT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.231 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0164 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 5.102 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4928 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1044.980000 445.480000 1045.080000 446.000000 ;
    END
  END BIAS_TIA_G_POT[12]
  PIN BIAS_TIA_G_POT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.2595 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5418 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1045.525000 445.480000 1045.625000 446.000000 ;
    END
  END BIAS_TIA_G_POT[11]
  PIN BIAS_TIA_G_POT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.473 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0812 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1046.070000 445.480000 1046.170000 446.000000 ;
    END
  END BIAS_TIA_G_POT[10]
  PIN BIAS_TIA_G_POT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.6435 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8314 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1046.615000 445.480000 1046.715000 446.000000 ;
    END
  END BIAS_TIA_G_POT[9]
  PIN BIAS_TIA_G_POT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1047.160000 445.480000 1047.260000 446.000000 ;
    END
  END BIAS_TIA_G_POT[8]
  PIN BIAS_TIA_G_POT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3965 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7446 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4112 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.84 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.228 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 32.702 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 143.933 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 5.276 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3024 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6  ;
    ANTENNAMAXAREACAR 199.834 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 883.09 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.33333 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 1047.705000 445.480000 1047.805000 446.000000 ;
    END
  END BIAS_TIA_G_POT[7]
  PIN BIAS_TIA_G_POT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.807 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5508 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.424 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3536 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.242 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5088 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 34.662 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 152.557 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0481 LAYER M5  ;
    ANTENNAMAXAREACAR 769.899 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 3390.14 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.4553 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1048.250000 445.480000 1048.350000 446.000000 ;
    END
  END BIAS_TIA_G_POT[6]
  PIN BIAS_TIA_G_POT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4574 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.446 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4064 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1048.795000 445.480000 1048.895000 446.000000 ;
    END
  END BIAS_TIA_G_POT[5]
  PIN BIAS_TIA_G_POT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.353 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5972 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1049.340000 445.480000 1049.440000 446.000000 ;
    END
  END BIAS_TIA_G_POT[4]
  PIN BIAS_TIA_G_POT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.0898 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.682 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4448 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4  ;
    ANTENNAMAXAREACAR 58.3424 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 259.053 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1049.885000 445.480000 1049.985000 446.000000 ;
    END
  END BIAS_TIA_G_POT[3]
  PIN BIAS_TIA_G_POT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.278 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1050.430000 445.480000 1050.530000 446.000000 ;
    END
  END BIAS_TIA_G_POT[2]
  PIN BIAS_TIA_G_POT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3385 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4894 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.898 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9952 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1050.975000 445.480000 1051.075000 446.000000 ;
    END
  END BIAS_TIA_G_POT[1]
  PIN BIAS_TIA_G_POT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.171 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7524 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.418 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2832 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 36.7551 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 162.799 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1051.520000 445.480000 1051.620000 446.000000 ;
    END
  END BIAS_TIA_G_POT[0]
  PIN BIAS_REV_POT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.558 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8992 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 607.010000 1139.520000 607.110000 ;
    END
  END BIAS_REV_POT[13]
  PIN BIAS_REV_POT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 607.555000 1139.520000 607.655000 ;
    END
  END BIAS_REV_POT[12]
  PIN BIAS_REV_POT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.147 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2908 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 608.100000 1139.520000 608.200000 ;
    END
  END BIAS_REV_POT[11]
  PIN BIAS_REV_POT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1675 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.737 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.986 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3824 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 608.645000 1139.520000 608.745000 ;
    END
  END BIAS_REV_POT[10]
  PIN BIAS_REV_POT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 609.190000 1139.520000 609.290000 ;
    END
  END BIAS_REV_POT[9]
  PIN BIAS_REV_POT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3105 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.4102 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.506 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2704 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 609.735000 1139.520000 609.835000 ;
    END
  END BIAS_REV_POT[8]
  PIN BIAS_REV_POT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.592 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6928 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 610.280000 1139.520000 610.380000 ;
    END
  END BIAS_REV_POT[7]
  PIN BIAS_REV_POT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0215 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0946 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.802 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5728 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 610.825000 1139.520000 610.925000 ;
    END
  END BIAS_REV_POT[6]
  PIN BIAS_REV_POT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.597 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6708 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 611.370000 1139.520000 611.470000 ;
    END
  END BIAS_REV_POT[5]
  PIN BIAS_REV_POT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.276 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 611.915000 1139.520000 612.015000 ;
    END
  END BIAS_REV_POT[4]
  PIN BIAS_REV_POT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.692 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.442 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 612.460000 1139.520000 612.560000 ;
    END
  END BIAS_REV_POT[3]
  PIN BIAS_REV_POT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.2425 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.155 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 613.005000 1139.520000 613.105000 ;
    END
  END BIAS_REV_POT[2]
  PIN BIAS_REV_POT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.838 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7312 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 613.550000 1139.520000 613.650000 ;
    END
  END BIAS_REV_POT[1]
  PIN BIAS_REV_POT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0395 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1738 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.862 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8368 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 614.095000 1139.520000 614.195000 ;
    END
  END BIAS_REV_POT[0]
  PIN BIAS_TC_DSADC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8755 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8522 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 10.7973 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 47.3247 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1019.335000 445.480000 1019.435000 446.000000 ;
    END
  END BIAS_TC_DSADC[5]
  PIN BIAS_TC_DSADC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.69 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.036 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1019.880000 445.480000 1019.980000 446.000000 ;
    END
  END BIAS_TC_DSADC[4]
  PIN BIAS_TC_DSADC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1135 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8994 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.982 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3648 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 25.956 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 113.198 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1020.425000 445.480000 1020.525000 446.000000 ;
    END
  END BIAS_TC_DSADC[3]
  PIN BIAS_TC_DSADC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.271 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1924 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1020.970000 445.480000 1021.070000 446.000000 ;
    END
  END BIAS_TC_DSADC[2]
  PIN BIAS_TC_DSADC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.3425 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.951 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1021.515000 445.480000 1021.615000 446.000000 ;
    END
  END BIAS_TC_DSADC[1]
  PIN BIAS_TC_DSADC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.646 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8424 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.518 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3232 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 17.601 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 77.4978 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.2886 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1022.060000 445.480000 1022.160000 446.000000 ;
    END
  END BIAS_TC_DSADC[0]
  PIN BIAS_LC_DSADC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.7179 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3018 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3  ;
    ANTENNAMAXAREACAR 17.1994 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 73.4401 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.647249 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1022.605000 445.480000 1022.705000 446.000000 ;
    END
  END BIAS_LC_DSADC[5]
  PIN BIAS_LC_DSADC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.471 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0724 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.838 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7312 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 2.47 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.912 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4  ;
    ANTENNAMAXAREACAR 120.551 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 530.337 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1023.150000 445.480000 1023.250000 446.000000 ;
    END
  END BIAS_LC_DSADC[4]
  PIN BIAS_LC_DSADC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7715 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3946 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.898 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3952 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3  ;
    ANTENNAMAXAREACAR 73.1254 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 318.498 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1023.695000 445.480000 1023.795000 446.000000 ;
    END
  END BIAS_LC_DSADC[3]
  PIN BIAS_LC_DSADC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.49 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1024.240000 445.480000 1024.340000 446.000000 ;
    END
  END BIAS_LC_DSADC[2]
  PIN BIAS_LC_DSADC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.0005 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4902 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1024.785000 445.480000 1024.885000 446.000000 ;
    END
  END BIAS_LC_DSADC[1]
  PIN BIAS_LC_DSADC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.416 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8304 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9152 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.646 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8864 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4  ;
    ANTENNAMAXAREACAR 35.1912 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 152.805 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1025.330000 445.480000 1025.430000 446.000000 ;
    END
  END BIAS_LC_DSADC[0]
  PIN BIAS_RIN_DSADC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2685 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5814 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.072 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3  ;
    ANTENNAMAXAREACAR 23.8091 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 106.466 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1016.065000 445.480000 1016.165000 446.000000 ;
    END
  END BIAS_RIN_DSADC[5]
  PIN BIAS_RIN_DSADC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.371 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6324 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.122 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9808 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.138 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6512 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4  ;
    ANTENNAMAXAREACAR 29.0906 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 130.641 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1016.610000 445.480000 1016.710000 446.000000 ;
    END
  END BIAS_RIN_DSADC[4]
  PIN BIAS_RIN_DSADC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.382 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1248 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.226 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4  ;
    ANTENNAMAXAREACAR 12.9094 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 59.4434 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAMAXCUTCAR 2.26537 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M5  ;
    ANTENNAGATEAREA 0.0309 LAYER M5  ;
    ANTENNAMAXAREACAR 20.6117 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 94.7573 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 1.546 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8464 LAYER M6  ;
    ANTENNAGATEAREA 0.0309 LAYER M6  ;
    ANTENNAMAXAREACAR 70.644 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 316.324 LAYER M6  ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 1017.155000 445.480000 1017.255000 446.000000 ;
    END
  END BIAS_RIN_DSADC[3]
  PIN BIAS_RIN_DSADC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.356 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9664 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.064 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1696 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 35.0595 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 155.974 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1017.700000 445.480000 1017.800000 446.000000 ;
    END
  END BIAS_RIN_DSADC[2]
  PIN BIAS_RIN_DSADC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3875 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.105 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.804 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0256 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3  ;
    ANTENNAMAXAREACAR 89.3495 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 395.78 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1018.245000 445.480000 1018.345000 446.000000 ;
    END
  END BIAS_RIN_DSADC[1]
  PIN BIAS_RIN_DSADC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.493 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2132 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1018.790000 445.480000 1018.890000 446.000000 ;
    END
  END BIAS_RIN_DSADC[0]
  PIN BIAS_RFB_DSADC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.2445 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5198 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 LAYER M2  ;
    ANTENNAMAXAREACAR 23.2979 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 102.273 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.35461 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 1012.795000 445.480000 1012.895000 446.000000 ;
    END
  END BIAS_RFB_DSADC[5]
  PIN BIAS_RFB_DSADC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.091 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 3.824 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9136 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.422 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9008 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 27.376 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 120.542 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 4.584 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 20.2576 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6  ;
    ANTENNAMAXAREACAR 179.329 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 791.265 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 1013.340000 445.480000 1013.440000 446.000000 ;
    END
  END BIAS_RFB_DSADC[4]
  PIN BIAS_RFB_DSADC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.693 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0932 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1013.885000 445.480000 1013.985000 446.000000 ;
    END
  END BIAS_RFB_DSADC[3]
  PIN BIAS_RFB_DSADC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.369 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6236 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 6.33 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.896 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 11.258 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 49.5792 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5  ;
    ANTENNAMAXAREACAR 232.015 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 1017.14 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1014.430000 445.480000 1014.530000 446.000000 ;
    END
  END BIAS_RFB_DSADC[2]
  PIN BIAS_RFB_DSADC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0945 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4158 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.118 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1014.975000 445.480000 1015.075000 446.000000 ;
    END
  END BIAS_RFB_DSADC[1]
  PIN BIAS_RFB_DSADC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.111 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4884 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.482 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1648 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 2.682 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8448 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M5  ;
    ANTENNAMAXAREACAR 463.304 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 2040.85 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.589 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1015.520000 445.480000 1015.620000 446.000000 ;
    END
  END BIAS_RFB_DSADC[0]
  PIN BIAS_DSADC_VCM[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.266 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2144 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 599.380000 1139.520000 599.480000 ;
    END
  END BIAS_DSADC_VCM[13]
  PIN BIAS_DSADC_VCM[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.338 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9312 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 599.925000 1139.520000 600.025000 ;
    END
  END BIAS_DSADC_VCM[12]
  PIN BIAS_DSADC_VCM[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.626 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.7984 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.586 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6224 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 600.470000 1139.520000 600.570000 ;
    END
  END BIAS_DSADC_VCM[11]
  PIN BIAS_DSADC_VCM[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 6.2835 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6474 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 601.015000 1139.520000 601.115000 ;
    END
  END BIAS_DSADC_VCM[10]
  PIN BIAS_DSADC_VCM[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.298 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3552 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 601.560000 1139.520000 601.660000 ;
    END
  END BIAS_DSADC_VCM[9]
  PIN BIAS_DSADC_VCM[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.564 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5696 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 602.105000 1139.520000 602.205000 ;
    END
  END BIAS_DSADC_VCM[8]
  PIN BIAS_DSADC_VCM[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 602.650000 1139.520000 602.750000 ;
    END
  END BIAS_DSADC_VCM[7]
  PIN BIAS_DSADC_VCM[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.522 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3408 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 603.195000 1139.520000 603.295000 ;
    END
  END BIAS_DSADC_VCM[6]
  PIN BIAS_DSADC_VCM[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 603.740000 1139.520000 603.840000 ;
    END
  END BIAS_DSADC_VCM[5]
  PIN BIAS_DSADC_VCM[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.692 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.482 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1648 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 604.285000 1139.520000 604.385000 ;
    END
  END BIAS_DSADC_VCM[4]
  PIN BIAS_DSADC_VCM[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 604.830000 1139.520000 604.930000 ;
    END
  END BIAS_DSADC_VCM[3]
  PIN BIAS_DSADC_VCM[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.318 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8432 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 605.375000 1139.520000 605.475000 ;
    END
  END BIAS_DSADC_VCM[2]
  PIN BIAS_DSADC_VCM[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.562 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5168 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 605.920000 1139.520000 606.020000 ;
    END
  END BIAS_DSADC_VCM[1]
  PIN BIAS_DSADC_VCM[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0275 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.165 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 606.465000 1139.520000 606.565000 ;
    END
  END BIAS_DSADC_VCM[0]
  PIN dsadc_conv_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.406 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7864 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 10.838 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.7312 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.718 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8032 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M5  ;
    ANTENNAMAXAREACAR 221.67 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 979.965 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.76322 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 998.030000 445.480000 998.130000 446.000000 ;
    END
  END dsadc_conv_done
  PIN dsadc_en
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.112 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 4.578 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1872 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1042.800000 445.480000 1042.900000 446.000000 ;
    END
  END dsadc_en
  PIN dsadc_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.94 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0934 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 33.144 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.6344 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1027.510000 445.480000 1027.610000 446.000000 ;
    END
  END dsadc_clk
  PIN dsadc_switch[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5095 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2418 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.798 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5552 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 4.902 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6128 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1025.875000 445.480000 1025.975000 446.000000 ;
    END
  END dsadc_switch[2]
  PIN dsadc_switch[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.284 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2496 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.002 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4528 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1026.420000 445.480000 1026.520000 446.000000 ;
    END
  END dsadc_switch[1]
  PIN dsadc_switch[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.9205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0942 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1026.965000 445.480000 1027.065000 446.000000 ;
    END
  END dsadc_switch[0]
  PIN dac_en_pot
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0445 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1958 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.0676 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 1.058 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6992 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 5.362 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 23.6368 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1042.255000 445.480000 1042.355000 446.000000 ;
    END
  END dac_en_pot
  PIN adc_ext_in
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1012.250000 445.480000 1012.350000 446.000000 ;
    END
  END adc_ext_in
  PIN atp_en
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9445 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1558 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 6.466 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.4944 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1010.615000 445.480000 1010.715000 446.000000 ;
    END
  END atp_en
  PIN atp_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.301 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3684 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.958 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6592 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1011.160000 445.480000 1011.260000 446.000000 ;
    END
  END atp_sel
  PIN adc_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0295 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1298 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 4.718 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8032 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1011.705000 445.480000 1011.805000 446.000000 ;
    END
  END adc_sel
  PIN saradc_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.291 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2804 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 874.605000 445.480000 874.705000 446.000000 ;
    END
  END saradc_clk
  PIN saradc_rdy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.571 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5124 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.3315 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9466 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 12.398 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 54.5952 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M5  ;
    ANTENNAMAXAREACAR 567.011 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 2498.6 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.95203 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 874.205000 445.480000 874.305000 446.000000 ;
    END
  END saradc_rdy
  PIN saradc_rst
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.265 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.21 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 873.805000 445.480000 873.905000 446.000000 ;
    END
  END saradc_rst
  PIN saradc_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3625 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.595 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 10.798 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.5552 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 404.566 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1781.88 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 873.405000 445.480000 873.505000 446.000000 ;
    END
  END saradc_data[9]
  PIN saradc_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.247 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0868 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 10.9335 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.1514 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 436.454 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1898.61 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 873.005000 445.480000 873.105000 446.000000 ;
    END
  END saradc_data[8]
  PIN saradc_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6515 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8666 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 6.542 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.8288 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.526 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M4  ;
    ANTENNAMAXAREACAR 225.83 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 992.59 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.84502 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 872.605000 445.480000 872.705000 446.000000 ;
    END
  END saradc_data[7]
  PIN saradc_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.231 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0164 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.266 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2144 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 13.042 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 57.4288 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M5  ;
    ANTENNAMAXAREACAR 578.672 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 2549.37 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.58303 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 872.205000 445.480000 872.305000 446.000000 ;
    END
  END saradc_data[6]
  PIN saradc_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7025 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.091 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 13.778 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.6672 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.518 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3232 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M4  ;
    ANTENNAMAXAREACAR 30.5535 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 136.295 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 871.805000 445.480000 871.905000 446.000000 ;
    END
  END saradc_data[5]
  PIN saradc_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8665 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8126 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 8.238 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.2912 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.706 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1504 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 5.218 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 23.0032 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M5  ;
    ANTENNAMAXAREACAR 246.199 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 1086.49 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.21402 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 871.405000 445.480000 871.505000 446.000000 ;
    END
  END saradc_data[4]
  PIN saradc_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.411 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8084 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 8.5575 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.697 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M3  ;
    ANTENNAMAXAREACAR 374.414 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1642.15 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.63265 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 871.005000 445.480000 871.105000 446.000000 ;
    END
  END saradc_data[3]
  PIN saradc_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.371 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6324 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.8335 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7114 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.246 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M4  ;
    ANTENNAMAXAREACAR 497.727 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 2139.04 LAYER M4  ;
    ANTENNAMAXCUTCAR 2.21402 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 870.605000 445.480000 870.705000 446.000000 ;
    END
  END saradc_data[2]
  PIN saradc_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2465 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0846 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 9.302 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.9728 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M3  ;
    ANTENNAMAXAREACAR 386.245 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1701.44 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.22449 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 870.205000 445.480000 870.305000 446.000000 ;
    END
  END saradc_data[1]
  PIN saradc_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8435 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7114 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 6.038 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.6112 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.526 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 7.478 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 32.9472 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M5  ;
    ANTENNAMAXAREACAR 313.506 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 1382.38 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.84502 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 869.805000 445.480000 869.905000 446.000000 ;
    END
  END saradc_data[0]
  PIN a0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[31]
  PIN a0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[30]
  PIN a0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[29]
  PIN a0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[28]
  PIN a0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[27]
  PIN a0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[26]
  PIN a0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[25]
  PIN a0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[24]
  PIN a0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[23]
  PIN a0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[22]
  PIN a0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[21]
  PIN a0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[20]
  PIN a0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[19]
  PIN a0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[18]
  PIN a0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[17]
  PIN a0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[16]
  PIN a0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[15]
  PIN a0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[14]
  PIN a0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[13]
  PIN a0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[12]
  PIN a0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[11]
  PIN a0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[10]
  PIN a0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[9]
  PIN a0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[8]
  PIN a0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[7]
  PIN a0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[6]
  PIN a0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[5]
  PIN a0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[4]
  PIN a0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[3]
  PIN a0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[2]
  PIN a0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[1]
  PIN a0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[0]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M7 ;
        RECT 51.000000 0.000000 56.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 51.000000 681.000000 56.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 101.000000 0.000000 106.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 101.000000 681.000000 106.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 151.000000 0.000000 156.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 151.000000 681.000000 156.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 201.000000 0.000000 206.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 201.000000 681.000000 206.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 251.000000 0.000000 256.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 251.000000 681.000000 256.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 301.000000 0.000000 306.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 301.000000 681.000000 306.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 351.000000 0.000000 356.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 351.000000 681.000000 356.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 401.000000 0.000000 406.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 401.000000 501.000000 406.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 401.000000 656.000000 406.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 401.000000 681.000000 406.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 451.000000 0.000000 456.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 451.000000 501.000000 456.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 451.000000 656.000000 456.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 451.000000 681.000000 456.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 501.000000 0.000000 506.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 501.000000 501.000000 506.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 501.000000 656.000000 506.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 501.000000 681.000000 506.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 551.000000 0.000000 556.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 551.000000 501.000000 556.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 551.000000 656.000000 556.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 551.000000 681.000000 556.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 601.000000 0.000000 606.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 601.000000 501.000000 606.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 601.000000 656.000000 606.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 601.000000 681.000000 606.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 651.000000 0.000000 656.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 651.000000 501.000000 656.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 651.000000 656.000000 656.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 651.000000 681.000000 656.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 701.000000 0.000000 706.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 701.000000 501.000000 706.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 751.000000 0.000000 756.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 751.000000 441.000000 756.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 801.000000 0.000000 806.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 801.000000 441.000000 806.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 851.000000 0.000000 856.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 851.000000 441.000000 856.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 901.000000 0.000000 906.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 901.000000 441.000000 906.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 951.000000 0.000000 956.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 951.000000 441.000000 956.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1001.000000 0.000000 1006.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1001.000000 441.000000 1006.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1051.000000 0.000000 1056.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1051.000000 441.000000 1056.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1101.000000 0.000000 1106.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1101.000000 441.000000 1106.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1151.000000 0.000000 1156.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1151.000000 681.000000 1156.000000 686.000000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER M2 ;
        RECT 4.000000 5.910000 14.000000 6.090000 ;
        RECT 51.000000 5.910000 56.000000 6.090000 ;
        RECT 51.000000 1.910000 56.000000 2.090000 ;
        RECT 101.000000 1.910000 106.000000 2.090000 ;
        RECT 101.000000 5.910000 106.000000 6.090000 ;
        RECT 151.000000 1.910000 156.000000 2.090000 ;
        RECT 151.000000 5.910000 156.000000 6.090000 ;
        RECT 201.000000 1.910000 206.000000 2.090000 ;
        RECT 201.000000 5.910000 206.000000 6.090000 ;
        RECT 251.000000 1.910000 256.000000 2.090000 ;
        RECT 251.000000 5.910000 256.000000 6.090000 ;
        RECT 301.000000 1.910000 306.000000 2.090000 ;
        RECT 301.000000 5.910000 306.000000 6.090000 ;
        RECT 351.000000 1.910000 356.000000 2.090000 ;
        RECT 351.000000 5.910000 356.000000 6.090000 ;
        RECT 401.000000 1.910000 406.000000 2.090000 ;
        RECT 401.000000 5.910000 406.000000 6.090000 ;
        RECT 451.000000 1.910000 456.000000 2.090000 ;
        RECT 451.000000 5.910000 456.000000 6.090000 ;
        RECT 501.000000 1.910000 506.000000 2.090000 ;
        RECT 501.000000 5.910000 506.000000 6.090000 ;
        RECT 551.000000 1.910000 556.000000 2.090000 ;
        RECT 551.000000 5.910000 556.000000 6.090000 ;
        RECT 4.000000 265.910000 14.000000 266.090000 ;
        RECT 4.000000 261.910000 14.000000 262.090000 ;
        RECT 51.000000 265.910000 56.000000 266.090000 ;
        RECT 51.000000 261.910000 56.000000 262.090000 ;
        RECT 101.000000 265.910000 106.000000 266.090000 ;
        RECT 101.000000 261.910000 106.000000 262.090000 ;
        RECT 51.000000 305.910000 56.000000 306.090000 ;
        RECT 4.000000 305.910000 14.000000 306.090000 ;
        RECT 4.000000 285.910000 14.000000 286.090000 ;
        RECT 4.000000 281.910000 14.000000 282.090000 ;
        RECT 4.000000 269.910000 14.000000 270.090000 ;
        RECT 4.000000 273.910000 14.000000 274.090000 ;
        RECT 4.000000 277.910000 14.000000 278.090000 ;
        RECT 4.000000 289.910000 14.000000 290.090000 ;
        RECT 4.000000 293.910000 14.000000 294.090000 ;
        RECT 4.000000 297.910000 14.000000 298.090000 ;
        RECT 4.000000 301.910000 14.000000 302.090000 ;
        RECT 51.000000 269.910000 56.000000 270.090000 ;
        RECT 51.000000 273.910000 56.000000 274.090000 ;
        RECT 51.000000 277.910000 56.000000 278.090000 ;
        RECT 51.000000 281.910000 56.000000 282.090000 ;
        RECT 51.000000 285.910000 56.000000 286.090000 ;
        RECT 51.000000 301.910000 56.000000 302.090000 ;
        RECT 51.000000 297.910000 56.000000 298.090000 ;
        RECT 51.000000 293.910000 56.000000 294.090000 ;
        RECT 51.000000 289.910000 56.000000 290.090000 ;
        RECT 4.000000 321.910000 14.000000 322.090000 ;
        RECT 4.000000 317.910000 14.000000 318.090000 ;
        RECT 4.000000 309.910000 14.000000 310.090000 ;
        RECT 4.000000 313.910000 14.000000 314.090000 ;
        RECT 4.000000 325.910000 14.000000 326.090000 ;
        RECT 4.000000 329.910000 14.000000 330.090000 ;
        RECT 4.000000 333.910000 14.000000 334.090000 ;
        RECT 4.000000 337.910000 14.000000 338.090000 ;
        RECT 4.000000 341.910000 14.000000 342.090000 ;
        RECT 51.000000 313.910000 56.000000 314.090000 ;
        RECT 51.000000 309.910000 56.000000 310.090000 ;
        RECT 51.000000 317.910000 56.000000 318.090000 ;
        RECT 51.000000 321.910000 56.000000 322.090000 ;
        RECT 51.000000 341.910000 56.000000 342.090000 ;
        RECT 51.000000 337.910000 56.000000 338.090000 ;
        RECT 51.000000 333.910000 56.000000 334.090000 ;
        RECT 51.000000 329.910000 56.000000 330.090000 ;
        RECT 51.000000 325.910000 56.000000 326.090000 ;
        RECT 101.000000 305.910000 106.000000 306.090000 ;
        RECT 101.000000 285.910000 106.000000 286.090000 ;
        RECT 101.000000 269.910000 106.000000 270.090000 ;
        RECT 101.000000 273.910000 106.000000 274.090000 ;
        RECT 101.000000 277.910000 106.000000 278.090000 ;
        RECT 101.000000 281.910000 106.000000 282.090000 ;
        RECT 101.000000 301.910000 106.000000 302.090000 ;
        RECT 101.000000 297.910000 106.000000 298.090000 ;
        RECT 101.000000 293.910000 106.000000 294.090000 ;
        RECT 101.000000 289.910000 106.000000 290.090000 ;
        RECT 101.000000 321.910000 106.000000 322.090000 ;
        RECT 101.000000 317.910000 106.000000 318.090000 ;
        RECT 101.000000 313.910000 106.000000 314.090000 ;
        RECT 101.000000 309.910000 106.000000 310.090000 ;
        RECT 101.000000 325.910000 106.000000 326.090000 ;
        RECT 101.000000 329.910000 106.000000 330.090000 ;
        RECT 101.000000 333.910000 106.000000 334.090000 ;
        RECT 101.000000 337.910000 106.000000 338.090000 ;
        RECT 101.000000 341.910000 106.000000 342.090000 ;
        RECT 151.000000 261.910000 156.000000 262.090000 ;
        RECT 151.000000 265.910000 156.000000 266.090000 ;
        RECT 201.000000 265.910000 206.000000 266.090000 ;
        RECT 201.000000 261.910000 206.000000 262.090000 ;
        RECT 251.000000 265.910000 256.000000 266.090000 ;
        RECT 251.000000 261.910000 256.000000 262.090000 ;
        RECT 201.000000 305.910000 206.000000 306.090000 ;
        RECT 151.000000 305.910000 156.000000 306.090000 ;
        RECT 151.000000 269.910000 156.000000 270.090000 ;
        RECT 151.000000 273.910000 156.000000 274.090000 ;
        RECT 151.000000 277.910000 156.000000 278.090000 ;
        RECT 151.000000 281.910000 156.000000 282.090000 ;
        RECT 151.000000 285.910000 156.000000 286.090000 ;
        RECT 151.000000 289.910000 156.000000 290.090000 ;
        RECT 151.000000 293.910000 156.000000 294.090000 ;
        RECT 151.000000 301.910000 156.000000 302.090000 ;
        RECT 151.000000 297.910000 156.000000 298.090000 ;
        RECT 201.000000 269.910000 206.000000 270.090000 ;
        RECT 201.000000 273.910000 206.000000 274.090000 ;
        RECT 201.000000 277.910000 206.000000 278.090000 ;
        RECT 201.000000 281.910000 206.000000 282.090000 ;
        RECT 201.000000 285.910000 206.000000 286.090000 ;
        RECT 201.000000 301.910000 206.000000 302.090000 ;
        RECT 201.000000 297.910000 206.000000 298.090000 ;
        RECT 201.000000 293.910000 206.000000 294.090000 ;
        RECT 201.000000 289.910000 206.000000 290.090000 ;
        RECT 151.000000 313.910000 156.000000 314.090000 ;
        RECT 151.000000 309.910000 156.000000 310.090000 ;
        RECT 151.000000 321.910000 156.000000 322.090000 ;
        RECT 151.000000 317.910000 156.000000 318.090000 ;
        RECT 151.000000 329.910000 156.000000 330.090000 ;
        RECT 151.000000 325.910000 156.000000 326.090000 ;
        RECT 151.000000 333.910000 156.000000 334.090000 ;
        RECT 151.000000 337.910000 156.000000 338.090000 ;
        RECT 151.000000 341.910000 156.000000 342.090000 ;
        RECT 201.000000 313.910000 206.000000 314.090000 ;
        RECT 201.000000 309.910000 206.000000 310.090000 ;
        RECT 201.000000 317.910000 206.000000 318.090000 ;
        RECT 201.000000 321.910000 206.000000 322.090000 ;
        RECT 201.000000 341.910000 206.000000 342.090000 ;
        RECT 201.000000 337.910000 206.000000 338.090000 ;
        RECT 201.000000 333.910000 206.000000 334.090000 ;
        RECT 201.000000 329.910000 206.000000 330.090000 ;
        RECT 201.000000 325.910000 206.000000 326.090000 ;
        RECT 251.000000 305.910000 256.000000 306.090000 ;
        RECT 251.000000 269.910000 256.000000 270.090000 ;
        RECT 251.000000 273.910000 256.000000 274.090000 ;
        RECT 251.000000 277.910000 256.000000 278.090000 ;
        RECT 251.000000 281.910000 256.000000 282.090000 ;
        RECT 251.000000 285.910000 256.000000 286.090000 ;
        RECT 251.000000 293.910000 256.000000 294.090000 ;
        RECT 251.000000 289.910000 256.000000 290.090000 ;
        RECT 251.000000 301.910000 256.000000 302.090000 ;
        RECT 251.000000 297.910000 256.000000 298.090000 ;
        RECT 251.000000 309.910000 256.000000 310.090000 ;
        RECT 251.000000 313.910000 256.000000 314.090000 ;
        RECT 251.000000 321.910000 256.000000 322.090000 ;
        RECT 251.000000 317.910000 256.000000 318.090000 ;
        RECT 251.000000 329.910000 256.000000 330.090000 ;
        RECT 251.000000 325.910000 256.000000 326.090000 ;
        RECT 251.000000 333.910000 256.000000 334.090000 ;
        RECT 251.000000 337.910000 256.000000 338.090000 ;
        RECT 251.000000 341.910000 256.000000 342.090000 ;
        RECT 301.000000 265.910000 306.000000 266.090000 ;
        RECT 301.000000 261.910000 306.000000 262.090000 ;
        RECT 351.000000 265.910000 356.000000 266.090000 ;
        RECT 351.000000 261.910000 356.000000 262.090000 ;
        RECT 401.000000 265.910000 406.000000 266.090000 ;
        RECT 401.000000 261.910000 406.000000 262.090000 ;
        RECT 351.000000 305.910000 356.000000 306.090000 ;
        RECT 301.000000 305.910000 306.000000 306.090000 ;
        RECT 301.000000 277.910000 306.000000 278.090000 ;
        RECT 301.000000 269.910000 306.000000 270.090000 ;
        RECT 301.000000 273.910000 306.000000 274.090000 ;
        RECT 301.000000 281.910000 306.000000 282.090000 ;
        RECT 301.000000 285.910000 306.000000 286.090000 ;
        RECT 301.000000 293.910000 306.000000 294.090000 ;
        RECT 301.000000 289.910000 306.000000 290.090000 ;
        RECT 301.000000 301.910000 306.000000 302.090000 ;
        RECT 301.000000 297.910000 306.000000 298.090000 ;
        RECT 351.000000 269.910000 356.000000 270.090000 ;
        RECT 351.000000 273.910000 356.000000 274.090000 ;
        RECT 351.000000 277.910000 356.000000 278.090000 ;
        RECT 351.000000 281.910000 356.000000 282.090000 ;
        RECT 351.000000 285.910000 356.000000 286.090000 ;
        RECT 351.000000 301.910000 356.000000 302.090000 ;
        RECT 351.000000 297.910000 356.000000 298.090000 ;
        RECT 351.000000 293.910000 356.000000 294.090000 ;
        RECT 351.000000 289.910000 356.000000 290.090000 ;
        RECT 301.000000 313.910000 306.000000 314.090000 ;
        RECT 301.000000 309.910000 306.000000 310.090000 ;
        RECT 301.000000 317.910000 306.000000 318.090000 ;
        RECT 301.000000 321.910000 306.000000 322.090000 ;
        RECT 301.000000 329.910000 306.000000 330.090000 ;
        RECT 301.000000 325.910000 306.000000 326.090000 ;
        RECT 301.000000 341.910000 306.000000 342.090000 ;
        RECT 301.000000 337.910000 306.000000 338.090000 ;
        RECT 301.000000 333.910000 306.000000 334.090000 ;
        RECT 351.000000 313.910000 356.000000 314.090000 ;
        RECT 351.000000 309.910000 356.000000 310.090000 ;
        RECT 351.000000 317.910000 356.000000 318.090000 ;
        RECT 351.000000 321.910000 356.000000 322.090000 ;
        RECT 351.000000 341.910000 356.000000 342.090000 ;
        RECT 351.000000 337.910000 356.000000 338.090000 ;
        RECT 351.000000 333.910000 356.000000 334.090000 ;
        RECT 351.000000 329.910000 356.000000 330.090000 ;
        RECT 351.000000 325.910000 356.000000 326.090000 ;
        RECT 401.000000 305.910000 406.000000 306.090000 ;
        RECT 401.000000 269.910000 406.000000 270.090000 ;
        RECT 401.000000 273.910000 406.000000 274.090000 ;
        RECT 401.000000 277.910000 406.000000 278.090000 ;
        RECT 401.000000 285.910000 406.000000 286.090000 ;
        RECT 401.000000 281.910000 406.000000 282.090000 ;
        RECT 401.000000 293.910000 406.000000 294.090000 ;
        RECT 401.000000 289.910000 406.000000 290.090000 ;
        RECT 401.000000 297.910000 406.000000 298.090000 ;
        RECT 401.000000 301.910000 406.000000 302.090000 ;
        RECT 401.000000 309.910000 406.000000 310.090000 ;
        RECT 401.000000 313.910000 406.000000 314.090000 ;
        RECT 401.000000 317.910000 406.000000 318.090000 ;
        RECT 401.000000 321.910000 406.000000 322.090000 ;
        RECT 401.000000 325.910000 406.000000 326.090000 ;
        RECT 401.000000 329.910000 406.000000 330.090000 ;
        RECT 401.000000 333.910000 406.000000 334.090000 ;
        RECT 401.000000 337.910000 406.000000 338.090000 ;
        RECT 401.000000 341.910000 406.000000 342.090000 ;
        RECT 451.000000 261.910000 456.000000 262.090000 ;
        RECT 451.000000 265.910000 456.000000 266.090000 ;
        RECT 501.000000 261.910000 506.000000 262.090000 ;
        RECT 501.000000 265.910000 506.000000 266.090000 ;
        RECT 551.000000 265.910000 556.000000 266.090000 ;
        RECT 551.000000 261.910000 556.000000 262.090000 ;
        RECT 501.000000 305.910000 506.000000 306.090000 ;
        RECT 451.000000 273.910000 456.000000 274.090000 ;
        RECT 451.000000 269.910000 456.000000 270.090000 ;
        RECT 451.000000 277.910000 456.000000 278.090000 ;
        RECT 451.000000 285.910000 456.000000 286.090000 ;
        RECT 451.000000 281.910000 456.000000 282.090000 ;
        RECT 451.000000 293.910000 456.000000 294.090000 ;
        RECT 451.000000 289.910000 456.000000 290.090000 ;
        RECT 451.000000 297.910000 456.000000 298.090000 ;
        RECT 501.000000 277.910000 506.000000 278.090000 ;
        RECT 501.000000 273.910000 506.000000 274.090000 ;
        RECT 501.000000 269.910000 506.000000 270.090000 ;
        RECT 501.000000 281.910000 506.000000 282.090000 ;
        RECT 501.000000 285.910000 506.000000 286.090000 ;
        RECT 501.000000 289.910000 506.000000 290.090000 ;
        RECT 501.000000 293.910000 506.000000 294.090000 ;
        RECT 501.000000 301.910000 506.000000 302.090000 ;
        RECT 501.000000 297.910000 506.000000 298.090000 ;
        RECT 451.000000 321.910000 456.000000 322.090000 ;
        RECT 451.000000 333.910000 456.000000 334.090000 ;
        RECT 451.000000 329.910000 456.000000 330.090000 ;
        RECT 451.000000 325.910000 456.000000 326.090000 ;
        RECT 451.000000 337.910000 456.000000 338.090000 ;
        RECT 451.000000 341.910000 456.000000 342.090000 ;
        RECT 501.000000 313.910000 506.000000 314.090000 ;
        RECT 501.000000 309.910000 506.000000 310.090000 ;
        RECT 501.000000 317.910000 506.000000 318.090000 ;
        RECT 501.000000 321.910000 506.000000 322.090000 ;
        RECT 501.000000 329.910000 506.000000 330.090000 ;
        RECT 501.000000 325.910000 506.000000 326.090000 ;
        RECT 501.000000 333.910000 506.000000 334.090000 ;
        RECT 501.000000 337.910000 506.000000 338.090000 ;
        RECT 501.000000 341.910000 506.000000 342.090000 ;
        RECT 551.000000 305.910000 556.000000 306.090000 ;
        RECT 551.000000 281.910000 556.000000 282.090000 ;
        RECT 551.000000 277.910000 556.000000 278.090000 ;
        RECT 551.000000 273.910000 556.000000 274.090000 ;
        RECT 551.000000 269.910000 556.000000 270.090000 ;
        RECT 551.000000 285.910000 556.000000 286.090000 ;
        RECT 551.000000 301.910000 556.000000 302.090000 ;
        RECT 551.000000 297.910000 556.000000 298.090000 ;
        RECT 551.000000 293.910000 556.000000 294.090000 ;
        RECT 551.000000 289.910000 556.000000 290.090000 ;
        RECT 551.000000 313.910000 556.000000 314.090000 ;
        RECT 551.000000 309.910000 556.000000 310.090000 ;
        RECT 551.000000 321.910000 556.000000 322.090000 ;
        RECT 551.000000 317.910000 556.000000 318.090000 ;
        RECT 551.000000 325.910000 556.000000 326.090000 ;
        RECT 551.000000 329.910000 556.000000 330.090000 ;
        RECT 551.000000 333.910000 556.000000 334.090000 ;
        RECT 551.000000 337.910000 556.000000 338.090000 ;
        RECT 551.000000 341.910000 556.000000 342.090000 ;
        RECT 601.000000 1.910000 606.000000 2.090000 ;
        RECT 601.000000 5.910000 606.000000 6.090000 ;
        RECT 651.000000 1.910000 656.000000 2.090000 ;
        RECT 651.000000 5.910000 656.000000 6.090000 ;
        RECT 701.000000 1.910000 706.000000 2.090000 ;
        RECT 701.000000 5.910000 706.000000 6.090000 ;
        RECT 751.000000 1.910000 756.000000 2.090000 ;
        RECT 751.000000 5.910000 756.000000 6.090000 ;
        RECT 801.000000 1.910000 806.000000 2.090000 ;
        RECT 801.000000 5.910000 806.000000 6.090000 ;
        RECT 851.000000 1.910000 856.000000 2.090000 ;
        RECT 851.000000 5.910000 856.000000 6.090000 ;
        RECT 901.000000 1.910000 906.000000 2.090000 ;
        RECT 901.000000 5.910000 906.000000 6.090000 ;
        RECT 951.000000 1.910000 956.000000 2.090000 ;
        RECT 951.000000 5.910000 956.000000 6.090000 ;
        RECT 1001.000000 1.910000 1006.000000 2.090000 ;
        RECT 1001.000000 5.910000 1006.000000 6.090000 ;
        RECT 1051.000000 1.910000 1056.000000 2.090000 ;
        RECT 1051.000000 5.910000 1056.000000 6.090000 ;
        RECT 1101.000000 1.910000 1106.000000 2.090000 ;
        RECT 1101.000000 5.910000 1106.000000 6.090000 ;
        RECT 1151.000000 5.910000 1156.000000 6.090000 ;
        RECT 1172.000000 5.910000 1182.000000 6.090000 ;
        RECT 1151.000000 1.910000 1156.000000 2.090000 ;
        RECT 1172.000000 17.910000 1182.000000 18.090000 ;
        RECT 1172.000000 13.910000 1182.000000 14.090000 ;
        RECT 1172.000000 9.910000 1182.000000 10.090000 ;
        RECT 1172.000000 21.910000 1182.000000 22.090000 ;
        RECT 1172.000000 25.910000 1182.000000 26.090000 ;
        RECT 1172.000000 33.910000 1182.000000 34.090000 ;
        RECT 1172.000000 29.910000 1182.000000 30.090000 ;
        RECT 1172.000000 41.910000 1182.000000 42.090000 ;
        RECT 1172.000000 37.910000 1182.000000 38.090000 ;
        RECT 1172.000000 45.910000 1182.000000 46.090000 ;
        RECT 601.000000 265.910000 606.000000 266.090000 ;
        RECT 601.000000 261.910000 606.000000 262.090000 ;
        RECT 651.000000 261.910000 656.000000 262.090000 ;
        RECT 651.000000 265.910000 656.000000 266.090000 ;
        RECT 701.000000 265.910000 706.000000 266.090000 ;
        RECT 701.000000 261.910000 706.000000 262.090000 ;
        RECT 601.000000 305.910000 606.000000 306.090000 ;
        RECT 651.000000 305.910000 656.000000 306.090000 ;
        RECT 601.000000 269.910000 606.000000 270.090000 ;
        RECT 601.000000 273.910000 606.000000 274.090000 ;
        RECT 601.000000 277.910000 606.000000 278.090000 ;
        RECT 601.000000 281.910000 606.000000 282.090000 ;
        RECT 601.000000 285.910000 606.000000 286.090000 ;
        RECT 601.000000 293.910000 606.000000 294.090000 ;
        RECT 601.000000 289.910000 606.000000 290.090000 ;
        RECT 601.000000 301.910000 606.000000 302.090000 ;
        RECT 601.000000 297.910000 606.000000 298.090000 ;
        RECT 651.000000 269.910000 656.000000 270.090000 ;
        RECT 651.000000 273.910000 656.000000 274.090000 ;
        RECT 651.000000 277.910000 656.000000 278.090000 ;
        RECT 651.000000 281.910000 656.000000 282.090000 ;
        RECT 651.000000 285.910000 656.000000 286.090000 ;
        RECT 651.000000 289.910000 656.000000 290.090000 ;
        RECT 651.000000 293.910000 656.000000 294.090000 ;
        RECT 651.000000 297.910000 656.000000 298.090000 ;
        RECT 651.000000 301.910000 656.000000 302.090000 ;
        RECT 601.000000 313.910000 606.000000 314.090000 ;
        RECT 601.000000 309.910000 606.000000 310.090000 ;
        RECT 601.000000 317.910000 606.000000 318.090000 ;
        RECT 601.000000 321.910000 606.000000 322.090000 ;
        RECT 601.000000 325.910000 606.000000 326.090000 ;
        RECT 601.000000 329.910000 606.000000 330.090000 ;
        RECT 601.000000 333.910000 606.000000 334.090000 ;
        RECT 601.000000 337.910000 606.000000 338.090000 ;
        RECT 601.000000 341.910000 606.000000 342.090000 ;
        RECT 651.000000 313.910000 656.000000 314.090000 ;
        RECT 651.000000 309.910000 656.000000 310.090000 ;
        RECT 651.000000 321.910000 656.000000 322.090000 ;
        RECT 651.000000 317.910000 656.000000 318.090000 ;
        RECT 651.000000 329.910000 656.000000 330.090000 ;
        RECT 651.000000 325.910000 656.000000 326.090000 ;
        RECT 651.000000 333.910000 656.000000 334.090000 ;
        RECT 651.000000 337.910000 656.000000 338.090000 ;
        RECT 651.000000 341.910000 656.000000 342.090000 ;
        RECT 701.000000 305.910000 706.000000 306.090000 ;
        RECT 701.000000 281.910000 706.000000 282.090000 ;
        RECT 701.000000 277.910000 706.000000 278.090000 ;
        RECT 701.000000 273.910000 706.000000 274.090000 ;
        RECT 701.000000 269.910000 706.000000 270.090000 ;
        RECT 701.000000 285.910000 706.000000 286.090000 ;
        RECT 701.000000 301.910000 706.000000 302.090000 ;
        RECT 701.000000 297.910000 706.000000 298.090000 ;
        RECT 701.000000 293.910000 706.000000 294.090000 ;
        RECT 701.000000 289.910000 706.000000 290.090000 ;
        RECT 701.000000 309.910000 706.000000 310.090000 ;
        RECT 701.000000 313.910000 706.000000 314.090000 ;
        RECT 701.000000 317.910000 706.000000 318.090000 ;
        RECT 701.000000 321.910000 706.000000 322.090000 ;
        RECT 701.000000 325.910000 706.000000 326.090000 ;
        RECT 701.000000 329.910000 706.000000 330.090000 ;
        RECT 701.000000 333.910000 706.000000 334.090000 ;
        RECT 701.000000 337.910000 706.000000 338.090000 ;
        RECT 701.000000 341.910000 706.000000 342.090000 ;
        RECT 751.000000 261.910000 756.000000 262.090000 ;
        RECT 751.000000 265.910000 756.000000 266.090000 ;
        RECT 801.000000 261.910000 806.000000 262.090000 ;
        RECT 801.000000 265.910000 806.000000 266.090000 ;
        RECT 851.000000 265.910000 856.000000 266.090000 ;
        RECT 851.000000 261.910000 856.000000 262.090000 ;
        RECT 801.000000 305.910000 806.000000 306.090000 ;
        RECT 751.000000 305.910000 756.000000 306.090000 ;
        RECT 751.000000 285.910000 756.000000 286.090000 ;
        RECT 751.000000 281.910000 756.000000 282.090000 ;
        RECT 751.000000 269.910000 756.000000 270.090000 ;
        RECT 751.000000 273.910000 756.000000 274.090000 ;
        RECT 751.000000 277.910000 756.000000 278.090000 ;
        RECT 751.000000 289.910000 756.000000 290.090000 ;
        RECT 751.000000 293.910000 756.000000 294.090000 ;
        RECT 751.000000 297.910000 756.000000 298.090000 ;
        RECT 751.000000 301.910000 756.000000 302.090000 ;
        RECT 801.000000 277.910000 806.000000 278.090000 ;
        RECT 801.000000 273.910000 806.000000 274.090000 ;
        RECT 801.000000 269.910000 806.000000 270.090000 ;
        RECT 801.000000 281.910000 806.000000 282.090000 ;
        RECT 801.000000 285.910000 806.000000 286.090000 ;
        RECT 801.000000 289.910000 806.000000 290.090000 ;
        RECT 801.000000 293.910000 806.000000 294.090000 ;
        RECT 801.000000 301.910000 806.000000 302.090000 ;
        RECT 801.000000 297.910000 806.000000 298.090000 ;
        RECT 751.000000 321.910000 756.000000 322.090000 ;
        RECT 751.000000 317.910000 756.000000 318.090000 ;
        RECT 751.000000 309.910000 756.000000 310.090000 ;
        RECT 751.000000 313.910000 756.000000 314.090000 ;
        RECT 751.000000 329.910000 756.000000 330.090000 ;
        RECT 751.000000 325.910000 756.000000 326.090000 ;
        RECT 751.000000 341.910000 756.000000 342.090000 ;
        RECT 751.000000 337.910000 756.000000 338.090000 ;
        RECT 751.000000 333.910000 756.000000 334.090000 ;
        RECT 801.000000 309.910000 806.000000 310.090000 ;
        RECT 801.000000 313.910000 806.000000 314.090000 ;
        RECT 801.000000 321.910000 806.000000 322.090000 ;
        RECT 801.000000 317.910000 806.000000 318.090000 ;
        RECT 801.000000 325.910000 806.000000 326.090000 ;
        RECT 801.000000 329.910000 806.000000 330.090000 ;
        RECT 801.000000 337.910000 806.000000 338.090000 ;
        RECT 801.000000 333.910000 806.000000 334.090000 ;
        RECT 801.000000 341.910000 806.000000 342.090000 ;
        RECT 851.000000 305.910000 856.000000 306.090000 ;
        RECT 851.000000 281.910000 856.000000 282.090000 ;
        RECT 851.000000 277.910000 856.000000 278.090000 ;
        RECT 851.000000 273.910000 856.000000 274.090000 ;
        RECT 851.000000 269.910000 856.000000 270.090000 ;
        RECT 851.000000 285.910000 856.000000 286.090000 ;
        RECT 851.000000 301.910000 856.000000 302.090000 ;
        RECT 851.000000 297.910000 856.000000 298.090000 ;
        RECT 851.000000 293.910000 856.000000 294.090000 ;
        RECT 851.000000 289.910000 856.000000 290.090000 ;
        RECT 851.000000 309.910000 856.000000 310.090000 ;
        RECT 851.000000 313.910000 856.000000 314.090000 ;
        RECT 851.000000 317.910000 856.000000 318.090000 ;
        RECT 851.000000 321.910000 856.000000 322.090000 ;
        RECT 851.000000 325.910000 856.000000 326.090000 ;
        RECT 851.000000 329.910000 856.000000 330.090000 ;
        RECT 851.000000 333.910000 856.000000 334.090000 ;
        RECT 851.000000 337.910000 856.000000 338.090000 ;
        RECT 851.000000 341.910000 856.000000 342.090000 ;
        RECT 1172.000000 61.910000 1182.000000 62.090000 ;
        RECT 1172.000000 57.910000 1182.000000 58.090000 ;
        RECT 1172.000000 53.910000 1182.000000 54.090000 ;
        RECT 1172.000000 49.910000 1182.000000 50.090000 ;
        RECT 1172.000000 73.910000 1182.000000 74.090000 ;
        RECT 1172.000000 69.910000 1182.000000 70.090000 ;
        RECT 1172.000000 65.910000 1182.000000 66.090000 ;
        RECT 1172.000000 77.910000 1182.000000 78.090000 ;
        RECT 1172.000000 81.910000 1182.000000 82.090000 ;
        RECT 1172.000000 85.910000 1182.000000 86.090000 ;
        RECT 1172.000000 89.910000 1182.000000 90.090000 ;
        RECT 1172.000000 97.910000 1182.000000 98.090000 ;
        RECT 1172.000000 93.910000 1182.000000 94.090000 ;
        RECT 1172.000000 101.910000 1182.000000 102.090000 ;
        RECT 1172.000000 117.910000 1182.000000 118.090000 ;
        RECT 1172.000000 113.910000 1182.000000 114.090000 ;
        RECT 1172.000000 105.910000 1182.000000 106.090000 ;
        RECT 1172.000000 109.910000 1182.000000 110.090000 ;
        RECT 1151.000000 133.910000 1156.000000 134.090000 ;
        RECT 1172.000000 125.910000 1182.000000 126.090000 ;
        RECT 1172.000000 121.910000 1182.000000 122.090000 ;
        RECT 1172.000000 129.910000 1182.000000 130.090000 ;
        RECT 1172.000000 133.910000 1182.000000 134.090000 ;
        RECT 1172.000000 137.910000 1182.000000 138.090000 ;
        RECT 1172.000000 141.910000 1182.000000 142.090000 ;
        RECT 1172.000000 145.910000 1182.000000 146.090000 ;
        RECT 1172.000000 149.910000 1182.000000 150.090000 ;
        RECT 1172.000000 153.910000 1182.000000 154.090000 ;
        RECT 1172.000000 165.910000 1182.000000 166.090000 ;
        RECT 1172.000000 161.910000 1182.000000 162.090000 ;
        RECT 1172.000000 157.910000 1182.000000 158.090000 ;
        RECT 1172.000000 169.910000 1182.000000 170.090000 ;
        RECT 1172.000000 173.910000 1182.000000 174.090000 ;
        RECT 1172.000000 177.910000 1182.000000 178.090000 ;
        RECT 1172.000000 181.910000 1182.000000 182.090000 ;
        RECT 1172.000000 185.910000 1182.000000 186.090000 ;
        RECT 1172.000000 189.910000 1182.000000 190.090000 ;
        RECT 1172.000000 193.910000 1182.000000 194.090000 ;
        RECT 901.000000 261.910000 906.000000 262.090000 ;
        RECT 901.000000 265.910000 906.000000 266.090000 ;
        RECT 951.000000 265.910000 956.000000 266.090000 ;
        RECT 951.000000 261.910000 956.000000 262.090000 ;
        RECT 1001.000000 261.910000 1006.000000 262.090000 ;
        RECT 1001.000000 265.910000 1006.000000 266.090000 ;
        RECT 951.000000 305.910000 956.000000 306.090000 ;
        RECT 901.000000 305.910000 906.000000 306.090000 ;
        RECT 901.000000 285.910000 906.000000 286.090000 ;
        RECT 901.000000 281.910000 906.000000 282.090000 ;
        RECT 901.000000 269.910000 906.000000 270.090000 ;
        RECT 901.000000 273.910000 906.000000 274.090000 ;
        RECT 901.000000 277.910000 906.000000 278.090000 ;
        RECT 901.000000 289.910000 906.000000 290.090000 ;
        RECT 901.000000 293.910000 906.000000 294.090000 ;
        RECT 901.000000 297.910000 906.000000 298.090000 ;
        RECT 901.000000 301.910000 906.000000 302.090000 ;
        RECT 951.000000 269.910000 956.000000 270.090000 ;
        RECT 951.000000 273.910000 956.000000 274.090000 ;
        RECT 951.000000 277.910000 956.000000 278.090000 ;
        RECT 951.000000 281.910000 956.000000 282.090000 ;
        RECT 951.000000 285.910000 956.000000 286.090000 ;
        RECT 951.000000 301.910000 956.000000 302.090000 ;
        RECT 951.000000 297.910000 956.000000 298.090000 ;
        RECT 951.000000 293.910000 956.000000 294.090000 ;
        RECT 951.000000 289.910000 956.000000 290.090000 ;
        RECT 901.000000 321.910000 906.000000 322.090000 ;
        RECT 901.000000 309.910000 906.000000 310.090000 ;
        RECT 901.000000 313.910000 906.000000 314.090000 ;
        RECT 901.000000 317.910000 906.000000 318.090000 ;
        RECT 901.000000 325.910000 906.000000 326.090000 ;
        RECT 901.000000 329.910000 906.000000 330.090000 ;
        RECT 901.000000 333.910000 906.000000 334.090000 ;
        RECT 901.000000 337.910000 906.000000 338.090000 ;
        RECT 901.000000 341.910000 906.000000 342.090000 ;
        RECT 951.000000 313.910000 956.000000 314.090000 ;
        RECT 951.000000 309.910000 956.000000 310.090000 ;
        RECT 951.000000 317.910000 956.000000 318.090000 ;
        RECT 951.000000 321.910000 956.000000 322.090000 ;
        RECT 951.000000 325.910000 956.000000 326.090000 ;
        RECT 951.000000 329.910000 956.000000 330.090000 ;
        RECT 951.000000 333.910000 956.000000 334.090000 ;
        RECT 951.000000 337.910000 956.000000 338.090000 ;
        RECT 951.000000 341.910000 956.000000 342.090000 ;
        RECT 1001.000000 305.910000 1006.000000 306.090000 ;
        RECT 1001.000000 277.910000 1006.000000 278.090000 ;
        RECT 1001.000000 273.910000 1006.000000 274.090000 ;
        RECT 1001.000000 269.910000 1006.000000 270.090000 ;
        RECT 1001.000000 285.910000 1006.000000 286.090000 ;
        RECT 1001.000000 281.910000 1006.000000 282.090000 ;
        RECT 1001.000000 289.910000 1006.000000 290.090000 ;
        RECT 1001.000000 293.910000 1006.000000 294.090000 ;
        RECT 1001.000000 301.910000 1006.000000 302.090000 ;
        RECT 1001.000000 297.910000 1006.000000 298.090000 ;
        RECT 1001.000000 313.910000 1006.000000 314.090000 ;
        RECT 1001.000000 309.910000 1006.000000 310.090000 ;
        RECT 1001.000000 317.910000 1006.000000 318.090000 ;
        RECT 1001.000000 321.910000 1006.000000 322.090000 ;
        RECT 1001.000000 329.910000 1006.000000 330.090000 ;
        RECT 1001.000000 325.910000 1006.000000 326.090000 ;
        RECT 1001.000000 333.910000 1006.000000 334.090000 ;
        RECT 1001.000000 337.910000 1006.000000 338.090000 ;
        RECT 1001.000000 341.910000 1006.000000 342.090000 ;
        RECT 1051.000000 261.910000 1056.000000 262.090000 ;
        RECT 1051.000000 265.910000 1056.000000 266.090000 ;
        RECT 1101.000000 265.910000 1106.000000 266.090000 ;
        RECT 1101.000000 261.910000 1106.000000 262.090000 ;
        RECT 1172.000000 197.910000 1182.000000 198.090000 ;
        RECT 1172.000000 201.910000 1182.000000 202.090000 ;
        RECT 1172.000000 205.910000 1182.000000 206.090000 ;
        RECT 1172.000000 209.910000 1182.000000 210.090000 ;
        RECT 1172.000000 221.910000 1182.000000 222.090000 ;
        RECT 1172.000000 217.910000 1182.000000 218.090000 ;
        RECT 1172.000000 213.910000 1182.000000 214.090000 ;
        RECT 1172.000000 225.910000 1182.000000 226.090000 ;
        RECT 1172.000000 229.910000 1182.000000 230.090000 ;
        RECT 1172.000000 233.910000 1182.000000 234.090000 ;
        RECT 1172.000000 237.910000 1182.000000 238.090000 ;
        RECT 1172.000000 241.910000 1182.000000 242.090000 ;
        RECT 1172.000000 245.910000 1182.000000 246.090000 ;
        RECT 1172.000000 249.910000 1182.000000 250.090000 ;
        RECT 1151.000000 257.910000 1156.000000 258.090000 ;
        RECT 1151.000000 265.910000 1156.000000 266.090000 ;
        RECT 1151.000000 261.910000 1156.000000 262.090000 ;
        RECT 1172.000000 265.910000 1182.000000 266.090000 ;
        RECT 1172.000000 253.910000 1182.000000 254.090000 ;
        RECT 1172.000000 257.910000 1182.000000 258.090000 ;
        RECT 1172.000000 261.910000 1182.000000 262.090000 ;
        RECT 1101.000000 305.910000 1106.000000 306.090000 ;
        RECT 1051.000000 305.910000 1056.000000 306.090000 ;
        RECT 1051.000000 285.910000 1056.000000 286.090000 ;
        RECT 1051.000000 281.910000 1056.000000 282.090000 ;
        RECT 1051.000000 273.910000 1056.000000 274.090000 ;
        RECT 1051.000000 269.910000 1056.000000 270.090000 ;
        RECT 1051.000000 277.910000 1056.000000 278.090000 ;
        RECT 1051.000000 289.910000 1056.000000 290.090000 ;
        RECT 1051.000000 293.910000 1056.000000 294.090000 ;
        RECT 1051.000000 297.910000 1056.000000 298.090000 ;
        RECT 1051.000000 301.910000 1056.000000 302.090000 ;
        RECT 1101.000000 269.910000 1106.000000 270.090000 ;
        RECT 1101.000000 273.910000 1106.000000 274.090000 ;
        RECT 1101.000000 277.910000 1106.000000 278.090000 ;
        RECT 1101.000000 281.910000 1106.000000 282.090000 ;
        RECT 1101.000000 285.910000 1106.000000 286.090000 ;
        RECT 1101.000000 301.910000 1106.000000 302.090000 ;
        RECT 1101.000000 297.910000 1106.000000 298.090000 ;
        RECT 1101.000000 293.910000 1106.000000 294.090000 ;
        RECT 1101.000000 289.910000 1106.000000 290.090000 ;
        RECT 1051.000000 321.910000 1056.000000 322.090000 ;
        RECT 1051.000000 309.910000 1056.000000 310.090000 ;
        RECT 1051.000000 313.910000 1056.000000 314.090000 ;
        RECT 1051.000000 317.910000 1056.000000 318.090000 ;
        RECT 1051.000000 325.910000 1056.000000 326.090000 ;
        RECT 1051.000000 329.910000 1056.000000 330.090000 ;
        RECT 1051.000000 333.910000 1056.000000 334.090000 ;
        RECT 1051.000000 337.910000 1056.000000 338.090000 ;
        RECT 1051.000000 341.910000 1056.000000 342.090000 ;
        RECT 1101.000000 313.910000 1106.000000 314.090000 ;
        RECT 1101.000000 309.910000 1106.000000 310.090000 ;
        RECT 1101.000000 317.910000 1106.000000 318.090000 ;
        RECT 1101.000000 321.910000 1106.000000 322.090000 ;
        RECT 1101.000000 325.910000 1106.000000 326.090000 ;
        RECT 1101.000000 329.910000 1106.000000 330.090000 ;
        RECT 1101.000000 333.910000 1106.000000 334.090000 ;
        RECT 1101.000000 337.910000 1106.000000 338.090000 ;
        RECT 1101.000000 341.910000 1106.000000 342.090000 ;
        RECT 1151.000000 305.910000 1156.000000 306.090000 ;
        RECT 1172.000000 305.910000 1182.000000 306.090000 ;
        RECT 1151.000000 269.910000 1156.000000 270.090000 ;
        RECT 1151.000000 273.910000 1156.000000 274.090000 ;
        RECT 1151.000000 277.910000 1156.000000 278.090000 ;
        RECT 1151.000000 281.910000 1156.000000 282.090000 ;
        RECT 1151.000000 285.910000 1156.000000 286.090000 ;
        RECT 1172.000000 277.910000 1182.000000 278.090000 ;
        RECT 1172.000000 269.910000 1182.000000 270.090000 ;
        RECT 1172.000000 273.910000 1182.000000 274.090000 ;
        RECT 1172.000000 281.910000 1182.000000 282.090000 ;
        RECT 1172.000000 285.910000 1182.000000 286.090000 ;
        RECT 1151.000000 301.910000 1156.000000 302.090000 ;
        RECT 1151.000000 297.910000 1156.000000 298.090000 ;
        RECT 1151.000000 289.910000 1156.000000 290.090000 ;
        RECT 1151.000000 293.910000 1156.000000 294.090000 ;
        RECT 1172.000000 301.910000 1182.000000 302.090000 ;
        RECT 1172.000000 289.910000 1182.000000 290.090000 ;
        RECT 1172.000000 293.910000 1182.000000 294.090000 ;
        RECT 1172.000000 297.910000 1182.000000 298.090000 ;
        RECT 1151.000000 321.910000 1156.000000 322.090000 ;
        RECT 1151.000000 317.910000 1156.000000 318.090000 ;
        RECT 1151.000000 309.910000 1156.000000 310.090000 ;
        RECT 1151.000000 313.910000 1156.000000 314.090000 ;
        RECT 1172.000000 321.910000 1182.000000 322.090000 ;
        RECT 1172.000000 309.910000 1182.000000 310.090000 ;
        RECT 1172.000000 313.910000 1182.000000 314.090000 ;
        RECT 1172.000000 317.910000 1182.000000 318.090000 ;
        RECT 1151.000000 329.910000 1156.000000 330.090000 ;
        RECT 1151.000000 325.910000 1156.000000 326.090000 ;
        RECT 1151.000000 333.910000 1156.000000 334.090000 ;
        RECT 1151.000000 337.910000 1156.000000 338.090000 ;
        RECT 1151.000000 341.910000 1156.000000 342.090000 ;
        RECT 1172.000000 329.910000 1182.000000 330.090000 ;
        RECT 1172.000000 325.910000 1182.000000 326.090000 ;
        RECT 1172.000000 333.910000 1182.000000 334.090000 ;
        RECT 1172.000000 337.910000 1182.000000 338.090000 ;
        RECT 1172.000000 341.910000 1182.000000 342.090000 ;
        RECT 4.000000 357.910000 14.000000 358.090000 ;
        RECT 4.000000 353.910000 14.000000 354.090000 ;
        RECT 4.000000 345.910000 14.000000 346.090000 ;
        RECT 4.000000 349.910000 14.000000 350.090000 ;
        RECT 4.000000 369.910000 14.000000 370.090000 ;
        RECT 4.000000 365.910000 14.000000 366.090000 ;
        RECT 4.000000 361.910000 14.000000 362.090000 ;
        RECT 4.000000 377.910000 14.000000 378.090000 ;
        RECT 4.000000 373.910000 14.000000 374.090000 ;
        RECT 51.000000 345.910000 56.000000 346.090000 ;
        RECT 51.000000 369.910000 56.000000 370.090000 ;
        RECT 51.000000 365.910000 56.000000 366.090000 ;
        RECT 51.000000 361.910000 56.000000 362.090000 ;
        RECT 51.000000 373.910000 56.000000 374.090000 ;
        RECT 51.000000 377.910000 56.000000 378.090000 ;
        RECT 4.000000 393.910000 14.000000 394.090000 ;
        RECT 4.000000 389.910000 14.000000 390.090000 ;
        RECT 4.000000 381.910000 14.000000 382.090000 ;
        RECT 4.000000 385.910000 14.000000 386.090000 ;
        RECT 4.000000 397.910000 14.000000 398.090000 ;
        RECT 4.000000 401.910000 14.000000 402.090000 ;
        RECT 4.000000 405.910000 14.000000 406.090000 ;
        RECT 4.000000 409.910000 14.000000 410.090000 ;
        RECT 4.000000 413.910000 14.000000 414.090000 ;
        RECT 51.000000 397.910000 56.000000 398.090000 ;
        RECT 51.000000 385.910000 56.000000 386.090000 ;
        RECT 51.000000 381.910000 56.000000 382.090000 ;
        RECT 51.000000 389.910000 56.000000 390.090000 ;
        RECT 51.000000 393.910000 56.000000 394.090000 ;
        RECT 51.000000 413.910000 56.000000 414.090000 ;
        RECT 51.000000 409.910000 56.000000 410.090000 ;
        RECT 51.000000 405.910000 56.000000 406.090000 ;
        RECT 51.000000 401.910000 56.000000 402.090000 ;
        RECT 101.000000 345.910000 106.000000 346.090000 ;
        RECT 101.000000 349.910000 106.000000 350.090000 ;
        RECT 101.000000 353.910000 106.000000 354.090000 ;
        RECT 101.000000 357.910000 106.000000 358.090000 ;
        RECT 101.000000 361.910000 106.000000 362.090000 ;
        RECT 101.000000 365.910000 106.000000 366.090000 ;
        RECT 101.000000 369.910000 106.000000 370.090000 ;
        RECT 101.000000 373.910000 106.000000 374.090000 ;
        RECT 101.000000 377.910000 106.000000 378.090000 ;
        RECT 101.000000 397.910000 106.000000 398.090000 ;
        RECT 101.000000 381.910000 106.000000 382.090000 ;
        RECT 101.000000 385.910000 106.000000 386.090000 ;
        RECT 101.000000 389.910000 106.000000 390.090000 ;
        RECT 101.000000 393.910000 106.000000 394.090000 ;
        RECT 101.000000 413.910000 106.000000 414.090000 ;
        RECT 101.000000 409.910000 106.000000 410.090000 ;
        RECT 101.000000 405.910000 106.000000 406.090000 ;
        RECT 101.000000 401.910000 106.000000 402.090000 ;
        RECT 4.000000 433.910000 14.000000 434.090000 ;
        RECT 4.000000 429.910000 14.000000 430.090000 ;
        RECT 4.000000 421.910000 14.000000 422.090000 ;
        RECT 4.000000 417.910000 14.000000 418.090000 ;
        RECT 4.000000 425.910000 14.000000 426.090000 ;
        RECT 4.000000 437.910000 14.000000 438.090000 ;
        RECT 4.000000 441.910000 14.000000 442.090000 ;
        RECT 4.000000 445.910000 14.000000 446.090000 ;
        RECT 4.000000 449.910000 14.000000 450.090000 ;
        RECT 4.000000 453.910000 14.000000 454.090000 ;
        RECT 51.000000 417.910000 56.000000 418.090000 ;
        RECT 51.000000 421.910000 56.000000 422.090000 ;
        RECT 51.000000 425.910000 56.000000 426.090000 ;
        RECT 51.000000 429.910000 56.000000 430.090000 ;
        RECT 51.000000 433.910000 56.000000 434.090000 ;
        RECT 51.000000 453.910000 56.000000 454.090000 ;
        RECT 51.000000 449.910000 56.000000 450.090000 ;
        RECT 51.000000 445.910000 56.000000 446.090000 ;
        RECT 51.000000 441.910000 56.000000 442.090000 ;
        RECT 51.000000 437.910000 56.000000 438.090000 ;
        RECT 4.000000 469.910000 14.000000 470.090000 ;
        RECT 4.000000 465.910000 14.000000 466.090000 ;
        RECT 4.000000 457.910000 14.000000 458.090000 ;
        RECT 4.000000 461.910000 14.000000 462.090000 ;
        RECT 4.000000 473.910000 14.000000 474.090000 ;
        RECT 4.000000 477.910000 14.000000 478.090000 ;
        RECT 4.000000 481.910000 14.000000 482.090000 ;
        RECT 4.000000 485.910000 14.000000 486.090000 ;
        RECT 4.000000 489.910000 14.000000 490.090000 ;
        RECT 51.000000 461.910000 56.000000 462.090000 ;
        RECT 51.000000 457.910000 56.000000 458.090000 ;
        RECT 51.000000 465.910000 56.000000 466.090000 ;
        RECT 51.000000 469.910000 56.000000 470.090000 ;
        RECT 51.000000 489.910000 56.000000 490.090000 ;
        RECT 51.000000 485.910000 56.000000 486.090000 ;
        RECT 51.000000 481.910000 56.000000 482.090000 ;
        RECT 51.000000 477.910000 56.000000 478.090000 ;
        RECT 51.000000 473.910000 56.000000 474.090000 ;
        RECT 101.000000 433.910000 106.000000 434.090000 ;
        RECT 101.000000 417.910000 106.000000 418.090000 ;
        RECT 101.000000 421.910000 106.000000 422.090000 ;
        RECT 101.000000 425.910000 106.000000 426.090000 ;
        RECT 101.000000 429.910000 106.000000 430.090000 ;
        RECT 101.000000 437.910000 106.000000 438.090000 ;
        RECT 101.000000 441.910000 106.000000 442.090000 ;
        RECT 101.000000 445.910000 106.000000 446.090000 ;
        RECT 101.000000 449.910000 106.000000 450.090000 ;
        RECT 101.000000 453.910000 106.000000 454.090000 ;
        RECT 101.000000 469.910000 106.000000 470.090000 ;
        RECT 101.000000 465.910000 106.000000 466.090000 ;
        RECT 101.000000 461.910000 106.000000 462.090000 ;
        RECT 101.000000 457.910000 106.000000 458.090000 ;
        RECT 101.000000 473.910000 106.000000 474.090000 ;
        RECT 101.000000 477.910000 106.000000 478.090000 ;
        RECT 101.000000 481.910000 106.000000 482.090000 ;
        RECT 101.000000 485.910000 106.000000 486.090000 ;
        RECT 101.000000 489.910000 106.000000 490.090000 ;
        RECT 151.000000 349.910000 156.000000 350.090000 ;
        RECT 151.000000 345.910000 156.000000 346.090000 ;
        RECT 151.000000 353.910000 156.000000 354.090000 ;
        RECT 151.000000 357.910000 156.000000 358.090000 ;
        RECT 151.000000 361.910000 156.000000 362.090000 ;
        RECT 151.000000 365.910000 156.000000 366.090000 ;
        RECT 151.000000 369.910000 156.000000 370.090000 ;
        RECT 151.000000 373.910000 156.000000 374.090000 ;
        RECT 151.000000 377.910000 156.000000 378.090000 ;
        RECT 201.000000 349.910000 206.000000 350.090000 ;
        RECT 201.000000 345.910000 206.000000 346.090000 ;
        RECT 201.000000 353.910000 206.000000 354.090000 ;
        RECT 201.000000 357.910000 206.000000 358.090000 ;
        RECT 201.000000 377.910000 206.000000 378.090000 ;
        RECT 201.000000 373.910000 206.000000 374.090000 ;
        RECT 201.000000 369.910000 206.000000 370.090000 ;
        RECT 201.000000 365.910000 206.000000 366.090000 ;
        RECT 201.000000 361.910000 206.000000 362.090000 ;
        RECT 151.000000 381.910000 156.000000 382.090000 ;
        RECT 151.000000 385.910000 156.000000 386.090000 ;
        RECT 151.000000 393.910000 156.000000 394.090000 ;
        RECT 151.000000 389.910000 156.000000 390.090000 ;
        RECT 151.000000 397.910000 156.000000 398.090000 ;
        RECT 151.000000 405.910000 156.000000 406.090000 ;
        RECT 151.000000 401.910000 156.000000 402.090000 ;
        RECT 201.000000 381.910000 206.000000 382.090000 ;
        RECT 201.000000 385.910000 206.000000 386.090000 ;
        RECT 201.000000 397.910000 206.000000 398.090000 ;
        RECT 201.000000 393.910000 206.000000 394.090000 ;
        RECT 201.000000 389.910000 206.000000 390.090000 ;
        RECT 201.000000 413.910000 206.000000 414.090000 ;
        RECT 201.000000 409.910000 206.000000 410.090000 ;
        RECT 201.000000 405.910000 206.000000 406.090000 ;
        RECT 201.000000 401.910000 206.000000 402.090000 ;
        RECT 251.000000 349.910000 256.000000 350.090000 ;
        RECT 251.000000 345.910000 256.000000 346.090000 ;
        RECT 251.000000 353.910000 256.000000 354.090000 ;
        RECT 251.000000 357.910000 256.000000 358.090000 ;
        RECT 251.000000 361.910000 256.000000 362.090000 ;
        RECT 251.000000 365.910000 256.000000 366.090000 ;
        RECT 251.000000 369.910000 256.000000 370.090000 ;
        RECT 251.000000 373.910000 256.000000 374.090000 ;
        RECT 251.000000 377.910000 256.000000 378.090000 ;
        RECT 251.000000 381.910000 256.000000 382.090000 ;
        RECT 251.000000 385.910000 256.000000 386.090000 ;
        RECT 251.000000 393.910000 256.000000 394.090000 ;
        RECT 251.000000 389.910000 256.000000 390.090000 ;
        RECT 251.000000 397.910000 256.000000 398.090000 ;
        RECT 251.000000 401.910000 256.000000 402.090000 ;
        RECT 251.000000 405.910000 256.000000 406.090000 ;
        RECT 151.000000 453.910000 156.000000 454.090000 ;
        RECT 201.000000 429.910000 206.000000 430.090000 ;
        RECT 201.000000 425.910000 206.000000 426.090000 ;
        RECT 201.000000 421.910000 206.000000 422.090000 ;
        RECT 201.000000 417.910000 206.000000 418.090000 ;
        RECT 201.000000 433.910000 206.000000 434.090000 ;
        RECT 201.000000 453.910000 206.000000 454.090000 ;
        RECT 201.000000 449.910000 206.000000 450.090000 ;
        RECT 201.000000 445.910000 206.000000 446.090000 ;
        RECT 201.000000 441.910000 206.000000 442.090000 ;
        RECT 201.000000 437.910000 206.000000 438.090000 ;
        RECT 151.000000 461.910000 156.000000 462.090000 ;
        RECT 151.000000 457.910000 156.000000 458.090000 ;
        RECT 151.000000 469.910000 156.000000 470.090000 ;
        RECT 151.000000 465.910000 156.000000 466.090000 ;
        RECT 151.000000 481.910000 156.000000 482.090000 ;
        RECT 151.000000 477.910000 156.000000 478.090000 ;
        RECT 151.000000 473.910000 156.000000 474.090000 ;
        RECT 151.000000 489.910000 156.000000 490.090000 ;
        RECT 151.000000 485.910000 156.000000 486.090000 ;
        RECT 201.000000 461.910000 206.000000 462.090000 ;
        RECT 201.000000 457.910000 206.000000 458.090000 ;
        RECT 201.000000 465.910000 206.000000 466.090000 ;
        RECT 201.000000 469.910000 206.000000 470.090000 ;
        RECT 201.000000 489.910000 206.000000 490.090000 ;
        RECT 201.000000 485.910000 206.000000 486.090000 ;
        RECT 201.000000 481.910000 206.000000 482.090000 ;
        RECT 201.000000 477.910000 206.000000 478.090000 ;
        RECT 201.000000 473.910000 206.000000 474.090000 ;
        RECT 251.000000 453.910000 256.000000 454.090000 ;
        RECT 251.000000 461.910000 256.000000 462.090000 ;
        RECT 251.000000 457.910000 256.000000 458.090000 ;
        RECT 251.000000 469.910000 256.000000 470.090000 ;
        RECT 251.000000 465.910000 256.000000 466.090000 ;
        RECT 251.000000 481.910000 256.000000 482.090000 ;
        RECT 251.000000 473.910000 256.000000 474.090000 ;
        RECT 251.000000 477.910000 256.000000 478.090000 ;
        RECT 251.000000 489.910000 256.000000 490.090000 ;
        RECT 251.000000 485.910000 256.000000 486.090000 ;
        RECT 4.000000 505.910000 14.000000 506.090000 ;
        RECT 4.000000 501.910000 14.000000 502.090000 ;
        RECT 4.000000 497.910000 14.000000 498.090000 ;
        RECT 4.000000 493.910000 14.000000 494.090000 ;
        RECT 4.000000 513.910000 14.000000 514.090000 ;
        RECT 4.000000 509.910000 14.000000 510.090000 ;
        RECT 51.000000 493.910000 56.000000 494.090000 ;
        RECT 51.000000 497.910000 56.000000 498.090000 ;
        RECT 51.000000 501.910000 56.000000 502.090000 ;
        RECT 51.000000 505.910000 56.000000 506.090000 ;
        RECT 51.000000 513.910000 56.000000 514.090000 ;
        RECT 51.000000 509.910000 56.000000 510.090000 ;
        RECT 101.000000 505.910000 106.000000 506.090000 ;
        RECT 101.000000 501.910000 106.000000 502.090000 ;
        RECT 101.000000 497.910000 106.000000 498.090000 ;
        RECT 101.000000 493.910000 106.000000 494.090000 ;
        RECT 101.000000 513.910000 106.000000 514.090000 ;
        RECT 101.000000 509.910000 106.000000 510.090000 ;
        RECT 151.000000 493.910000 156.000000 494.090000 ;
        RECT 151.000000 497.910000 156.000000 498.090000 ;
        RECT 151.000000 501.910000 156.000000 502.090000 ;
        RECT 151.000000 505.910000 156.000000 506.090000 ;
        RECT 151.000000 509.910000 156.000000 510.090000 ;
        RECT 151.000000 513.910000 156.000000 514.090000 ;
        RECT 201.000000 497.910000 206.000000 498.090000 ;
        RECT 201.000000 493.910000 206.000000 494.090000 ;
        RECT 201.000000 501.910000 206.000000 502.090000 ;
        RECT 201.000000 505.910000 206.000000 506.090000 ;
        RECT 201.000000 513.910000 206.000000 514.090000 ;
        RECT 201.000000 509.910000 206.000000 510.090000 ;
        RECT 251.000000 493.910000 256.000000 494.090000 ;
        RECT 251.000000 497.910000 256.000000 498.090000 ;
        RECT 251.000000 501.910000 256.000000 502.090000 ;
        RECT 251.000000 505.910000 256.000000 506.090000 ;
        RECT 251.000000 509.910000 256.000000 510.090000 ;
        RECT 251.000000 513.910000 256.000000 514.090000 ;
        RECT 301.000000 345.910000 306.000000 346.090000 ;
        RECT 301.000000 349.910000 306.000000 350.090000 ;
        RECT 301.000000 353.910000 306.000000 354.090000 ;
        RECT 301.000000 357.910000 306.000000 358.090000 ;
        RECT 301.000000 369.910000 306.000000 370.090000 ;
        RECT 301.000000 365.910000 306.000000 366.090000 ;
        RECT 301.000000 361.910000 306.000000 362.090000 ;
        RECT 301.000000 377.910000 306.000000 378.090000 ;
        RECT 301.000000 373.910000 306.000000 374.090000 ;
        RECT 351.000000 349.910000 356.000000 350.090000 ;
        RECT 351.000000 345.910000 356.000000 346.090000 ;
        RECT 351.000000 353.910000 356.000000 354.090000 ;
        RECT 351.000000 357.910000 356.000000 358.090000 ;
        RECT 351.000000 361.910000 356.000000 362.090000 ;
        RECT 351.000000 365.910000 356.000000 366.090000 ;
        RECT 351.000000 369.910000 356.000000 370.090000 ;
        RECT 351.000000 373.910000 356.000000 374.090000 ;
        RECT 351.000000 377.910000 356.000000 378.090000 ;
        RECT 301.000000 385.910000 306.000000 386.090000 ;
        RECT 301.000000 381.910000 306.000000 382.090000 ;
        RECT 301.000000 397.910000 306.000000 398.090000 ;
        RECT 301.000000 389.910000 306.000000 390.090000 ;
        RECT 301.000000 393.910000 306.000000 394.090000 ;
        RECT 301.000000 405.910000 306.000000 406.090000 ;
        RECT 301.000000 401.910000 306.000000 402.090000 ;
        RECT 301.000000 413.910000 306.000000 414.090000 ;
        RECT 301.000000 409.910000 306.000000 410.090000 ;
        RECT 351.000000 381.910000 356.000000 382.090000 ;
        RECT 351.000000 385.910000 356.000000 386.090000 ;
        RECT 351.000000 393.910000 356.000000 394.090000 ;
        RECT 351.000000 389.910000 356.000000 390.090000 ;
        RECT 351.000000 397.910000 356.000000 398.090000 ;
        RECT 351.000000 413.910000 356.000000 414.090000 ;
        RECT 351.000000 409.910000 356.000000 410.090000 ;
        RECT 351.000000 405.910000 356.000000 406.090000 ;
        RECT 351.000000 401.910000 356.000000 402.090000 ;
        RECT 401.000000 345.910000 406.000000 346.090000 ;
        RECT 401.000000 349.910000 406.000000 350.090000 ;
        RECT 401.000000 353.910000 406.000000 354.090000 ;
        RECT 401.000000 357.910000 406.000000 358.090000 ;
        RECT 401.000000 369.910000 406.000000 370.090000 ;
        RECT 401.000000 365.910000 406.000000 366.090000 ;
        RECT 401.000000 361.910000 406.000000 362.090000 ;
        RECT 401.000000 373.910000 406.000000 374.090000 ;
        RECT 401.000000 377.910000 406.000000 378.090000 ;
        RECT 401.000000 381.910000 406.000000 382.090000 ;
        RECT 401.000000 385.910000 406.000000 386.090000 ;
        RECT 401.000000 393.910000 406.000000 394.090000 ;
        RECT 401.000000 389.910000 406.000000 390.090000 ;
        RECT 401.000000 397.910000 406.000000 398.090000 ;
        RECT 401.000000 401.910000 406.000000 402.090000 ;
        RECT 401.000000 405.910000 406.000000 406.090000 ;
        RECT 401.000000 413.910000 406.000000 414.090000 ;
        RECT 401.000000 409.910000 406.000000 410.090000 ;
        RECT 301.000000 425.910000 306.000000 426.090000 ;
        RECT 301.000000 417.910000 306.000000 418.090000 ;
        RECT 301.000000 421.910000 306.000000 422.090000 ;
        RECT 301.000000 429.910000 306.000000 430.090000 ;
        RECT 301.000000 433.910000 306.000000 434.090000 ;
        RECT 301.000000 441.910000 306.000000 442.090000 ;
        RECT 301.000000 437.910000 306.000000 438.090000 ;
        RECT 301.000000 453.910000 306.000000 454.090000 ;
        RECT 301.000000 449.910000 306.000000 450.090000 ;
        RECT 301.000000 445.910000 306.000000 446.090000 ;
        RECT 351.000000 425.910000 356.000000 426.090000 ;
        RECT 351.000000 421.910000 356.000000 422.090000 ;
        RECT 351.000000 417.910000 356.000000 418.090000 ;
        RECT 351.000000 433.910000 356.000000 434.090000 ;
        RECT 351.000000 429.910000 356.000000 430.090000 ;
        RECT 351.000000 437.910000 356.000000 438.090000 ;
        RECT 351.000000 441.910000 356.000000 442.090000 ;
        RECT 351.000000 445.910000 356.000000 446.090000 ;
        RECT 351.000000 449.910000 356.000000 450.090000 ;
        RECT 351.000000 453.910000 356.000000 454.090000 ;
        RECT 301.000000 461.910000 306.000000 462.090000 ;
        RECT 301.000000 457.910000 306.000000 458.090000 ;
        RECT 301.000000 465.910000 306.000000 466.090000 ;
        RECT 301.000000 469.910000 306.000000 470.090000 ;
        RECT 301.000000 481.910000 306.000000 482.090000 ;
        RECT 301.000000 477.910000 306.000000 478.090000 ;
        RECT 301.000000 473.910000 306.000000 474.090000 ;
        RECT 301.000000 489.910000 306.000000 490.090000 ;
        RECT 301.000000 485.910000 306.000000 486.090000 ;
        RECT 351.000000 457.910000 356.000000 458.090000 ;
        RECT 351.000000 461.910000 356.000000 462.090000 ;
        RECT 351.000000 469.910000 356.000000 470.090000 ;
        RECT 351.000000 465.910000 356.000000 466.090000 ;
        RECT 351.000000 481.910000 356.000000 482.090000 ;
        RECT 351.000000 473.910000 356.000000 474.090000 ;
        RECT 351.000000 477.910000 356.000000 478.090000 ;
        RECT 351.000000 485.910000 356.000000 486.090000 ;
        RECT 351.000000 489.910000 356.000000 490.090000 ;
        RECT 401.000000 417.910000 406.000000 418.090000 ;
        RECT 401.000000 421.910000 406.000000 422.090000 ;
        RECT 401.000000 425.910000 406.000000 426.090000 ;
        RECT 401.000000 429.910000 406.000000 430.090000 ;
        RECT 401.000000 433.910000 406.000000 434.090000 ;
        RECT 401.000000 437.910000 406.000000 438.090000 ;
        RECT 401.000000 441.910000 406.000000 442.090000 ;
        RECT 401.000000 445.910000 406.000000 446.090000 ;
        RECT 401.000000 453.910000 406.000000 454.090000 ;
        RECT 401.000000 449.910000 406.000000 450.090000 ;
        RECT 401.000000 457.910000 406.000000 458.090000 ;
        RECT 401.000000 461.910000 406.000000 462.090000 ;
        RECT 401.000000 465.910000 406.000000 466.090000 ;
        RECT 401.000000 469.910000 406.000000 470.090000 ;
        RECT 401.000000 481.910000 406.000000 482.090000 ;
        RECT 401.000000 473.910000 406.000000 474.090000 ;
        RECT 401.000000 477.910000 406.000000 478.090000 ;
        RECT 401.000000 485.910000 406.000000 486.090000 ;
        RECT 401.000000 489.910000 406.000000 490.090000 ;
        RECT 451.000000 345.910000 456.000000 346.090000 ;
        RECT 451.000000 369.910000 456.000000 370.090000 ;
        RECT 451.000000 373.910000 456.000000 374.090000 ;
        RECT 451.000000 377.910000 456.000000 378.090000 ;
        RECT 501.000000 345.910000 506.000000 346.090000 ;
        RECT 501.000000 349.910000 506.000000 350.090000 ;
        RECT 501.000000 353.910000 506.000000 354.090000 ;
        RECT 501.000000 357.910000 506.000000 358.090000 ;
        RECT 501.000000 361.910000 506.000000 362.090000 ;
        RECT 501.000000 365.910000 506.000000 366.090000 ;
        RECT 501.000000 369.910000 506.000000 370.090000 ;
        RECT 501.000000 377.910000 506.000000 378.090000 ;
        RECT 501.000000 373.910000 506.000000 374.090000 ;
        RECT 451.000000 381.910000 456.000000 382.090000 ;
        RECT 451.000000 385.910000 456.000000 386.090000 ;
        RECT 451.000000 397.910000 456.000000 398.090000 ;
        RECT 451.000000 393.910000 456.000000 394.090000 ;
        RECT 451.000000 389.910000 456.000000 390.090000 ;
        RECT 501.000000 381.910000 506.000000 382.090000 ;
        RECT 501.000000 385.910000 506.000000 386.090000 ;
        RECT 501.000000 393.910000 506.000000 394.090000 ;
        RECT 501.000000 389.910000 506.000000 390.090000 ;
        RECT 501.000000 397.910000 506.000000 398.090000 ;
        RECT 501.000000 401.910000 506.000000 402.090000 ;
        RECT 501.000000 405.910000 506.000000 406.090000 ;
        RECT 501.000000 409.910000 506.000000 410.090000 ;
        RECT 501.000000 413.910000 506.000000 414.090000 ;
        RECT 551.000000 357.910000 556.000000 358.090000 ;
        RECT 551.000000 353.910000 556.000000 354.090000 ;
        RECT 551.000000 349.910000 556.000000 350.090000 ;
        RECT 551.000000 345.910000 556.000000 346.090000 ;
        RECT 551.000000 361.910000 556.000000 362.090000 ;
        RECT 551.000000 365.910000 556.000000 366.090000 ;
        RECT 551.000000 369.910000 556.000000 370.090000 ;
        RECT 551.000000 373.910000 556.000000 374.090000 ;
        RECT 551.000000 377.910000 556.000000 378.090000 ;
        RECT 551.000000 385.910000 556.000000 386.090000 ;
        RECT 551.000000 381.910000 556.000000 382.090000 ;
        RECT 551.000000 397.910000 556.000000 398.090000 ;
        RECT 551.000000 393.910000 556.000000 394.090000 ;
        RECT 551.000000 389.910000 556.000000 390.090000 ;
        RECT 551.000000 401.910000 556.000000 402.090000 ;
        RECT 551.000000 405.910000 556.000000 406.090000 ;
        RECT 551.000000 409.910000 556.000000 410.090000 ;
        RECT 551.000000 413.910000 556.000000 414.090000 ;
        RECT 451.000000 425.910000 456.000000 426.090000 ;
        RECT 451.000000 421.910000 456.000000 422.090000 ;
        RECT 451.000000 429.910000 456.000000 430.090000 ;
        RECT 451.000000 433.910000 456.000000 434.090000 ;
        RECT 451.000000 441.910000 456.000000 442.090000 ;
        RECT 451.000000 437.910000 456.000000 438.090000 ;
        RECT 451.000000 453.910000 456.000000 454.090000 ;
        RECT 451.000000 449.910000 456.000000 450.090000 ;
        RECT 451.000000 445.910000 456.000000 446.090000 ;
        RECT 501.000000 425.910000 506.000000 426.090000 ;
        RECT 501.000000 421.910000 506.000000 422.090000 ;
        RECT 501.000000 417.910000 506.000000 418.090000 ;
        RECT 501.000000 429.910000 506.000000 430.090000 ;
        RECT 501.000000 433.910000 506.000000 434.090000 ;
        RECT 501.000000 437.910000 506.000000 438.090000 ;
        RECT 501.000000 441.910000 506.000000 442.090000 ;
        RECT 501.000000 445.910000 506.000000 446.090000 ;
        RECT 501.000000 449.910000 506.000000 450.090000 ;
        RECT 501.000000 453.910000 506.000000 454.090000 ;
        RECT 451.000000 461.910000 456.000000 462.090000 ;
        RECT 451.000000 457.910000 456.000000 458.090000 ;
        RECT 451.000000 465.910000 456.000000 466.090000 ;
        RECT 451.000000 469.910000 456.000000 470.090000 ;
        RECT 451.000000 481.910000 456.000000 482.090000 ;
        RECT 451.000000 477.910000 456.000000 478.090000 ;
        RECT 451.000000 473.910000 456.000000 474.090000 ;
        RECT 451.000000 489.910000 456.000000 490.090000 ;
        RECT 451.000000 485.910000 456.000000 486.090000 ;
        RECT 501.000000 461.910000 506.000000 462.090000 ;
        RECT 501.000000 457.910000 506.000000 458.090000 ;
        RECT 501.000000 469.910000 506.000000 470.090000 ;
        RECT 501.000000 465.910000 506.000000 466.090000 ;
        RECT 501.000000 481.910000 506.000000 482.090000 ;
        RECT 501.000000 477.910000 506.000000 478.090000 ;
        RECT 501.000000 473.910000 506.000000 474.090000 ;
        RECT 501.000000 489.910000 506.000000 490.090000 ;
        RECT 501.000000 485.910000 506.000000 486.090000 ;
        RECT 551.000000 417.910000 556.000000 418.090000 ;
        RECT 551.000000 425.910000 556.000000 426.090000 ;
        RECT 551.000000 421.910000 556.000000 422.090000 ;
        RECT 551.000000 433.910000 556.000000 434.090000 ;
        RECT 551.000000 429.910000 556.000000 430.090000 ;
        RECT 551.000000 437.910000 556.000000 438.090000 ;
        RECT 551.000000 441.910000 556.000000 442.090000 ;
        RECT 551.000000 445.910000 556.000000 446.090000 ;
        RECT 551.000000 449.910000 556.000000 450.090000 ;
        RECT 551.000000 453.910000 556.000000 454.090000 ;
        RECT 551.000000 461.910000 556.000000 462.090000 ;
        RECT 551.000000 457.910000 556.000000 458.090000 ;
        RECT 551.000000 469.910000 556.000000 470.090000 ;
        RECT 551.000000 465.910000 556.000000 466.090000 ;
        RECT 551.000000 481.910000 556.000000 482.090000 ;
        RECT 551.000000 473.910000 556.000000 474.090000 ;
        RECT 551.000000 477.910000 556.000000 478.090000 ;
        RECT 551.000000 485.910000 556.000000 486.090000 ;
        RECT 551.000000 489.910000 556.000000 490.090000 ;
        RECT 301.000000 497.910000 306.000000 498.090000 ;
        RECT 301.000000 493.910000 306.000000 494.090000 ;
        RECT 301.000000 501.910000 306.000000 502.090000 ;
        RECT 301.000000 505.910000 306.000000 506.090000 ;
        RECT 301.000000 517.910000 306.000000 518.090000 ;
        RECT 301.000000 513.910000 306.000000 514.090000 ;
        RECT 301.000000 509.910000 306.000000 510.090000 ;
        RECT 351.000000 493.910000 356.000000 494.090000 ;
        RECT 351.000000 497.910000 356.000000 498.090000 ;
        RECT 351.000000 505.910000 356.000000 506.090000 ;
        RECT 351.000000 501.910000 356.000000 502.090000 ;
        RECT 351.000000 509.910000 356.000000 510.090000 ;
        RECT 351.000000 513.910000 356.000000 514.090000 ;
        RECT 351.000000 517.910000 356.000000 518.090000 ;
        RECT 351.000000 521.910000 356.000000 522.090000 ;
        RECT 351.000000 525.910000 356.000000 526.090000 ;
        RECT 351.000000 533.910000 356.000000 534.090000 ;
        RECT 351.000000 529.910000 356.000000 530.090000 ;
        RECT 351.000000 537.910000 356.000000 538.090000 ;
        RECT 351.000000 541.910000 356.000000 542.090000 ;
        RECT 351.000000 545.910000 356.000000 546.090000 ;
        RECT 351.000000 549.910000 356.000000 550.090000 ;
        RECT 351.000000 553.910000 356.000000 554.090000 ;
        RECT 351.000000 557.910000 356.000000 558.090000 ;
        RECT 351.000000 561.910000 356.000000 562.090000 ;
        RECT 375.000000 493.910000 385.000000 494.090000 ;
        RECT 375.000000 497.910000 385.000000 498.090000 ;
        RECT 375.000000 501.910000 385.000000 502.090000 ;
        RECT 375.000000 505.910000 385.000000 506.090000 ;
        RECT 401.000000 493.910000 406.000000 494.090000 ;
        RECT 401.000000 497.910000 406.000000 498.090000 ;
        RECT 401.000000 501.910000 406.000000 502.090000 ;
        RECT 375.000000 517.910000 385.000000 518.090000 ;
        RECT 375.000000 513.910000 385.000000 514.090000 ;
        RECT 375.000000 509.910000 385.000000 510.090000 ;
        RECT 375.000000 525.910000 385.000000 526.090000 ;
        RECT 375.000000 521.910000 385.000000 522.090000 ;
        RECT 375.000000 533.910000 385.000000 534.090000 ;
        RECT 375.000000 529.910000 385.000000 530.090000 ;
        RECT 375.000000 545.910000 385.000000 546.090000 ;
        RECT 375.000000 541.910000 385.000000 542.090000 ;
        RECT 375.000000 537.910000 385.000000 538.090000 ;
        RECT 375.000000 553.910000 385.000000 554.090000 ;
        RECT 375.000000 549.910000 385.000000 550.090000 ;
        RECT 375.000000 561.910000 385.000000 562.090000 ;
        RECT 375.000000 557.910000 385.000000 558.090000 ;
        RECT 351.000000 581.910000 356.000000 582.090000 ;
        RECT 351.000000 577.910000 356.000000 578.090000 ;
        RECT 351.000000 573.910000 356.000000 574.090000 ;
        RECT 351.000000 569.910000 356.000000 570.090000 ;
        RECT 351.000000 565.910000 356.000000 566.090000 ;
        RECT 351.000000 601.910000 356.000000 602.090000 ;
        RECT 351.000000 597.910000 356.000000 598.090000 ;
        RECT 351.000000 593.910000 356.000000 594.090000 ;
        RECT 351.000000 589.910000 356.000000 590.090000 ;
        RECT 351.000000 585.910000 356.000000 586.090000 ;
        RECT 351.000000 609.910000 356.000000 610.090000 ;
        RECT 351.000000 605.910000 356.000000 606.090000 ;
        RECT 351.000000 613.910000 356.000000 614.090000 ;
        RECT 351.000000 617.910000 356.000000 618.090000 ;
        RECT 351.000000 637.910000 356.000000 638.090000 ;
        RECT 351.000000 633.910000 356.000000 634.090000 ;
        RECT 351.000000 629.910000 356.000000 630.090000 ;
        RECT 351.000000 625.910000 356.000000 626.090000 ;
        RECT 351.000000 621.910000 356.000000 622.090000 ;
        RECT 375.000000 565.910000 385.000000 566.090000 ;
        RECT 375.000000 569.910000 385.000000 570.090000 ;
        RECT 375.000000 573.910000 385.000000 574.090000 ;
        RECT 375.000000 577.910000 385.000000 578.090000 ;
        RECT 375.000000 581.910000 385.000000 582.090000 ;
        RECT 375.000000 589.910000 385.000000 590.090000 ;
        RECT 375.000000 585.910000 385.000000 586.090000 ;
        RECT 375.000000 601.910000 385.000000 602.090000 ;
        RECT 375.000000 597.910000 385.000000 598.090000 ;
        RECT 375.000000 593.910000 385.000000 594.090000 ;
        RECT 375.000000 609.910000 385.000000 610.090000 ;
        RECT 375.000000 605.910000 385.000000 606.090000 ;
        RECT 375.000000 617.910000 385.000000 618.090000 ;
        RECT 375.000000 613.910000 385.000000 614.090000 ;
        RECT 375.000000 629.910000 385.000000 630.090000 ;
        RECT 375.000000 625.910000 385.000000 626.090000 ;
        RECT 375.000000 621.910000 385.000000 622.090000 ;
        RECT 375.000000 637.910000 385.000000 638.090000 ;
        RECT 375.000000 633.910000 385.000000 634.090000 ;
        RECT 451.000000 493.910000 456.000000 494.090000 ;
        RECT 451.000000 497.910000 456.000000 498.090000 ;
        RECT 451.000000 501.910000 456.000000 502.090000 ;
        RECT 501.000000 497.910000 506.000000 498.090000 ;
        RECT 501.000000 493.910000 506.000000 494.090000 ;
        RECT 501.000000 501.910000 506.000000 502.090000 ;
        RECT 551.000000 493.910000 556.000000 494.090000 ;
        RECT 551.000000 497.910000 556.000000 498.090000 ;
        RECT 551.000000 501.910000 556.000000 502.090000 ;
        RECT 351.000000 657.910000 356.000000 658.090000 ;
        RECT 351.000000 641.910000 356.000000 642.090000 ;
        RECT 351.000000 645.910000 356.000000 646.090000 ;
        RECT 351.000000 649.910000 356.000000 650.090000 ;
        RECT 351.000000 653.910000 356.000000 654.090000 ;
        RECT 351.000000 673.910000 356.000000 674.090000 ;
        RECT 351.000000 669.910000 356.000000 670.090000 ;
        RECT 351.000000 665.910000 356.000000 666.090000 ;
        RECT 351.000000 661.910000 356.000000 662.090000 ;
        RECT 301.000000 677.910000 306.000000 678.090000 ;
        RECT 301.000000 681.910000 306.000000 682.090000 ;
        RECT 351.000000 681.910000 356.000000 682.090000 ;
        RECT 351.000000 677.910000 356.000000 678.090000 ;
        RECT 375.000000 657.910000 385.000000 658.090000 ;
        RECT 401.000000 657.910000 406.000000 658.090000 ;
        RECT 375.000000 641.910000 385.000000 642.090000 ;
        RECT 375.000000 645.910000 385.000000 646.090000 ;
        RECT 375.000000 649.910000 385.000000 650.090000 ;
        RECT 375.000000 653.910000 385.000000 654.090000 ;
        RECT 375.000000 665.910000 385.000000 666.090000 ;
        RECT 375.000000 661.910000 385.000000 662.090000 ;
        RECT 375.000000 669.910000 385.000000 670.090000 ;
        RECT 375.000000 673.910000 385.000000 674.090000 ;
        RECT 401.000000 673.910000 406.000000 674.090000 ;
        RECT 401.000000 661.910000 406.000000 662.090000 ;
        RECT 401.000000 665.910000 406.000000 666.090000 ;
        RECT 401.000000 669.910000 406.000000 670.090000 ;
        RECT 375.000000 681.910000 385.000000 682.090000 ;
        RECT 375.000000 677.910000 385.000000 678.090000 ;
        RECT 401.000000 677.910000 406.000000 678.090000 ;
        RECT 401.000000 681.910000 406.000000 682.090000 ;
        RECT 451.000000 657.910000 456.000000 658.090000 ;
        RECT 451.000000 673.910000 456.000000 674.090000 ;
        RECT 451.000000 669.910000 456.000000 670.090000 ;
        RECT 451.000000 665.910000 456.000000 666.090000 ;
        RECT 451.000000 661.910000 456.000000 662.090000 ;
        RECT 501.000000 657.910000 506.000000 658.090000 ;
        RECT 501.000000 665.910000 506.000000 666.090000 ;
        RECT 501.000000 661.910000 506.000000 662.090000 ;
        RECT 501.000000 673.910000 506.000000 674.090000 ;
        RECT 501.000000 669.910000 506.000000 670.090000 ;
        RECT 451.000000 677.910000 456.000000 678.090000 ;
        RECT 451.000000 681.910000 456.000000 682.090000 ;
        RECT 501.000000 677.910000 506.000000 678.090000 ;
        RECT 501.000000 681.910000 506.000000 682.090000 ;
        RECT 551.000000 673.910000 556.000000 674.090000 ;
        RECT 551.000000 657.910000 556.000000 658.090000 ;
        RECT 551.000000 661.910000 556.000000 662.090000 ;
        RECT 551.000000 665.910000 556.000000 666.090000 ;
        RECT 551.000000 669.910000 556.000000 670.090000 ;
        RECT 551.000000 681.910000 556.000000 682.090000 ;
        RECT 551.000000 677.910000 556.000000 678.090000 ;
        RECT 601.000000 349.910000 606.000000 350.090000 ;
        RECT 601.000000 345.910000 606.000000 346.090000 ;
        RECT 601.000000 353.910000 606.000000 354.090000 ;
        RECT 601.000000 357.910000 606.000000 358.090000 ;
        RECT 601.000000 369.910000 606.000000 370.090000 ;
        RECT 601.000000 365.910000 606.000000 366.090000 ;
        RECT 601.000000 361.910000 606.000000 362.090000 ;
        RECT 601.000000 377.910000 606.000000 378.090000 ;
        RECT 601.000000 373.910000 606.000000 374.090000 ;
        RECT 651.000000 349.910000 656.000000 350.090000 ;
        RECT 651.000000 345.910000 656.000000 346.090000 ;
        RECT 651.000000 357.910000 656.000000 358.090000 ;
        RECT 651.000000 353.910000 656.000000 354.090000 ;
        RECT 651.000000 361.910000 656.000000 362.090000 ;
        RECT 651.000000 365.910000 656.000000 366.090000 ;
        RECT 651.000000 369.910000 656.000000 370.090000 ;
        RECT 651.000000 373.910000 656.000000 374.090000 ;
        RECT 651.000000 377.910000 656.000000 378.090000 ;
        RECT 601.000000 385.910000 606.000000 386.090000 ;
        RECT 601.000000 381.910000 606.000000 382.090000 ;
        RECT 601.000000 397.910000 606.000000 398.090000 ;
        RECT 601.000000 389.910000 606.000000 390.090000 ;
        RECT 601.000000 393.910000 606.000000 394.090000 ;
        RECT 601.000000 405.910000 606.000000 406.090000 ;
        RECT 601.000000 401.910000 606.000000 402.090000 ;
        RECT 601.000000 413.910000 606.000000 414.090000 ;
        RECT 601.000000 409.910000 606.000000 410.090000 ;
        RECT 651.000000 381.910000 656.000000 382.090000 ;
        RECT 651.000000 385.910000 656.000000 386.090000 ;
        RECT 651.000000 393.910000 656.000000 394.090000 ;
        RECT 651.000000 389.910000 656.000000 390.090000 ;
        RECT 651.000000 397.910000 656.000000 398.090000 ;
        RECT 651.000000 405.910000 656.000000 406.090000 ;
        RECT 651.000000 401.910000 656.000000 402.090000 ;
        RECT 651.000000 409.910000 656.000000 410.090000 ;
        RECT 651.000000 413.910000 656.000000 414.090000 ;
        RECT 701.000000 357.910000 706.000000 358.090000 ;
        RECT 701.000000 353.910000 706.000000 354.090000 ;
        RECT 701.000000 349.910000 706.000000 350.090000 ;
        RECT 701.000000 345.910000 706.000000 346.090000 ;
        RECT 701.000000 361.910000 706.000000 362.090000 ;
        RECT 701.000000 365.910000 706.000000 366.090000 ;
        RECT 701.000000 369.910000 706.000000 370.090000 ;
        RECT 701.000000 373.910000 706.000000 374.090000 ;
        RECT 701.000000 377.910000 706.000000 378.090000 ;
        RECT 701.000000 385.910000 706.000000 386.090000 ;
        RECT 701.000000 381.910000 706.000000 382.090000 ;
        RECT 701.000000 397.910000 706.000000 398.090000 ;
        RECT 701.000000 393.910000 706.000000 394.090000 ;
        RECT 701.000000 389.910000 706.000000 390.090000 ;
        RECT 701.000000 413.910000 706.000000 414.090000 ;
        RECT 701.000000 409.910000 706.000000 410.090000 ;
        RECT 701.000000 405.910000 706.000000 406.090000 ;
        RECT 701.000000 401.910000 706.000000 402.090000 ;
        RECT 601.000000 417.910000 606.000000 418.090000 ;
        RECT 601.000000 421.910000 606.000000 422.090000 ;
        RECT 601.000000 425.910000 606.000000 426.090000 ;
        RECT 601.000000 429.910000 606.000000 430.090000 ;
        RECT 601.000000 433.910000 606.000000 434.090000 ;
        RECT 601.000000 441.910000 606.000000 442.090000 ;
        RECT 601.000000 437.910000 606.000000 438.090000 ;
        RECT 601.000000 453.910000 606.000000 454.090000 ;
        RECT 601.000000 449.910000 606.000000 450.090000 ;
        RECT 601.000000 445.910000 606.000000 446.090000 ;
        RECT 651.000000 421.910000 656.000000 422.090000 ;
        RECT 651.000000 417.910000 656.000000 418.090000 ;
        RECT 651.000000 425.910000 656.000000 426.090000 ;
        RECT 651.000000 429.910000 656.000000 430.090000 ;
        RECT 651.000000 433.910000 656.000000 434.090000 ;
        RECT 651.000000 437.910000 656.000000 438.090000 ;
        RECT 651.000000 441.910000 656.000000 442.090000 ;
        RECT 651.000000 445.910000 656.000000 446.090000 ;
        RECT 651.000000 449.910000 656.000000 450.090000 ;
        RECT 651.000000 453.910000 656.000000 454.090000 ;
        RECT 601.000000 461.910000 606.000000 462.090000 ;
        RECT 601.000000 457.910000 606.000000 458.090000 ;
        RECT 601.000000 465.910000 606.000000 466.090000 ;
        RECT 601.000000 469.910000 606.000000 470.090000 ;
        RECT 601.000000 481.910000 606.000000 482.090000 ;
        RECT 601.000000 477.910000 606.000000 478.090000 ;
        RECT 601.000000 473.910000 606.000000 474.090000 ;
        RECT 601.000000 489.910000 606.000000 490.090000 ;
        RECT 601.000000 485.910000 606.000000 486.090000 ;
        RECT 651.000000 461.910000 656.000000 462.090000 ;
        RECT 651.000000 457.910000 656.000000 458.090000 ;
        RECT 651.000000 469.910000 656.000000 470.090000 ;
        RECT 651.000000 465.910000 656.000000 466.090000 ;
        RECT 651.000000 481.910000 656.000000 482.090000 ;
        RECT 651.000000 477.910000 656.000000 478.090000 ;
        RECT 651.000000 473.910000 656.000000 474.090000 ;
        RECT 651.000000 489.910000 656.000000 490.090000 ;
        RECT 651.000000 485.910000 656.000000 486.090000 ;
        RECT 701.000000 417.910000 706.000000 418.090000 ;
        RECT 701.000000 421.910000 706.000000 422.090000 ;
        RECT 701.000000 425.910000 706.000000 426.090000 ;
        RECT 701.000000 433.910000 706.000000 434.090000 ;
        RECT 701.000000 429.910000 706.000000 430.090000 ;
        RECT 701.000000 437.910000 706.000000 438.090000 ;
        RECT 701.000000 441.910000 706.000000 442.090000 ;
        RECT 701.000000 445.910000 706.000000 446.090000 ;
        RECT 701.000000 449.910000 706.000000 450.090000 ;
        RECT 701.000000 453.910000 706.000000 454.090000 ;
        RECT 725.000000 433.910000 735.000000 434.090000 ;
        RECT 725.000000 437.910000 735.000000 438.090000 ;
        RECT 725.000000 441.910000 735.000000 442.090000 ;
        RECT 725.000000 453.910000 735.000000 454.090000 ;
        RECT 725.000000 449.910000 735.000000 450.090000 ;
        RECT 725.000000 445.910000 735.000000 446.090000 ;
        RECT 701.000000 457.910000 706.000000 458.090000 ;
        RECT 701.000000 461.910000 706.000000 462.090000 ;
        RECT 701.000000 465.910000 706.000000 466.090000 ;
        RECT 701.000000 469.910000 706.000000 470.090000 ;
        RECT 701.000000 481.910000 706.000000 482.090000 ;
        RECT 701.000000 473.910000 706.000000 474.090000 ;
        RECT 701.000000 477.910000 706.000000 478.090000 ;
        RECT 701.000000 485.910000 706.000000 486.090000 ;
        RECT 701.000000 489.910000 706.000000 490.090000 ;
        RECT 725.000000 469.910000 735.000000 470.090000 ;
        RECT 725.000000 465.910000 735.000000 466.090000 ;
        RECT 725.000000 457.910000 735.000000 458.090000 ;
        RECT 725.000000 461.910000 735.000000 462.090000 ;
        RECT 725.000000 481.910000 735.000000 482.090000 ;
        RECT 725.000000 477.910000 735.000000 478.090000 ;
        RECT 725.000000 473.910000 735.000000 474.090000 ;
        RECT 725.000000 489.910000 735.000000 490.090000 ;
        RECT 725.000000 485.910000 735.000000 486.090000 ;
        RECT 751.000000 349.910000 756.000000 350.090000 ;
        RECT 751.000000 345.910000 756.000000 346.090000 ;
        RECT 751.000000 353.910000 756.000000 354.090000 ;
        RECT 751.000000 357.910000 756.000000 358.090000 ;
        RECT 751.000000 369.910000 756.000000 370.090000 ;
        RECT 751.000000 365.910000 756.000000 366.090000 ;
        RECT 751.000000 361.910000 756.000000 362.090000 ;
        RECT 751.000000 373.910000 756.000000 374.090000 ;
        RECT 751.000000 377.910000 756.000000 378.090000 ;
        RECT 801.000000 345.910000 806.000000 346.090000 ;
        RECT 801.000000 349.910000 806.000000 350.090000 ;
        RECT 801.000000 353.910000 806.000000 354.090000 ;
        RECT 801.000000 357.910000 806.000000 358.090000 ;
        RECT 801.000000 361.910000 806.000000 362.090000 ;
        RECT 801.000000 365.910000 806.000000 366.090000 ;
        RECT 801.000000 369.910000 806.000000 370.090000 ;
        RECT 801.000000 373.910000 806.000000 374.090000 ;
        RECT 801.000000 377.910000 806.000000 378.090000 ;
        RECT 751.000000 393.910000 756.000000 394.090000 ;
        RECT 751.000000 389.910000 756.000000 390.090000 ;
        RECT 751.000000 381.910000 756.000000 382.090000 ;
        RECT 751.000000 385.910000 756.000000 386.090000 ;
        RECT 751.000000 397.910000 756.000000 398.090000 ;
        RECT 751.000000 401.910000 756.000000 402.090000 ;
        RECT 751.000000 405.910000 756.000000 406.090000 ;
        RECT 751.000000 409.910000 756.000000 410.090000 ;
        RECT 751.000000 413.910000 756.000000 414.090000 ;
        RECT 801.000000 385.910000 806.000000 386.090000 ;
        RECT 801.000000 381.910000 806.000000 382.090000 ;
        RECT 801.000000 393.910000 806.000000 394.090000 ;
        RECT 801.000000 389.910000 806.000000 390.090000 ;
        RECT 801.000000 397.910000 806.000000 398.090000 ;
        RECT 801.000000 405.910000 806.000000 406.090000 ;
        RECT 801.000000 401.910000 806.000000 402.090000 ;
        RECT 801.000000 409.910000 806.000000 410.090000 ;
        RECT 801.000000 413.910000 806.000000 414.090000 ;
        RECT 851.000000 357.910000 856.000000 358.090000 ;
        RECT 851.000000 353.910000 856.000000 354.090000 ;
        RECT 851.000000 349.910000 856.000000 350.090000 ;
        RECT 851.000000 345.910000 856.000000 346.090000 ;
        RECT 851.000000 361.910000 856.000000 362.090000 ;
        RECT 851.000000 365.910000 856.000000 366.090000 ;
        RECT 851.000000 369.910000 856.000000 370.090000 ;
        RECT 851.000000 373.910000 856.000000 374.090000 ;
        RECT 851.000000 377.910000 856.000000 378.090000 ;
        RECT 851.000000 385.910000 856.000000 386.090000 ;
        RECT 851.000000 381.910000 856.000000 382.090000 ;
        RECT 851.000000 397.910000 856.000000 398.090000 ;
        RECT 851.000000 393.910000 856.000000 394.090000 ;
        RECT 851.000000 389.910000 856.000000 390.090000 ;
        RECT 851.000000 413.910000 856.000000 414.090000 ;
        RECT 851.000000 409.910000 856.000000 410.090000 ;
        RECT 851.000000 405.910000 856.000000 406.090000 ;
        RECT 851.000000 401.910000 856.000000 402.090000 ;
        RECT 751.000000 421.910000 756.000000 422.090000 ;
        RECT 751.000000 417.910000 756.000000 418.090000 ;
        RECT 751.000000 425.910000 756.000000 426.090000 ;
        RECT 751.000000 429.910000 756.000000 430.090000 ;
        RECT 751.000000 433.910000 756.000000 434.090000 ;
        RECT 751.000000 437.910000 756.000000 438.090000 ;
        RECT 751.000000 441.910000 756.000000 442.090000 ;
        RECT 801.000000 425.910000 806.000000 426.090000 ;
        RECT 801.000000 421.910000 806.000000 422.090000 ;
        RECT 801.000000 417.910000 806.000000 418.090000 ;
        RECT 801.000000 433.910000 806.000000 434.090000 ;
        RECT 801.000000 429.910000 806.000000 430.090000 ;
        RECT 801.000000 437.910000 806.000000 438.090000 ;
        RECT 801.000000 441.910000 806.000000 442.090000 ;
        RECT 851.000000 417.910000 856.000000 418.090000 ;
        RECT 851.000000 421.910000 856.000000 422.090000 ;
        RECT 851.000000 425.910000 856.000000 426.090000 ;
        RECT 851.000000 433.910000 856.000000 434.090000 ;
        RECT 851.000000 429.910000 856.000000 430.090000 ;
        RECT 851.000000 441.910000 856.000000 442.090000 ;
        RECT 851.000000 437.910000 856.000000 438.090000 ;
        RECT 601.000000 493.910000 606.000000 494.090000 ;
        RECT 601.000000 497.910000 606.000000 498.090000 ;
        RECT 601.000000 501.910000 606.000000 502.090000 ;
        RECT 651.000000 497.910000 656.000000 498.090000 ;
        RECT 651.000000 493.910000 656.000000 494.090000 ;
        RECT 651.000000 501.910000 656.000000 502.090000 ;
        RECT 701.000000 501.910000 706.000000 502.090000 ;
        RECT 701.000000 493.910000 706.000000 494.090000 ;
        RECT 701.000000 497.910000 706.000000 498.090000 ;
        RECT 725.000000 497.910000 735.000000 498.090000 ;
        RECT 725.000000 493.910000 735.000000 494.090000 ;
        RECT 725.000000 501.910000 735.000000 502.090000 ;
        RECT 901.000000 357.910000 906.000000 358.090000 ;
        RECT 901.000000 353.910000 906.000000 354.090000 ;
        RECT 901.000000 349.910000 906.000000 350.090000 ;
        RECT 901.000000 345.910000 906.000000 346.090000 ;
        RECT 901.000000 369.910000 906.000000 370.090000 ;
        RECT 901.000000 365.910000 906.000000 366.090000 ;
        RECT 901.000000 361.910000 906.000000 362.090000 ;
        RECT 901.000000 373.910000 906.000000 374.090000 ;
        RECT 901.000000 377.910000 906.000000 378.090000 ;
        RECT 951.000000 345.910000 956.000000 346.090000 ;
        RECT 951.000000 349.910000 956.000000 350.090000 ;
        RECT 951.000000 353.910000 956.000000 354.090000 ;
        RECT 951.000000 357.910000 956.000000 358.090000 ;
        RECT 951.000000 369.910000 956.000000 370.090000 ;
        RECT 951.000000 365.910000 956.000000 366.090000 ;
        RECT 951.000000 361.910000 956.000000 362.090000 ;
        RECT 951.000000 377.910000 956.000000 378.090000 ;
        RECT 951.000000 373.910000 956.000000 374.090000 ;
        RECT 901.000000 393.910000 906.000000 394.090000 ;
        RECT 901.000000 389.910000 906.000000 390.090000 ;
        RECT 901.000000 381.910000 906.000000 382.090000 ;
        RECT 901.000000 385.910000 906.000000 386.090000 ;
        RECT 901.000000 397.910000 906.000000 398.090000 ;
        RECT 901.000000 401.910000 906.000000 402.090000 ;
        RECT 901.000000 405.910000 906.000000 406.090000 ;
        RECT 901.000000 413.910000 906.000000 414.090000 ;
        RECT 901.000000 409.910000 906.000000 410.090000 ;
        RECT 951.000000 397.910000 956.000000 398.090000 ;
        RECT 951.000000 393.910000 956.000000 394.090000 ;
        RECT 951.000000 389.910000 956.000000 390.090000 ;
        RECT 951.000000 381.910000 956.000000 382.090000 ;
        RECT 951.000000 385.910000 956.000000 386.090000 ;
        RECT 951.000000 405.910000 956.000000 406.090000 ;
        RECT 951.000000 401.910000 956.000000 402.090000 ;
        RECT 951.000000 413.910000 956.000000 414.090000 ;
        RECT 951.000000 409.910000 956.000000 410.090000 ;
        RECT 1001.000000 349.910000 1006.000000 350.090000 ;
        RECT 1001.000000 345.910000 1006.000000 346.090000 ;
        RECT 1001.000000 353.910000 1006.000000 354.090000 ;
        RECT 1001.000000 357.910000 1006.000000 358.090000 ;
        RECT 1001.000000 361.910000 1006.000000 362.090000 ;
        RECT 1001.000000 365.910000 1006.000000 366.090000 ;
        RECT 1001.000000 369.910000 1006.000000 370.090000 ;
        RECT 1001.000000 373.910000 1006.000000 374.090000 ;
        RECT 1001.000000 377.910000 1006.000000 378.090000 ;
        RECT 1001.000000 385.910000 1006.000000 386.090000 ;
        RECT 1001.000000 381.910000 1006.000000 382.090000 ;
        RECT 1001.000000 397.910000 1006.000000 398.090000 ;
        RECT 1001.000000 389.910000 1006.000000 390.090000 ;
        RECT 1001.000000 393.910000 1006.000000 394.090000 ;
        RECT 1001.000000 401.910000 1006.000000 402.090000 ;
        RECT 1001.000000 405.910000 1006.000000 406.090000 ;
        RECT 1001.000000 409.910000 1006.000000 410.090000 ;
        RECT 1001.000000 413.910000 1006.000000 414.090000 ;
        RECT 901.000000 417.910000 906.000000 418.090000 ;
        RECT 901.000000 421.910000 906.000000 422.090000 ;
        RECT 901.000000 425.910000 906.000000 426.090000 ;
        RECT 901.000000 429.910000 906.000000 430.090000 ;
        RECT 901.000000 433.910000 906.000000 434.090000 ;
        RECT 901.000000 437.910000 906.000000 438.090000 ;
        RECT 901.000000 441.910000 906.000000 442.090000 ;
        RECT 951.000000 433.910000 956.000000 434.090000 ;
        RECT 951.000000 429.910000 956.000000 430.090000 ;
        RECT 951.000000 425.910000 956.000000 426.090000 ;
        RECT 951.000000 421.910000 956.000000 422.090000 ;
        RECT 951.000000 417.910000 956.000000 418.090000 ;
        RECT 951.000000 437.910000 956.000000 438.090000 ;
        RECT 951.000000 441.910000 956.000000 442.090000 ;
        RECT 1001.000000 425.910000 1006.000000 426.090000 ;
        RECT 1001.000000 421.910000 1006.000000 422.090000 ;
        RECT 1001.000000 417.910000 1006.000000 418.090000 ;
        RECT 1001.000000 429.910000 1006.000000 430.090000 ;
        RECT 1001.000000 433.910000 1006.000000 434.090000 ;
        RECT 1001.000000 437.910000 1006.000000 438.090000 ;
        RECT 1001.000000 441.910000 1006.000000 442.090000 ;
        RECT 1051.000000 357.910000 1056.000000 358.090000 ;
        RECT 1051.000000 353.910000 1056.000000 354.090000 ;
        RECT 1051.000000 349.910000 1056.000000 350.090000 ;
        RECT 1051.000000 345.910000 1056.000000 346.090000 ;
        RECT 1051.000000 369.910000 1056.000000 370.090000 ;
        RECT 1051.000000 365.910000 1056.000000 366.090000 ;
        RECT 1051.000000 361.910000 1056.000000 362.090000 ;
        RECT 1051.000000 373.910000 1056.000000 374.090000 ;
        RECT 1051.000000 377.910000 1056.000000 378.090000 ;
        RECT 1101.000000 345.910000 1106.000000 346.090000 ;
        RECT 1101.000000 349.910000 1106.000000 350.090000 ;
        RECT 1101.000000 353.910000 1106.000000 354.090000 ;
        RECT 1101.000000 357.910000 1106.000000 358.090000 ;
        RECT 1101.000000 369.910000 1106.000000 370.090000 ;
        RECT 1101.000000 365.910000 1106.000000 366.090000 ;
        RECT 1101.000000 361.910000 1106.000000 362.090000 ;
        RECT 1101.000000 377.910000 1106.000000 378.090000 ;
        RECT 1101.000000 373.910000 1106.000000 374.090000 ;
        RECT 1051.000000 393.910000 1056.000000 394.090000 ;
        RECT 1051.000000 389.910000 1056.000000 390.090000 ;
        RECT 1051.000000 381.910000 1056.000000 382.090000 ;
        RECT 1051.000000 385.910000 1056.000000 386.090000 ;
        RECT 1051.000000 397.910000 1056.000000 398.090000 ;
        RECT 1051.000000 405.910000 1056.000000 406.090000 ;
        RECT 1051.000000 401.910000 1056.000000 402.090000 ;
        RECT 1051.000000 413.910000 1056.000000 414.090000 ;
        RECT 1051.000000 409.910000 1056.000000 410.090000 ;
        RECT 1101.000000 397.910000 1106.000000 398.090000 ;
        RECT 1101.000000 393.910000 1106.000000 394.090000 ;
        RECT 1101.000000 389.910000 1106.000000 390.090000 ;
        RECT 1101.000000 381.910000 1106.000000 382.090000 ;
        RECT 1101.000000 385.910000 1106.000000 386.090000 ;
        RECT 1101.000000 405.910000 1106.000000 406.090000 ;
        RECT 1101.000000 401.910000 1106.000000 402.090000 ;
        RECT 1101.000000 413.910000 1106.000000 414.090000 ;
        RECT 1101.000000 409.910000 1106.000000 410.090000 ;
        RECT 1151.000000 357.910000 1156.000000 358.090000 ;
        RECT 1151.000000 353.910000 1156.000000 354.090000 ;
        RECT 1151.000000 349.910000 1156.000000 350.090000 ;
        RECT 1151.000000 345.910000 1156.000000 346.090000 ;
        RECT 1172.000000 357.910000 1182.000000 358.090000 ;
        RECT 1172.000000 349.910000 1182.000000 350.090000 ;
        RECT 1172.000000 345.910000 1182.000000 346.090000 ;
        RECT 1172.000000 353.910000 1182.000000 354.090000 ;
        RECT 1151.000000 365.910000 1156.000000 366.090000 ;
        RECT 1151.000000 361.910000 1156.000000 362.090000 ;
        RECT 1151.000000 369.910000 1156.000000 370.090000 ;
        RECT 1151.000000 377.910000 1156.000000 378.090000 ;
        RECT 1151.000000 373.910000 1156.000000 374.090000 ;
        RECT 1172.000000 369.910000 1182.000000 370.090000 ;
        RECT 1172.000000 365.910000 1182.000000 366.090000 ;
        RECT 1172.000000 361.910000 1182.000000 362.090000 ;
        RECT 1172.000000 373.910000 1182.000000 374.090000 ;
        RECT 1172.000000 377.910000 1182.000000 378.090000 ;
        RECT 1151.000000 385.910000 1156.000000 386.090000 ;
        RECT 1151.000000 381.910000 1156.000000 382.090000 ;
        RECT 1151.000000 389.910000 1156.000000 390.090000 ;
        RECT 1151.000000 393.910000 1156.000000 394.090000 ;
        RECT 1151.000000 397.910000 1156.000000 398.090000 ;
        RECT 1172.000000 385.910000 1182.000000 386.090000 ;
        RECT 1172.000000 381.910000 1182.000000 382.090000 ;
        RECT 1172.000000 389.910000 1182.000000 390.090000 ;
        RECT 1172.000000 393.910000 1182.000000 394.090000 ;
        RECT 1172.000000 397.910000 1182.000000 398.090000 ;
        RECT 1151.000000 405.910000 1156.000000 406.090000 ;
        RECT 1151.000000 401.910000 1156.000000 402.090000 ;
        RECT 1151.000000 409.910000 1156.000000 410.090000 ;
        RECT 1151.000000 413.910000 1156.000000 414.090000 ;
        RECT 1172.000000 405.910000 1182.000000 406.090000 ;
        RECT 1172.000000 401.910000 1182.000000 402.090000 ;
        RECT 1172.000000 409.910000 1182.000000 410.090000 ;
        RECT 1172.000000 413.910000 1182.000000 414.090000 ;
        RECT 1051.000000 417.910000 1056.000000 418.090000 ;
        RECT 1051.000000 421.910000 1056.000000 422.090000 ;
        RECT 1051.000000 425.910000 1056.000000 426.090000 ;
        RECT 1051.000000 429.910000 1056.000000 430.090000 ;
        RECT 1051.000000 433.910000 1056.000000 434.090000 ;
        RECT 1051.000000 437.910000 1056.000000 438.090000 ;
        RECT 1051.000000 441.910000 1056.000000 442.090000 ;
        RECT 1101.000000 433.910000 1106.000000 434.090000 ;
        RECT 1101.000000 429.910000 1106.000000 430.090000 ;
        RECT 1101.000000 425.910000 1106.000000 426.090000 ;
        RECT 1101.000000 421.910000 1106.000000 422.090000 ;
        RECT 1101.000000 417.910000 1106.000000 418.090000 ;
        RECT 1101.000000 441.910000 1106.000000 442.090000 ;
        RECT 1101.000000 437.910000 1106.000000 438.090000 ;
        RECT 1151.000000 417.910000 1156.000000 418.090000 ;
        RECT 1151.000000 421.910000 1156.000000 422.090000 ;
        RECT 1151.000000 425.910000 1156.000000 426.090000 ;
        RECT 1151.000000 429.910000 1156.000000 430.090000 ;
        RECT 1151.000000 433.910000 1156.000000 434.090000 ;
        RECT 1172.000000 417.910000 1182.000000 418.090000 ;
        RECT 1172.000000 421.910000 1182.000000 422.090000 ;
        RECT 1172.000000 425.910000 1182.000000 426.090000 ;
        RECT 1172.000000 429.910000 1182.000000 430.090000 ;
        RECT 1172.000000 433.910000 1182.000000 434.090000 ;
        RECT 1151.000000 437.910000 1156.000000 438.090000 ;
        RECT 1151.000000 441.910000 1156.000000 442.090000 ;
        RECT 1151.000000 453.910000 1156.000000 454.090000 ;
        RECT 1151.000000 449.910000 1156.000000 450.090000 ;
        RECT 1151.000000 445.910000 1156.000000 446.090000 ;
        RECT 1172.000000 437.910000 1182.000000 438.090000 ;
        RECT 1172.000000 441.910000 1182.000000 442.090000 ;
        RECT 1151.000000 461.910000 1156.000000 462.090000 ;
        RECT 1151.000000 457.910000 1156.000000 458.090000 ;
        RECT 1151.000000 465.910000 1156.000000 466.090000 ;
        RECT 1151.000000 469.910000 1156.000000 470.090000 ;
        RECT 1151.000000 481.910000 1156.000000 482.090000 ;
        RECT 1151.000000 477.910000 1156.000000 478.090000 ;
        RECT 1151.000000 473.910000 1156.000000 474.090000 ;
        RECT 1151.000000 489.910000 1156.000000 490.090000 ;
        RECT 1151.000000 485.910000 1156.000000 486.090000 ;
        RECT 1151.000000 493.910000 1156.000000 494.090000 ;
        RECT 1151.000000 497.910000 1156.000000 498.090000 ;
        RECT 1151.000000 505.910000 1156.000000 506.090000 ;
        RECT 1151.000000 501.910000 1156.000000 502.090000 ;
        RECT 1151.000000 509.910000 1156.000000 510.090000 ;
        RECT 1151.000000 513.910000 1156.000000 514.090000 ;
        RECT 1151.000000 517.910000 1156.000000 518.090000 ;
        RECT 1151.000000 521.910000 1156.000000 522.090000 ;
        RECT 1151.000000 525.910000 1156.000000 526.090000 ;
        RECT 1151.000000 533.910000 1156.000000 534.090000 ;
        RECT 1151.000000 529.910000 1156.000000 530.090000 ;
        RECT 1151.000000 545.910000 1156.000000 546.090000 ;
        RECT 1151.000000 537.910000 1156.000000 538.090000 ;
        RECT 1151.000000 541.910000 1156.000000 542.090000 ;
        RECT 1151.000000 549.910000 1156.000000 550.090000 ;
        RECT 1151.000000 553.910000 1156.000000 554.090000 ;
        RECT 1151.000000 561.910000 1156.000000 562.090000 ;
        RECT 1151.000000 557.910000 1156.000000 558.090000 ;
        RECT 1151.000000 565.910000 1156.000000 566.090000 ;
        RECT 1151.000000 569.910000 1156.000000 570.090000 ;
        RECT 1151.000000 573.910000 1156.000000 574.090000 ;
        RECT 1151.000000 577.910000 1156.000000 578.090000 ;
        RECT 1151.000000 581.910000 1156.000000 582.090000 ;
        RECT 1151.000000 585.910000 1156.000000 586.090000 ;
        RECT 1151.000000 589.910000 1156.000000 590.090000 ;
        RECT 1151.000000 593.910000 1156.000000 594.090000 ;
        RECT 1151.000000 597.910000 1156.000000 598.090000 ;
        RECT 1151.000000 601.910000 1156.000000 602.090000 ;
        RECT 1151.000000 609.910000 1156.000000 610.090000 ;
        RECT 1151.000000 605.910000 1156.000000 606.090000 ;
        RECT 1151.000000 613.910000 1156.000000 614.090000 ;
        RECT 1151.000000 617.910000 1156.000000 618.090000 ;
        RECT 1151.000000 621.910000 1156.000000 622.090000 ;
        RECT 1151.000000 625.910000 1156.000000 626.090000 ;
        RECT 1151.000000 629.910000 1156.000000 630.090000 ;
        RECT 1151.000000 637.910000 1156.000000 638.090000 ;
        RECT 1151.000000 633.910000 1156.000000 634.090000 ;
        RECT 601.000000 657.910000 606.000000 658.090000 ;
        RECT 601.000000 673.910000 606.000000 674.090000 ;
        RECT 601.000000 669.910000 606.000000 670.090000 ;
        RECT 601.000000 665.910000 606.000000 666.090000 ;
        RECT 601.000000 661.910000 606.000000 662.090000 ;
        RECT 651.000000 657.910000 656.000000 658.090000 ;
        RECT 651.000000 665.910000 656.000000 666.090000 ;
        RECT 651.000000 661.910000 656.000000 662.090000 ;
        RECT 651.000000 673.910000 656.000000 674.090000 ;
        RECT 651.000000 669.910000 656.000000 670.090000 ;
        RECT 601.000000 677.910000 606.000000 678.090000 ;
        RECT 601.000000 681.910000 606.000000 682.090000 ;
        RECT 651.000000 677.910000 656.000000 678.090000 ;
        RECT 651.000000 681.910000 656.000000 682.090000 ;
        RECT 1151.000000 657.910000 1156.000000 658.090000 ;
        RECT 1151.000000 641.910000 1156.000000 642.090000 ;
        RECT 1151.000000 645.910000 1156.000000 646.090000 ;
        RECT 1151.000000 649.910000 1156.000000 650.090000 ;
        RECT 1151.000000 653.910000 1156.000000 654.090000 ;
        RECT 1151.000000 665.910000 1156.000000 666.090000 ;
        RECT 1151.000000 661.910000 1156.000000 662.090000 ;
        RECT 1151.000000 669.910000 1156.000000 670.090000 ;
        RECT 1151.000000 673.910000 1156.000000 674.090000 ;
        RECT 1151.000000 681.910000 1156.000000 682.090000 ;
        RECT 1151.000000 677.910000 1156.000000 678.090000 ;
      LAYER M3 ;
        RECT 4.000000 5.910000 14.000000 6.090000 ;
        RECT 51.000000 5.910000 56.000000 6.090000 ;
        RECT 51.000000 1.910000 56.000000 2.090000 ;
        RECT 101.000000 1.910000 106.000000 2.090000 ;
        RECT 101.000000 5.910000 106.000000 6.090000 ;
        RECT 151.000000 1.910000 156.000000 2.090000 ;
        RECT 151.000000 5.910000 156.000000 6.090000 ;
        RECT 201.000000 1.910000 206.000000 2.090000 ;
        RECT 201.000000 5.910000 206.000000 6.090000 ;
        RECT 251.000000 1.910000 256.000000 2.090000 ;
        RECT 251.000000 5.910000 256.000000 6.090000 ;
        RECT 301.000000 1.910000 306.000000 2.090000 ;
        RECT 301.000000 5.910000 306.000000 6.090000 ;
        RECT 351.000000 1.910000 356.000000 2.090000 ;
        RECT 351.000000 5.910000 356.000000 6.090000 ;
        RECT 401.000000 1.910000 406.000000 2.090000 ;
        RECT 401.000000 5.910000 406.000000 6.090000 ;
        RECT 451.000000 1.910000 456.000000 2.090000 ;
        RECT 451.000000 5.910000 456.000000 6.090000 ;
        RECT 501.000000 1.910000 506.000000 2.090000 ;
        RECT 501.000000 5.910000 506.000000 6.090000 ;
        RECT 551.000000 1.910000 556.000000 2.090000 ;
        RECT 551.000000 5.910000 556.000000 6.090000 ;
        RECT 4.000000 265.910000 14.000000 266.090000 ;
        RECT 4.000000 261.910000 14.000000 262.090000 ;
        RECT 51.000000 265.910000 56.000000 266.090000 ;
        RECT 51.000000 261.910000 56.000000 262.090000 ;
        RECT 101.000000 265.910000 106.000000 266.090000 ;
        RECT 101.000000 261.910000 106.000000 262.090000 ;
        RECT 51.000000 305.910000 56.000000 306.090000 ;
        RECT 4.000000 305.910000 14.000000 306.090000 ;
        RECT 4.000000 285.910000 14.000000 286.090000 ;
        RECT 4.000000 281.910000 14.000000 282.090000 ;
        RECT 4.000000 269.910000 14.000000 270.090000 ;
        RECT 4.000000 273.910000 14.000000 274.090000 ;
        RECT 4.000000 277.910000 14.000000 278.090000 ;
        RECT 4.000000 289.910000 14.000000 290.090000 ;
        RECT 4.000000 293.910000 14.000000 294.090000 ;
        RECT 4.000000 297.910000 14.000000 298.090000 ;
        RECT 4.000000 301.910000 14.000000 302.090000 ;
        RECT 51.000000 269.910000 56.000000 270.090000 ;
        RECT 51.000000 273.910000 56.000000 274.090000 ;
        RECT 51.000000 277.910000 56.000000 278.090000 ;
        RECT 51.000000 281.910000 56.000000 282.090000 ;
        RECT 51.000000 285.910000 56.000000 286.090000 ;
        RECT 51.000000 301.910000 56.000000 302.090000 ;
        RECT 51.000000 297.910000 56.000000 298.090000 ;
        RECT 51.000000 293.910000 56.000000 294.090000 ;
        RECT 51.000000 289.910000 56.000000 290.090000 ;
        RECT 4.000000 321.910000 14.000000 322.090000 ;
        RECT 4.000000 309.910000 14.000000 310.090000 ;
        RECT 4.000000 313.910000 14.000000 314.090000 ;
        RECT 4.000000 317.910000 14.000000 318.090000 ;
        RECT 4.000000 325.910000 14.000000 326.090000 ;
        RECT 4.000000 329.910000 14.000000 330.090000 ;
        RECT 4.000000 333.910000 14.000000 334.090000 ;
        RECT 4.000000 337.910000 14.000000 338.090000 ;
        RECT 4.000000 341.910000 14.000000 342.090000 ;
        RECT 51.000000 313.910000 56.000000 314.090000 ;
        RECT 51.000000 309.910000 56.000000 310.090000 ;
        RECT 51.000000 317.910000 56.000000 318.090000 ;
        RECT 51.000000 321.910000 56.000000 322.090000 ;
        RECT 51.000000 341.910000 56.000000 342.090000 ;
        RECT 51.000000 337.910000 56.000000 338.090000 ;
        RECT 51.000000 333.910000 56.000000 334.090000 ;
        RECT 51.000000 329.910000 56.000000 330.090000 ;
        RECT 51.000000 325.910000 56.000000 326.090000 ;
        RECT 101.000000 305.910000 106.000000 306.090000 ;
        RECT 101.000000 269.910000 106.000000 270.090000 ;
        RECT 101.000000 273.910000 106.000000 274.090000 ;
        RECT 101.000000 277.910000 106.000000 278.090000 ;
        RECT 101.000000 281.910000 106.000000 282.090000 ;
        RECT 101.000000 285.910000 106.000000 286.090000 ;
        RECT 101.000000 301.910000 106.000000 302.090000 ;
        RECT 101.000000 297.910000 106.000000 298.090000 ;
        RECT 101.000000 293.910000 106.000000 294.090000 ;
        RECT 101.000000 289.910000 106.000000 290.090000 ;
        RECT 101.000000 321.910000 106.000000 322.090000 ;
        RECT 101.000000 317.910000 106.000000 318.090000 ;
        RECT 101.000000 313.910000 106.000000 314.090000 ;
        RECT 101.000000 309.910000 106.000000 310.090000 ;
        RECT 101.000000 325.910000 106.000000 326.090000 ;
        RECT 101.000000 329.910000 106.000000 330.090000 ;
        RECT 101.000000 333.910000 106.000000 334.090000 ;
        RECT 101.000000 337.910000 106.000000 338.090000 ;
        RECT 101.000000 341.910000 106.000000 342.090000 ;
        RECT 151.000000 261.910000 156.000000 262.090000 ;
        RECT 151.000000 265.910000 156.000000 266.090000 ;
        RECT 201.000000 265.910000 206.000000 266.090000 ;
        RECT 201.000000 261.910000 206.000000 262.090000 ;
        RECT 251.000000 265.910000 256.000000 266.090000 ;
        RECT 251.000000 261.910000 256.000000 262.090000 ;
        RECT 201.000000 305.910000 206.000000 306.090000 ;
        RECT 151.000000 305.910000 156.000000 306.090000 ;
        RECT 151.000000 269.910000 156.000000 270.090000 ;
        RECT 151.000000 273.910000 156.000000 274.090000 ;
        RECT 151.000000 277.910000 156.000000 278.090000 ;
        RECT 151.000000 281.910000 156.000000 282.090000 ;
        RECT 151.000000 285.910000 156.000000 286.090000 ;
        RECT 151.000000 289.910000 156.000000 290.090000 ;
        RECT 151.000000 293.910000 156.000000 294.090000 ;
        RECT 151.000000 301.910000 156.000000 302.090000 ;
        RECT 151.000000 297.910000 156.000000 298.090000 ;
        RECT 201.000000 269.910000 206.000000 270.090000 ;
        RECT 201.000000 273.910000 206.000000 274.090000 ;
        RECT 201.000000 277.910000 206.000000 278.090000 ;
        RECT 201.000000 281.910000 206.000000 282.090000 ;
        RECT 201.000000 285.910000 206.000000 286.090000 ;
        RECT 201.000000 301.910000 206.000000 302.090000 ;
        RECT 201.000000 297.910000 206.000000 298.090000 ;
        RECT 201.000000 293.910000 206.000000 294.090000 ;
        RECT 201.000000 289.910000 206.000000 290.090000 ;
        RECT 151.000000 313.910000 156.000000 314.090000 ;
        RECT 151.000000 309.910000 156.000000 310.090000 ;
        RECT 151.000000 321.910000 156.000000 322.090000 ;
        RECT 151.000000 317.910000 156.000000 318.090000 ;
        RECT 151.000000 329.910000 156.000000 330.090000 ;
        RECT 151.000000 325.910000 156.000000 326.090000 ;
        RECT 151.000000 333.910000 156.000000 334.090000 ;
        RECT 151.000000 337.910000 156.000000 338.090000 ;
        RECT 151.000000 341.910000 156.000000 342.090000 ;
        RECT 201.000000 313.910000 206.000000 314.090000 ;
        RECT 201.000000 309.910000 206.000000 310.090000 ;
        RECT 201.000000 317.910000 206.000000 318.090000 ;
        RECT 201.000000 321.910000 206.000000 322.090000 ;
        RECT 201.000000 341.910000 206.000000 342.090000 ;
        RECT 201.000000 337.910000 206.000000 338.090000 ;
        RECT 201.000000 333.910000 206.000000 334.090000 ;
        RECT 201.000000 329.910000 206.000000 330.090000 ;
        RECT 201.000000 325.910000 206.000000 326.090000 ;
        RECT 251.000000 305.910000 256.000000 306.090000 ;
        RECT 251.000000 269.910000 256.000000 270.090000 ;
        RECT 251.000000 273.910000 256.000000 274.090000 ;
        RECT 251.000000 277.910000 256.000000 278.090000 ;
        RECT 251.000000 281.910000 256.000000 282.090000 ;
        RECT 251.000000 285.910000 256.000000 286.090000 ;
        RECT 251.000000 293.910000 256.000000 294.090000 ;
        RECT 251.000000 289.910000 256.000000 290.090000 ;
        RECT 251.000000 301.910000 256.000000 302.090000 ;
        RECT 251.000000 297.910000 256.000000 298.090000 ;
        RECT 251.000000 309.910000 256.000000 310.090000 ;
        RECT 251.000000 313.910000 256.000000 314.090000 ;
        RECT 251.000000 321.910000 256.000000 322.090000 ;
        RECT 251.000000 317.910000 256.000000 318.090000 ;
        RECT 251.000000 329.910000 256.000000 330.090000 ;
        RECT 251.000000 325.910000 256.000000 326.090000 ;
        RECT 251.000000 333.910000 256.000000 334.090000 ;
        RECT 251.000000 337.910000 256.000000 338.090000 ;
        RECT 251.000000 341.910000 256.000000 342.090000 ;
        RECT 301.000000 265.910000 306.000000 266.090000 ;
        RECT 301.000000 261.910000 306.000000 262.090000 ;
        RECT 351.000000 265.910000 356.000000 266.090000 ;
        RECT 351.000000 261.910000 356.000000 262.090000 ;
        RECT 401.000000 265.910000 406.000000 266.090000 ;
        RECT 401.000000 261.910000 406.000000 262.090000 ;
        RECT 351.000000 305.910000 356.000000 306.090000 ;
        RECT 301.000000 305.910000 306.000000 306.090000 ;
        RECT 301.000000 277.910000 306.000000 278.090000 ;
        RECT 301.000000 269.910000 306.000000 270.090000 ;
        RECT 301.000000 273.910000 306.000000 274.090000 ;
        RECT 301.000000 281.910000 306.000000 282.090000 ;
        RECT 301.000000 285.910000 306.000000 286.090000 ;
        RECT 301.000000 293.910000 306.000000 294.090000 ;
        RECT 301.000000 289.910000 306.000000 290.090000 ;
        RECT 301.000000 301.910000 306.000000 302.090000 ;
        RECT 301.000000 297.910000 306.000000 298.090000 ;
        RECT 351.000000 269.910000 356.000000 270.090000 ;
        RECT 351.000000 273.910000 356.000000 274.090000 ;
        RECT 351.000000 277.910000 356.000000 278.090000 ;
        RECT 351.000000 281.910000 356.000000 282.090000 ;
        RECT 351.000000 285.910000 356.000000 286.090000 ;
        RECT 351.000000 301.910000 356.000000 302.090000 ;
        RECT 351.000000 297.910000 356.000000 298.090000 ;
        RECT 351.000000 293.910000 356.000000 294.090000 ;
        RECT 351.000000 289.910000 356.000000 290.090000 ;
        RECT 301.000000 313.910000 306.000000 314.090000 ;
        RECT 301.000000 309.910000 306.000000 310.090000 ;
        RECT 301.000000 317.910000 306.000000 318.090000 ;
        RECT 301.000000 321.910000 306.000000 322.090000 ;
        RECT 301.000000 329.910000 306.000000 330.090000 ;
        RECT 301.000000 325.910000 306.000000 326.090000 ;
        RECT 301.000000 341.910000 306.000000 342.090000 ;
        RECT 301.000000 337.910000 306.000000 338.090000 ;
        RECT 301.000000 333.910000 306.000000 334.090000 ;
        RECT 351.000000 313.910000 356.000000 314.090000 ;
        RECT 351.000000 309.910000 356.000000 310.090000 ;
        RECT 351.000000 317.910000 356.000000 318.090000 ;
        RECT 351.000000 321.910000 356.000000 322.090000 ;
        RECT 351.000000 341.910000 356.000000 342.090000 ;
        RECT 351.000000 337.910000 356.000000 338.090000 ;
        RECT 351.000000 333.910000 356.000000 334.090000 ;
        RECT 351.000000 329.910000 356.000000 330.090000 ;
        RECT 351.000000 325.910000 356.000000 326.090000 ;
        RECT 401.000000 305.910000 406.000000 306.090000 ;
        RECT 401.000000 269.910000 406.000000 270.090000 ;
        RECT 401.000000 273.910000 406.000000 274.090000 ;
        RECT 401.000000 277.910000 406.000000 278.090000 ;
        RECT 401.000000 281.910000 406.000000 282.090000 ;
        RECT 401.000000 285.910000 406.000000 286.090000 ;
        RECT 401.000000 293.910000 406.000000 294.090000 ;
        RECT 401.000000 289.910000 406.000000 290.090000 ;
        RECT 401.000000 297.910000 406.000000 298.090000 ;
        RECT 401.000000 301.910000 406.000000 302.090000 ;
        RECT 401.000000 309.910000 406.000000 310.090000 ;
        RECT 401.000000 313.910000 406.000000 314.090000 ;
        RECT 401.000000 317.910000 406.000000 318.090000 ;
        RECT 401.000000 321.910000 406.000000 322.090000 ;
        RECT 401.000000 325.910000 406.000000 326.090000 ;
        RECT 401.000000 329.910000 406.000000 330.090000 ;
        RECT 401.000000 333.910000 406.000000 334.090000 ;
        RECT 401.000000 337.910000 406.000000 338.090000 ;
        RECT 401.000000 341.910000 406.000000 342.090000 ;
        RECT 451.000000 261.910000 456.000000 262.090000 ;
        RECT 451.000000 265.910000 456.000000 266.090000 ;
        RECT 501.000000 261.910000 506.000000 262.090000 ;
        RECT 501.000000 265.910000 506.000000 266.090000 ;
        RECT 551.000000 265.910000 556.000000 266.090000 ;
        RECT 551.000000 261.910000 556.000000 262.090000 ;
        RECT 501.000000 305.910000 506.000000 306.090000 ;
        RECT 451.000000 273.910000 456.000000 274.090000 ;
        RECT 451.000000 269.910000 456.000000 270.090000 ;
        RECT 451.000000 277.910000 456.000000 278.090000 ;
        RECT 451.000000 285.910000 456.000000 286.090000 ;
        RECT 451.000000 281.910000 456.000000 282.090000 ;
        RECT 451.000000 293.910000 456.000000 294.090000 ;
        RECT 451.000000 289.910000 456.000000 290.090000 ;
        RECT 451.000000 297.910000 456.000000 298.090000 ;
        RECT 501.000000 277.910000 506.000000 278.090000 ;
        RECT 501.000000 273.910000 506.000000 274.090000 ;
        RECT 501.000000 269.910000 506.000000 270.090000 ;
        RECT 501.000000 281.910000 506.000000 282.090000 ;
        RECT 501.000000 285.910000 506.000000 286.090000 ;
        RECT 501.000000 289.910000 506.000000 290.090000 ;
        RECT 501.000000 293.910000 506.000000 294.090000 ;
        RECT 501.000000 301.910000 506.000000 302.090000 ;
        RECT 501.000000 297.910000 506.000000 298.090000 ;
        RECT 451.000000 321.910000 456.000000 322.090000 ;
        RECT 451.000000 316.105000 456.000000 317.105000 ;
        RECT 451.000000 333.910000 456.000000 334.090000 ;
        RECT 451.000000 329.910000 456.000000 330.090000 ;
        RECT 451.000000 325.910000 456.000000 326.090000 ;
        RECT 451.000000 337.910000 456.000000 338.090000 ;
        RECT 451.000000 341.910000 456.000000 342.090000 ;
        RECT 501.000000 313.910000 506.000000 314.090000 ;
        RECT 501.000000 309.910000 506.000000 310.090000 ;
        RECT 501.000000 317.910000 506.000000 318.090000 ;
        RECT 501.000000 321.910000 506.000000 322.090000 ;
        RECT 501.000000 329.910000 506.000000 330.090000 ;
        RECT 501.000000 325.910000 506.000000 326.090000 ;
        RECT 501.000000 333.910000 506.000000 334.090000 ;
        RECT 501.000000 337.910000 506.000000 338.090000 ;
        RECT 501.000000 341.910000 506.000000 342.090000 ;
        RECT 551.000000 305.910000 556.000000 306.090000 ;
        RECT 551.000000 285.910000 556.000000 286.090000 ;
        RECT 551.000000 281.910000 556.000000 282.090000 ;
        RECT 551.000000 277.910000 556.000000 278.090000 ;
        RECT 551.000000 273.910000 556.000000 274.090000 ;
        RECT 551.000000 269.910000 556.000000 270.090000 ;
        RECT 551.000000 301.910000 556.000000 302.090000 ;
        RECT 551.000000 297.910000 556.000000 298.090000 ;
        RECT 551.000000 293.910000 556.000000 294.090000 ;
        RECT 551.000000 289.910000 556.000000 290.090000 ;
        RECT 551.000000 313.910000 556.000000 314.090000 ;
        RECT 551.000000 309.910000 556.000000 310.090000 ;
        RECT 551.000000 321.910000 556.000000 322.090000 ;
        RECT 551.000000 317.910000 556.000000 318.090000 ;
        RECT 551.000000 325.910000 556.000000 326.090000 ;
        RECT 551.000000 329.910000 556.000000 330.090000 ;
        RECT 551.000000 333.910000 556.000000 334.090000 ;
        RECT 551.000000 337.910000 556.000000 338.090000 ;
        RECT 551.000000 341.910000 556.000000 342.090000 ;
        RECT 601.000000 1.910000 606.000000 2.090000 ;
        RECT 601.000000 5.910000 606.000000 6.090000 ;
        RECT 651.000000 1.910000 656.000000 2.090000 ;
        RECT 651.000000 5.910000 656.000000 6.090000 ;
        RECT 701.000000 1.910000 706.000000 2.090000 ;
        RECT 701.000000 5.910000 706.000000 6.090000 ;
        RECT 751.000000 1.910000 756.000000 2.090000 ;
        RECT 751.000000 5.910000 756.000000 6.090000 ;
        RECT 801.000000 1.910000 806.000000 2.090000 ;
        RECT 801.000000 5.910000 806.000000 6.090000 ;
        RECT 851.000000 1.910000 856.000000 2.090000 ;
        RECT 851.000000 5.910000 856.000000 6.090000 ;
        RECT 901.000000 1.910000 906.000000 2.090000 ;
        RECT 901.000000 5.910000 906.000000 6.090000 ;
        RECT 951.000000 1.910000 956.000000 2.090000 ;
        RECT 951.000000 5.910000 956.000000 6.090000 ;
        RECT 1001.000000 1.910000 1006.000000 2.090000 ;
        RECT 1001.000000 5.910000 1006.000000 6.090000 ;
        RECT 1051.000000 1.910000 1056.000000 2.090000 ;
        RECT 1051.000000 5.910000 1056.000000 6.090000 ;
        RECT 1101.000000 1.910000 1106.000000 2.090000 ;
        RECT 1101.000000 5.910000 1106.000000 6.090000 ;
        RECT 1151.000000 5.910000 1156.000000 6.090000 ;
        RECT 1172.000000 5.910000 1182.000000 6.090000 ;
        RECT 1151.000000 1.910000 1156.000000 2.090000 ;
        RECT 1172.000000 17.910000 1182.000000 18.090000 ;
        RECT 1172.000000 13.910000 1182.000000 14.090000 ;
        RECT 1172.000000 9.910000 1182.000000 10.090000 ;
        RECT 1172.000000 21.910000 1182.000000 22.090000 ;
        RECT 1172.000000 25.910000 1182.000000 26.090000 ;
        RECT 1172.000000 33.910000 1182.000000 34.090000 ;
        RECT 1172.000000 29.910000 1182.000000 30.090000 ;
        RECT 1172.000000 41.910000 1182.000000 42.090000 ;
        RECT 1172.000000 37.910000 1182.000000 38.090000 ;
        RECT 1172.000000 45.910000 1182.000000 46.090000 ;
        RECT 601.000000 265.910000 606.000000 266.090000 ;
        RECT 601.000000 261.910000 606.000000 262.090000 ;
        RECT 651.000000 261.910000 656.000000 262.090000 ;
        RECT 651.000000 265.910000 656.000000 266.090000 ;
        RECT 701.000000 265.910000 706.000000 266.090000 ;
        RECT 701.000000 261.910000 706.000000 262.090000 ;
        RECT 601.000000 305.910000 606.000000 306.090000 ;
        RECT 651.000000 305.910000 656.000000 306.090000 ;
        RECT 601.000000 269.910000 606.000000 270.090000 ;
        RECT 601.000000 273.910000 606.000000 274.090000 ;
        RECT 601.000000 277.910000 606.000000 278.090000 ;
        RECT 601.000000 281.910000 606.000000 282.090000 ;
        RECT 601.000000 285.910000 606.000000 286.090000 ;
        RECT 601.000000 293.910000 606.000000 294.090000 ;
        RECT 601.000000 289.910000 606.000000 290.090000 ;
        RECT 601.000000 301.910000 606.000000 302.090000 ;
        RECT 601.000000 297.910000 606.000000 298.090000 ;
        RECT 651.000000 269.910000 656.000000 270.090000 ;
        RECT 651.000000 273.910000 656.000000 274.090000 ;
        RECT 651.000000 277.910000 656.000000 278.090000 ;
        RECT 651.000000 281.910000 656.000000 282.090000 ;
        RECT 651.000000 285.910000 656.000000 286.090000 ;
        RECT 651.000000 289.910000 656.000000 290.090000 ;
        RECT 651.000000 293.910000 656.000000 294.090000 ;
        RECT 651.000000 297.910000 656.000000 298.090000 ;
        RECT 651.000000 301.910000 656.000000 302.090000 ;
        RECT 601.000000 313.910000 606.000000 314.090000 ;
        RECT 601.000000 309.910000 606.000000 310.090000 ;
        RECT 601.000000 317.910000 606.000000 318.090000 ;
        RECT 601.000000 321.910000 606.000000 322.090000 ;
        RECT 601.000000 325.910000 606.000000 326.090000 ;
        RECT 601.000000 329.910000 606.000000 330.090000 ;
        RECT 601.000000 333.910000 606.000000 334.090000 ;
        RECT 601.000000 337.910000 606.000000 338.090000 ;
        RECT 601.000000 341.910000 606.000000 342.090000 ;
        RECT 651.000000 313.910000 656.000000 314.090000 ;
        RECT 651.000000 309.910000 656.000000 310.090000 ;
        RECT 651.000000 321.910000 656.000000 322.090000 ;
        RECT 651.000000 317.910000 656.000000 318.090000 ;
        RECT 651.000000 329.910000 656.000000 330.090000 ;
        RECT 651.000000 325.910000 656.000000 326.090000 ;
        RECT 651.000000 333.910000 656.000000 334.090000 ;
        RECT 651.000000 337.910000 656.000000 338.090000 ;
        RECT 651.000000 341.910000 656.000000 342.090000 ;
        RECT 701.000000 305.910000 706.000000 306.090000 ;
        RECT 701.000000 285.910000 706.000000 286.090000 ;
        RECT 701.000000 281.910000 706.000000 282.090000 ;
        RECT 701.000000 277.910000 706.000000 278.090000 ;
        RECT 701.000000 273.910000 706.000000 274.090000 ;
        RECT 701.000000 269.910000 706.000000 270.090000 ;
        RECT 701.000000 301.910000 706.000000 302.090000 ;
        RECT 701.000000 297.910000 706.000000 298.090000 ;
        RECT 701.000000 293.910000 706.000000 294.090000 ;
        RECT 701.000000 289.910000 706.000000 290.090000 ;
        RECT 701.000000 309.910000 706.000000 310.090000 ;
        RECT 701.000000 313.910000 706.000000 314.090000 ;
        RECT 701.000000 317.910000 706.000000 318.090000 ;
        RECT 701.000000 321.910000 706.000000 322.090000 ;
        RECT 701.000000 325.910000 706.000000 326.090000 ;
        RECT 701.000000 329.910000 706.000000 330.090000 ;
        RECT 701.000000 333.910000 706.000000 334.090000 ;
        RECT 701.000000 337.910000 706.000000 338.090000 ;
        RECT 701.000000 341.910000 706.000000 342.090000 ;
        RECT 751.000000 261.910000 756.000000 262.090000 ;
        RECT 751.000000 265.910000 756.000000 266.090000 ;
        RECT 801.000000 261.910000 806.000000 262.090000 ;
        RECT 801.000000 265.910000 806.000000 266.090000 ;
        RECT 851.000000 265.910000 856.000000 266.090000 ;
        RECT 851.000000 261.910000 856.000000 262.090000 ;
        RECT 801.000000 305.910000 806.000000 306.090000 ;
        RECT 751.000000 305.910000 756.000000 306.090000 ;
        RECT 751.000000 285.910000 756.000000 286.090000 ;
        RECT 751.000000 281.910000 756.000000 282.090000 ;
        RECT 751.000000 269.910000 756.000000 270.090000 ;
        RECT 751.000000 273.910000 756.000000 274.090000 ;
        RECT 751.000000 277.910000 756.000000 278.090000 ;
        RECT 751.000000 289.910000 756.000000 290.090000 ;
        RECT 751.000000 293.910000 756.000000 294.090000 ;
        RECT 751.000000 297.910000 756.000000 298.090000 ;
        RECT 751.000000 301.910000 756.000000 302.090000 ;
        RECT 801.000000 277.910000 806.000000 278.090000 ;
        RECT 801.000000 273.910000 806.000000 274.090000 ;
        RECT 801.000000 269.910000 806.000000 270.090000 ;
        RECT 801.000000 281.910000 806.000000 282.090000 ;
        RECT 801.000000 285.910000 806.000000 286.090000 ;
        RECT 801.000000 289.910000 806.000000 290.090000 ;
        RECT 801.000000 293.910000 806.000000 294.090000 ;
        RECT 801.000000 301.910000 806.000000 302.090000 ;
        RECT 801.000000 297.910000 806.000000 298.090000 ;
        RECT 751.000000 321.910000 756.000000 322.090000 ;
        RECT 751.000000 309.910000 756.000000 310.090000 ;
        RECT 751.000000 313.910000 756.000000 314.090000 ;
        RECT 751.000000 317.910000 756.000000 318.090000 ;
        RECT 751.000000 329.910000 756.000000 330.090000 ;
        RECT 751.000000 325.910000 756.000000 326.090000 ;
        RECT 751.000000 341.910000 756.000000 342.090000 ;
        RECT 751.000000 337.910000 756.000000 338.090000 ;
        RECT 751.000000 333.910000 756.000000 334.090000 ;
        RECT 801.000000 309.910000 806.000000 310.090000 ;
        RECT 801.000000 313.910000 806.000000 314.090000 ;
        RECT 801.000000 321.910000 806.000000 322.090000 ;
        RECT 801.000000 317.910000 806.000000 318.090000 ;
        RECT 801.000000 325.910000 806.000000 326.090000 ;
        RECT 801.000000 329.910000 806.000000 330.090000 ;
        RECT 801.000000 337.910000 806.000000 338.090000 ;
        RECT 801.000000 333.910000 806.000000 334.090000 ;
        RECT 801.000000 341.910000 806.000000 342.090000 ;
        RECT 851.000000 305.910000 856.000000 306.090000 ;
        RECT 851.000000 285.910000 856.000000 286.090000 ;
        RECT 851.000000 281.910000 856.000000 282.090000 ;
        RECT 851.000000 277.910000 856.000000 278.090000 ;
        RECT 851.000000 273.910000 856.000000 274.090000 ;
        RECT 851.000000 269.910000 856.000000 270.090000 ;
        RECT 851.000000 301.910000 856.000000 302.090000 ;
        RECT 851.000000 297.910000 856.000000 298.090000 ;
        RECT 851.000000 293.910000 856.000000 294.090000 ;
        RECT 851.000000 289.910000 856.000000 290.090000 ;
        RECT 851.000000 309.910000 856.000000 310.090000 ;
        RECT 851.000000 313.910000 856.000000 314.090000 ;
        RECT 851.000000 317.910000 856.000000 318.090000 ;
        RECT 851.000000 321.910000 856.000000 322.090000 ;
        RECT 851.000000 325.910000 856.000000 326.090000 ;
        RECT 851.000000 329.910000 856.000000 330.090000 ;
        RECT 851.000000 333.910000 856.000000 334.090000 ;
        RECT 851.000000 337.910000 856.000000 338.090000 ;
        RECT 851.000000 341.910000 856.000000 342.090000 ;
        RECT 1172.000000 61.910000 1182.000000 62.090000 ;
        RECT 1172.000000 57.910000 1182.000000 58.090000 ;
        RECT 1172.000000 53.910000 1182.000000 54.090000 ;
        RECT 1172.000000 49.910000 1182.000000 50.090000 ;
        RECT 1172.000000 73.910000 1182.000000 74.090000 ;
        RECT 1172.000000 69.910000 1182.000000 70.090000 ;
        RECT 1172.000000 65.910000 1182.000000 66.090000 ;
        RECT 1172.000000 77.910000 1182.000000 78.090000 ;
        RECT 1172.000000 81.910000 1182.000000 82.090000 ;
        RECT 1172.000000 89.910000 1182.000000 90.090000 ;
        RECT 1172.000000 85.910000 1182.000000 86.090000 ;
        RECT 1172.000000 97.910000 1182.000000 98.090000 ;
        RECT 1172.000000 93.910000 1182.000000 94.090000 ;
        RECT 1172.000000 101.910000 1182.000000 102.090000 ;
        RECT 1172.000000 117.910000 1182.000000 118.090000 ;
        RECT 1172.000000 113.910000 1182.000000 114.090000 ;
        RECT 1172.000000 105.910000 1182.000000 106.090000 ;
        RECT 1172.000000 109.910000 1182.000000 110.090000 ;
        RECT 1151.000000 133.910000 1156.000000 134.090000 ;
        RECT 1172.000000 125.910000 1182.000000 126.090000 ;
        RECT 1172.000000 121.910000 1182.000000 122.090000 ;
        RECT 1172.000000 129.910000 1182.000000 130.090000 ;
        RECT 1172.000000 133.910000 1182.000000 134.090000 ;
        RECT 1172.000000 137.910000 1182.000000 138.090000 ;
        RECT 1172.000000 141.910000 1182.000000 142.090000 ;
        RECT 1172.000000 145.910000 1182.000000 146.090000 ;
        RECT 1172.000000 149.910000 1182.000000 150.090000 ;
        RECT 1172.000000 153.910000 1182.000000 154.090000 ;
        RECT 1172.000000 165.910000 1182.000000 166.090000 ;
        RECT 1172.000000 161.910000 1182.000000 162.090000 ;
        RECT 1172.000000 157.910000 1182.000000 158.090000 ;
        RECT 1172.000000 169.910000 1182.000000 170.090000 ;
        RECT 1172.000000 173.910000 1182.000000 174.090000 ;
        RECT 1172.000000 177.910000 1182.000000 178.090000 ;
        RECT 1172.000000 181.910000 1182.000000 182.090000 ;
        RECT 1172.000000 185.910000 1182.000000 186.090000 ;
        RECT 1172.000000 189.910000 1182.000000 190.090000 ;
        RECT 1172.000000 193.910000 1182.000000 194.090000 ;
        RECT 901.000000 261.910000 906.000000 262.090000 ;
        RECT 901.000000 265.910000 906.000000 266.090000 ;
        RECT 951.000000 265.910000 956.000000 266.090000 ;
        RECT 951.000000 261.910000 956.000000 262.090000 ;
        RECT 1001.000000 261.910000 1006.000000 262.090000 ;
        RECT 1001.000000 265.910000 1006.000000 266.090000 ;
        RECT 951.000000 305.910000 956.000000 306.090000 ;
        RECT 901.000000 305.910000 906.000000 306.090000 ;
        RECT 901.000000 285.910000 906.000000 286.090000 ;
        RECT 901.000000 281.910000 906.000000 282.090000 ;
        RECT 901.000000 269.910000 906.000000 270.090000 ;
        RECT 901.000000 273.910000 906.000000 274.090000 ;
        RECT 901.000000 277.910000 906.000000 278.090000 ;
        RECT 901.000000 289.910000 906.000000 290.090000 ;
        RECT 901.000000 293.910000 906.000000 294.090000 ;
        RECT 901.000000 297.910000 906.000000 298.090000 ;
        RECT 901.000000 301.910000 906.000000 302.090000 ;
        RECT 951.000000 269.910000 956.000000 270.090000 ;
        RECT 951.000000 273.910000 956.000000 274.090000 ;
        RECT 951.000000 277.910000 956.000000 278.090000 ;
        RECT 951.000000 281.910000 956.000000 282.090000 ;
        RECT 951.000000 285.910000 956.000000 286.090000 ;
        RECT 951.000000 301.910000 956.000000 302.090000 ;
        RECT 951.000000 297.910000 956.000000 298.090000 ;
        RECT 951.000000 293.910000 956.000000 294.090000 ;
        RECT 951.000000 289.910000 956.000000 290.090000 ;
        RECT 901.000000 321.910000 906.000000 322.090000 ;
        RECT 901.000000 309.910000 906.000000 310.090000 ;
        RECT 901.000000 313.910000 906.000000 314.090000 ;
        RECT 901.000000 317.910000 906.000000 318.090000 ;
        RECT 901.000000 325.910000 906.000000 326.090000 ;
        RECT 901.000000 329.910000 906.000000 330.090000 ;
        RECT 901.000000 333.910000 906.000000 334.090000 ;
        RECT 901.000000 337.910000 906.000000 338.090000 ;
        RECT 901.000000 341.910000 906.000000 342.090000 ;
        RECT 951.000000 313.910000 956.000000 314.090000 ;
        RECT 951.000000 309.910000 956.000000 310.090000 ;
        RECT 951.000000 317.910000 956.000000 318.090000 ;
        RECT 951.000000 321.910000 956.000000 322.090000 ;
        RECT 951.000000 325.910000 956.000000 326.090000 ;
        RECT 951.000000 329.910000 956.000000 330.090000 ;
        RECT 951.000000 333.910000 956.000000 334.090000 ;
        RECT 951.000000 337.910000 956.000000 338.090000 ;
        RECT 951.000000 341.910000 956.000000 342.090000 ;
        RECT 1001.000000 305.910000 1006.000000 306.090000 ;
        RECT 1001.000000 277.910000 1006.000000 278.090000 ;
        RECT 1001.000000 273.910000 1006.000000 274.090000 ;
        RECT 1001.000000 269.910000 1006.000000 270.090000 ;
        RECT 1001.000000 281.910000 1006.000000 282.090000 ;
        RECT 1001.000000 285.910000 1006.000000 286.090000 ;
        RECT 1001.000000 289.910000 1006.000000 290.090000 ;
        RECT 1001.000000 293.910000 1006.000000 294.090000 ;
        RECT 1001.000000 301.910000 1006.000000 302.090000 ;
        RECT 1001.000000 297.910000 1006.000000 298.090000 ;
        RECT 1001.000000 313.910000 1006.000000 314.090000 ;
        RECT 1001.000000 309.910000 1006.000000 310.090000 ;
        RECT 1001.000000 317.910000 1006.000000 318.090000 ;
        RECT 1001.000000 321.910000 1006.000000 322.090000 ;
        RECT 1001.000000 329.910000 1006.000000 330.090000 ;
        RECT 1001.000000 325.910000 1006.000000 326.090000 ;
        RECT 1001.000000 333.910000 1006.000000 334.090000 ;
        RECT 1001.000000 337.910000 1006.000000 338.090000 ;
        RECT 1001.000000 341.910000 1006.000000 342.090000 ;
        RECT 1051.000000 261.910000 1056.000000 262.090000 ;
        RECT 1051.000000 265.910000 1056.000000 266.090000 ;
        RECT 1101.000000 265.910000 1106.000000 266.090000 ;
        RECT 1101.000000 261.910000 1106.000000 262.090000 ;
        RECT 1172.000000 197.910000 1182.000000 198.090000 ;
        RECT 1172.000000 201.910000 1182.000000 202.090000 ;
        RECT 1172.000000 205.910000 1182.000000 206.090000 ;
        RECT 1172.000000 209.910000 1182.000000 210.090000 ;
        RECT 1172.000000 221.910000 1182.000000 222.090000 ;
        RECT 1172.000000 217.910000 1182.000000 218.090000 ;
        RECT 1172.000000 213.910000 1182.000000 214.090000 ;
        RECT 1172.000000 225.910000 1182.000000 226.090000 ;
        RECT 1172.000000 229.910000 1182.000000 230.090000 ;
        RECT 1172.000000 237.910000 1182.000000 238.090000 ;
        RECT 1172.000000 233.910000 1182.000000 234.090000 ;
        RECT 1172.000000 241.910000 1182.000000 242.090000 ;
        RECT 1172.000000 245.910000 1182.000000 246.090000 ;
        RECT 1172.000000 249.910000 1182.000000 250.090000 ;
        RECT 1151.000000 257.910000 1156.000000 258.090000 ;
        RECT 1151.000000 265.910000 1156.000000 266.090000 ;
        RECT 1151.000000 261.910000 1156.000000 262.090000 ;
        RECT 1172.000000 265.910000 1182.000000 266.090000 ;
        RECT 1172.000000 253.910000 1182.000000 254.090000 ;
        RECT 1172.000000 257.910000 1182.000000 258.090000 ;
        RECT 1172.000000 261.910000 1182.000000 262.090000 ;
        RECT 1101.000000 305.910000 1106.000000 306.090000 ;
        RECT 1051.000000 305.910000 1056.000000 306.090000 ;
        RECT 1051.000000 285.910000 1056.000000 286.090000 ;
        RECT 1051.000000 281.910000 1056.000000 282.090000 ;
        RECT 1051.000000 273.910000 1056.000000 274.090000 ;
        RECT 1051.000000 269.910000 1056.000000 270.090000 ;
        RECT 1051.000000 277.910000 1056.000000 278.090000 ;
        RECT 1051.000000 289.910000 1056.000000 290.090000 ;
        RECT 1051.000000 293.910000 1056.000000 294.090000 ;
        RECT 1051.000000 297.910000 1056.000000 298.090000 ;
        RECT 1051.000000 301.910000 1056.000000 302.090000 ;
        RECT 1101.000000 269.910000 1106.000000 270.090000 ;
        RECT 1101.000000 273.910000 1106.000000 274.090000 ;
        RECT 1101.000000 277.910000 1106.000000 278.090000 ;
        RECT 1101.000000 281.910000 1106.000000 282.090000 ;
        RECT 1101.000000 285.910000 1106.000000 286.090000 ;
        RECT 1101.000000 301.910000 1106.000000 302.090000 ;
        RECT 1101.000000 297.910000 1106.000000 298.090000 ;
        RECT 1101.000000 293.910000 1106.000000 294.090000 ;
        RECT 1101.000000 289.910000 1106.000000 290.090000 ;
        RECT 1051.000000 321.910000 1056.000000 322.090000 ;
        RECT 1051.000000 309.910000 1056.000000 310.090000 ;
        RECT 1051.000000 313.910000 1056.000000 314.090000 ;
        RECT 1051.000000 317.910000 1056.000000 318.090000 ;
        RECT 1051.000000 325.910000 1056.000000 326.090000 ;
        RECT 1051.000000 329.910000 1056.000000 330.090000 ;
        RECT 1051.000000 333.910000 1056.000000 334.090000 ;
        RECT 1051.000000 337.910000 1056.000000 338.090000 ;
        RECT 1051.000000 341.910000 1056.000000 342.090000 ;
        RECT 1101.000000 313.910000 1106.000000 314.090000 ;
        RECT 1101.000000 309.910000 1106.000000 310.090000 ;
        RECT 1101.000000 317.910000 1106.000000 318.090000 ;
        RECT 1101.000000 321.910000 1106.000000 322.090000 ;
        RECT 1101.000000 325.910000 1106.000000 326.090000 ;
        RECT 1101.000000 329.910000 1106.000000 330.090000 ;
        RECT 1101.000000 333.910000 1106.000000 334.090000 ;
        RECT 1101.000000 337.910000 1106.000000 338.090000 ;
        RECT 1101.000000 341.910000 1106.000000 342.090000 ;
        RECT 1151.000000 305.910000 1156.000000 306.090000 ;
        RECT 1172.000000 305.910000 1182.000000 306.090000 ;
        RECT 1151.000000 269.910000 1156.000000 270.090000 ;
        RECT 1151.000000 273.910000 1156.000000 274.090000 ;
        RECT 1151.000000 277.910000 1156.000000 278.090000 ;
        RECT 1151.000000 281.910000 1156.000000 282.090000 ;
        RECT 1151.000000 285.910000 1156.000000 286.090000 ;
        RECT 1172.000000 277.910000 1182.000000 278.090000 ;
        RECT 1172.000000 269.910000 1182.000000 270.090000 ;
        RECT 1172.000000 273.910000 1182.000000 274.090000 ;
        RECT 1172.000000 281.910000 1182.000000 282.090000 ;
        RECT 1172.000000 285.910000 1182.000000 286.090000 ;
        RECT 1151.000000 301.910000 1156.000000 302.090000 ;
        RECT 1151.000000 297.910000 1156.000000 298.090000 ;
        RECT 1151.000000 289.910000 1156.000000 290.090000 ;
        RECT 1151.000000 293.910000 1156.000000 294.090000 ;
        RECT 1172.000000 301.910000 1182.000000 302.090000 ;
        RECT 1172.000000 289.910000 1182.000000 290.090000 ;
        RECT 1172.000000 293.910000 1182.000000 294.090000 ;
        RECT 1172.000000 297.910000 1182.000000 298.090000 ;
        RECT 1151.000000 321.910000 1156.000000 322.090000 ;
        RECT 1151.000000 317.910000 1156.000000 318.090000 ;
        RECT 1151.000000 309.910000 1156.000000 310.090000 ;
        RECT 1151.000000 313.910000 1156.000000 314.090000 ;
        RECT 1172.000000 321.910000 1182.000000 322.090000 ;
        RECT 1172.000000 309.910000 1182.000000 310.090000 ;
        RECT 1172.000000 313.910000 1182.000000 314.090000 ;
        RECT 1172.000000 317.910000 1182.000000 318.090000 ;
        RECT 1151.000000 329.910000 1156.000000 330.090000 ;
        RECT 1151.000000 325.910000 1156.000000 326.090000 ;
        RECT 1151.000000 333.910000 1156.000000 334.090000 ;
        RECT 1151.000000 337.910000 1156.000000 338.090000 ;
        RECT 1151.000000 341.910000 1156.000000 342.090000 ;
        RECT 1172.000000 329.910000 1182.000000 330.090000 ;
        RECT 1172.000000 325.910000 1182.000000 326.090000 ;
        RECT 1172.000000 333.910000 1182.000000 334.090000 ;
        RECT 1172.000000 337.910000 1182.000000 338.090000 ;
        RECT 1172.000000 341.910000 1182.000000 342.090000 ;
        RECT 4.000000 357.910000 14.000000 358.090000 ;
        RECT 4.000000 353.910000 14.000000 354.090000 ;
        RECT 4.000000 345.910000 14.000000 346.090000 ;
        RECT 4.000000 349.910000 14.000000 350.090000 ;
        RECT 4.000000 369.910000 14.000000 370.090000 ;
        RECT 4.000000 365.910000 14.000000 366.090000 ;
        RECT 4.000000 361.910000 14.000000 362.090000 ;
        RECT 4.000000 377.910000 14.000000 378.090000 ;
        RECT 4.000000 373.910000 14.000000 374.090000 ;
        RECT 51.000000 354.445000 56.000000 354.745000 ;
        RECT 51.000000 345.910000 56.000000 346.090000 ;
        RECT 51.000000 369.910000 56.000000 370.090000 ;
        RECT 51.000000 365.910000 56.000000 366.090000 ;
        RECT 51.000000 361.910000 56.000000 362.090000 ;
        RECT 51.000000 373.910000 56.000000 374.090000 ;
        RECT 51.000000 377.910000 56.000000 378.090000 ;
        RECT 4.000000 397.910000 14.000000 398.090000 ;
        RECT 4.000000 393.910000 14.000000 394.090000 ;
        RECT 4.000000 389.910000 14.000000 390.090000 ;
        RECT 4.000000 381.910000 14.000000 382.090000 ;
        RECT 4.000000 385.910000 14.000000 386.090000 ;
        RECT 4.000000 401.910000 14.000000 402.090000 ;
        RECT 4.000000 405.910000 14.000000 406.090000 ;
        RECT 4.000000 409.910000 14.000000 410.090000 ;
        RECT 4.000000 413.910000 14.000000 414.090000 ;
        RECT 51.000000 385.910000 56.000000 386.090000 ;
        RECT 51.000000 381.910000 56.000000 382.090000 ;
        RECT 51.000000 389.910000 56.000000 390.090000 ;
        RECT 51.000000 393.910000 56.000000 394.090000 ;
        RECT 51.000000 397.910000 56.000000 398.090000 ;
        RECT 51.000000 413.910000 56.000000 414.090000 ;
        RECT 51.000000 409.910000 56.000000 410.090000 ;
        RECT 51.000000 405.910000 56.000000 406.090000 ;
        RECT 51.000000 401.910000 56.000000 402.090000 ;
        RECT 101.000000 345.910000 106.000000 346.090000 ;
        RECT 101.000000 349.910000 106.000000 350.090000 ;
        RECT 101.000000 353.910000 106.000000 354.090000 ;
        RECT 101.000000 357.910000 106.000000 358.090000 ;
        RECT 101.000000 361.910000 106.000000 362.090000 ;
        RECT 101.000000 365.910000 106.000000 366.090000 ;
        RECT 101.000000 369.910000 106.000000 370.090000 ;
        RECT 101.000000 373.910000 106.000000 374.090000 ;
        RECT 101.000000 377.910000 106.000000 378.090000 ;
        RECT 101.000000 381.910000 106.000000 382.090000 ;
        RECT 101.000000 385.910000 106.000000 386.090000 ;
        RECT 101.000000 389.910000 106.000000 390.090000 ;
        RECT 101.000000 393.910000 106.000000 394.090000 ;
        RECT 101.000000 397.910000 106.000000 398.090000 ;
        RECT 101.000000 413.910000 106.000000 414.090000 ;
        RECT 101.000000 409.910000 106.000000 410.090000 ;
        RECT 101.000000 405.910000 106.000000 406.090000 ;
        RECT 101.000000 401.910000 106.000000 402.090000 ;
        RECT 4.000000 433.910000 14.000000 434.090000 ;
        RECT 4.000000 429.910000 14.000000 430.090000 ;
        RECT 4.000000 417.910000 14.000000 418.090000 ;
        RECT 4.000000 421.910000 14.000000 422.090000 ;
        RECT 4.000000 425.910000 14.000000 426.090000 ;
        RECT 4.000000 437.910000 14.000000 438.090000 ;
        RECT 4.000000 441.910000 14.000000 442.090000 ;
        RECT 4.000000 445.910000 14.000000 446.090000 ;
        RECT 4.000000 449.910000 14.000000 450.090000 ;
        RECT 4.000000 453.910000 14.000000 454.090000 ;
        RECT 51.000000 417.910000 56.000000 418.090000 ;
        RECT 51.000000 421.910000 56.000000 422.090000 ;
        RECT 51.000000 425.910000 56.000000 426.090000 ;
        RECT 51.000000 429.910000 56.000000 430.090000 ;
        RECT 51.000000 433.910000 56.000000 434.090000 ;
        RECT 51.000000 453.910000 56.000000 454.090000 ;
        RECT 51.000000 449.910000 56.000000 450.090000 ;
        RECT 51.000000 445.910000 56.000000 446.090000 ;
        RECT 51.000000 441.910000 56.000000 442.090000 ;
        RECT 51.000000 437.910000 56.000000 438.090000 ;
        RECT 4.000000 469.910000 14.000000 470.090000 ;
        RECT 4.000000 457.910000 14.000000 458.090000 ;
        RECT 4.000000 461.910000 14.000000 462.090000 ;
        RECT 4.000000 465.910000 14.000000 466.090000 ;
        RECT 4.000000 473.910000 14.000000 474.090000 ;
        RECT 4.000000 477.910000 14.000000 478.090000 ;
        RECT 4.000000 481.910000 14.000000 482.090000 ;
        RECT 4.000000 485.910000 14.000000 486.090000 ;
        RECT 4.000000 489.910000 14.000000 490.090000 ;
        RECT 51.000000 461.910000 56.000000 462.090000 ;
        RECT 51.000000 457.910000 56.000000 458.090000 ;
        RECT 51.000000 465.910000 56.000000 466.090000 ;
        RECT 51.000000 469.910000 56.000000 470.090000 ;
        RECT 51.000000 489.910000 56.000000 490.090000 ;
        RECT 51.000000 485.910000 56.000000 486.090000 ;
        RECT 51.000000 481.910000 56.000000 482.090000 ;
        RECT 51.000000 477.910000 56.000000 478.090000 ;
        RECT 51.000000 473.910000 56.000000 474.090000 ;
        RECT 101.000000 417.910000 106.000000 418.090000 ;
        RECT 101.000000 421.910000 106.000000 422.090000 ;
        RECT 101.000000 425.910000 106.000000 426.090000 ;
        RECT 101.000000 429.910000 106.000000 430.090000 ;
        RECT 101.000000 433.910000 106.000000 434.090000 ;
        RECT 101.000000 437.910000 106.000000 438.090000 ;
        RECT 101.000000 441.910000 106.000000 442.090000 ;
        RECT 101.000000 445.910000 106.000000 446.090000 ;
        RECT 101.000000 449.910000 106.000000 450.090000 ;
        RECT 101.000000 453.910000 106.000000 454.090000 ;
        RECT 101.000000 469.910000 106.000000 470.090000 ;
        RECT 101.000000 465.910000 106.000000 466.090000 ;
        RECT 101.000000 461.910000 106.000000 462.090000 ;
        RECT 101.000000 457.910000 106.000000 458.090000 ;
        RECT 101.000000 473.910000 106.000000 474.090000 ;
        RECT 101.000000 477.910000 106.000000 478.090000 ;
        RECT 101.000000 481.910000 106.000000 482.090000 ;
        RECT 101.000000 485.910000 106.000000 486.090000 ;
        RECT 101.000000 489.910000 106.000000 490.090000 ;
        RECT 151.000000 349.910000 156.000000 350.090000 ;
        RECT 151.000000 345.910000 156.000000 346.090000 ;
        RECT 151.000000 353.910000 156.000000 354.090000 ;
        RECT 151.000000 357.910000 156.000000 358.090000 ;
        RECT 151.000000 361.910000 156.000000 362.090000 ;
        RECT 151.000000 365.910000 156.000000 366.090000 ;
        RECT 151.000000 369.910000 156.000000 370.090000 ;
        RECT 151.000000 373.910000 156.000000 374.090000 ;
        RECT 151.000000 377.910000 156.000000 378.090000 ;
        RECT 201.000000 349.910000 206.000000 350.090000 ;
        RECT 201.000000 345.910000 206.000000 346.090000 ;
        RECT 201.000000 353.910000 206.000000 354.090000 ;
        RECT 201.000000 357.910000 206.000000 358.090000 ;
        RECT 201.000000 377.910000 206.000000 378.090000 ;
        RECT 201.000000 373.910000 206.000000 374.090000 ;
        RECT 201.000000 369.910000 206.000000 370.090000 ;
        RECT 201.000000 365.910000 206.000000 366.090000 ;
        RECT 201.000000 361.910000 206.000000 362.090000 ;
        RECT 151.000000 381.910000 156.000000 382.090000 ;
        RECT 151.000000 385.910000 156.000000 386.090000 ;
        RECT 151.000000 393.910000 156.000000 394.090000 ;
        RECT 151.000000 389.910000 156.000000 390.090000 ;
        RECT 151.000000 397.910000 156.000000 398.090000 ;
        RECT 151.000000 405.910000 156.000000 406.090000 ;
        RECT 151.000000 401.910000 156.000000 402.090000 ;
        RECT 201.000000 381.910000 206.000000 382.090000 ;
        RECT 201.000000 385.910000 206.000000 386.090000 ;
        RECT 201.000000 397.910000 206.000000 398.090000 ;
        RECT 201.000000 393.910000 206.000000 394.090000 ;
        RECT 201.000000 389.910000 206.000000 390.090000 ;
        RECT 201.000000 413.910000 206.000000 414.090000 ;
        RECT 201.000000 409.910000 206.000000 410.090000 ;
        RECT 201.000000 405.910000 206.000000 406.090000 ;
        RECT 201.000000 401.910000 206.000000 402.090000 ;
        RECT 251.000000 349.910000 256.000000 350.090000 ;
        RECT 251.000000 345.910000 256.000000 346.090000 ;
        RECT 251.000000 353.910000 256.000000 354.090000 ;
        RECT 251.000000 357.910000 256.000000 358.090000 ;
        RECT 251.000000 361.910000 256.000000 362.090000 ;
        RECT 251.000000 365.910000 256.000000 366.090000 ;
        RECT 251.000000 369.910000 256.000000 370.090000 ;
        RECT 251.000000 373.910000 256.000000 374.090000 ;
        RECT 251.000000 377.910000 256.000000 378.090000 ;
        RECT 251.000000 381.910000 256.000000 382.090000 ;
        RECT 251.000000 385.910000 256.000000 386.090000 ;
        RECT 251.000000 393.910000 256.000000 394.090000 ;
        RECT 251.000000 389.910000 256.000000 390.090000 ;
        RECT 251.000000 397.910000 256.000000 398.090000 ;
        RECT 251.000000 401.910000 256.000000 402.090000 ;
        RECT 251.000000 405.910000 256.000000 406.090000 ;
        RECT 151.000000 453.910000 156.000000 454.090000 ;
        RECT 201.000000 425.910000 206.000000 426.090000 ;
        RECT 201.000000 421.910000 206.000000 422.090000 ;
        RECT 201.000000 417.910000 206.000000 418.090000 ;
        RECT 201.000000 429.910000 206.000000 430.090000 ;
        RECT 201.000000 433.910000 206.000000 434.090000 ;
        RECT 201.000000 453.910000 206.000000 454.090000 ;
        RECT 201.000000 449.910000 206.000000 450.090000 ;
        RECT 201.000000 445.910000 206.000000 446.090000 ;
        RECT 201.000000 441.910000 206.000000 442.090000 ;
        RECT 201.000000 437.910000 206.000000 438.090000 ;
        RECT 151.000000 461.910000 156.000000 462.090000 ;
        RECT 151.000000 457.910000 156.000000 458.090000 ;
        RECT 151.000000 469.910000 156.000000 470.090000 ;
        RECT 151.000000 465.910000 156.000000 466.090000 ;
        RECT 151.000000 481.910000 156.000000 482.090000 ;
        RECT 151.000000 477.910000 156.000000 478.090000 ;
        RECT 151.000000 473.910000 156.000000 474.090000 ;
        RECT 151.000000 489.910000 156.000000 490.090000 ;
        RECT 151.000000 485.910000 156.000000 486.090000 ;
        RECT 201.000000 461.910000 206.000000 462.090000 ;
        RECT 201.000000 457.910000 206.000000 458.090000 ;
        RECT 201.000000 465.910000 206.000000 466.090000 ;
        RECT 201.000000 469.910000 206.000000 470.090000 ;
        RECT 201.000000 489.910000 206.000000 490.090000 ;
        RECT 201.000000 485.910000 206.000000 486.090000 ;
        RECT 201.000000 481.910000 206.000000 482.090000 ;
        RECT 201.000000 477.910000 206.000000 478.090000 ;
        RECT 201.000000 473.910000 206.000000 474.090000 ;
        RECT 251.000000 453.910000 256.000000 454.090000 ;
        RECT 251.000000 461.910000 256.000000 462.090000 ;
        RECT 251.000000 457.910000 256.000000 458.090000 ;
        RECT 251.000000 465.910000 256.000000 466.090000 ;
        RECT 251.000000 469.910000 256.000000 470.090000 ;
        RECT 251.000000 481.910000 256.000000 482.090000 ;
        RECT 251.000000 473.910000 256.000000 474.090000 ;
        RECT 251.000000 477.910000 256.000000 478.090000 ;
        RECT 251.000000 489.910000 256.000000 490.090000 ;
        RECT 251.000000 485.910000 256.000000 486.090000 ;
        RECT 4.000000 505.910000 14.000000 506.090000 ;
        RECT 4.000000 497.910000 14.000000 498.090000 ;
        RECT 4.000000 493.910000 14.000000 494.090000 ;
        RECT 4.000000 501.910000 14.000000 502.090000 ;
        RECT 4.000000 513.910000 14.000000 514.090000 ;
        RECT 4.000000 509.910000 14.000000 510.090000 ;
        RECT 51.000000 493.910000 56.000000 494.090000 ;
        RECT 51.000000 497.910000 56.000000 498.090000 ;
        RECT 51.000000 501.910000 56.000000 502.090000 ;
        RECT 51.000000 505.910000 56.000000 506.090000 ;
        RECT 51.000000 513.910000 56.000000 514.090000 ;
        RECT 51.000000 509.910000 56.000000 510.090000 ;
        RECT 101.000000 505.910000 106.000000 506.090000 ;
        RECT 101.000000 501.910000 106.000000 502.090000 ;
        RECT 101.000000 497.910000 106.000000 498.090000 ;
        RECT 101.000000 493.910000 106.000000 494.090000 ;
        RECT 101.000000 513.910000 106.000000 514.090000 ;
        RECT 101.000000 509.910000 106.000000 510.090000 ;
        RECT 151.000000 493.910000 156.000000 494.090000 ;
        RECT 151.000000 497.910000 156.000000 498.090000 ;
        RECT 151.000000 501.910000 156.000000 502.090000 ;
        RECT 151.000000 505.910000 156.000000 506.090000 ;
        RECT 151.000000 509.910000 156.000000 510.090000 ;
        RECT 151.000000 513.910000 156.000000 514.090000 ;
        RECT 201.000000 497.910000 206.000000 498.090000 ;
        RECT 201.000000 493.910000 206.000000 494.090000 ;
        RECT 201.000000 501.910000 206.000000 502.090000 ;
        RECT 201.000000 505.910000 206.000000 506.090000 ;
        RECT 201.000000 513.910000 206.000000 514.090000 ;
        RECT 201.000000 509.910000 206.000000 510.090000 ;
        RECT 251.000000 493.910000 256.000000 494.090000 ;
        RECT 251.000000 497.910000 256.000000 498.090000 ;
        RECT 251.000000 501.910000 256.000000 502.090000 ;
        RECT 251.000000 505.910000 256.000000 506.090000 ;
        RECT 251.000000 509.910000 256.000000 510.090000 ;
        RECT 251.000000 513.910000 256.000000 514.090000 ;
        RECT 301.000000 345.910000 306.000000 346.090000 ;
        RECT 301.000000 349.910000 306.000000 350.090000 ;
        RECT 301.000000 353.910000 306.000000 354.090000 ;
        RECT 301.000000 357.910000 306.000000 358.090000 ;
        RECT 301.000000 369.910000 306.000000 370.090000 ;
        RECT 301.000000 365.910000 306.000000 366.090000 ;
        RECT 301.000000 361.910000 306.000000 362.090000 ;
        RECT 301.000000 377.910000 306.000000 378.090000 ;
        RECT 301.000000 373.910000 306.000000 374.090000 ;
        RECT 351.000000 345.910000 356.000000 346.090000 ;
        RECT 351.000000 349.910000 356.000000 350.090000 ;
        RECT 351.000000 353.910000 356.000000 354.090000 ;
        RECT 351.000000 357.910000 356.000000 358.090000 ;
        RECT 351.000000 361.910000 356.000000 362.090000 ;
        RECT 351.000000 365.910000 356.000000 366.090000 ;
        RECT 351.000000 369.910000 356.000000 370.090000 ;
        RECT 351.000000 373.910000 356.000000 374.090000 ;
        RECT 351.000000 377.910000 356.000000 378.090000 ;
        RECT 301.000000 385.910000 306.000000 386.090000 ;
        RECT 301.000000 381.910000 306.000000 382.090000 ;
        RECT 301.000000 389.910000 306.000000 390.090000 ;
        RECT 301.000000 393.910000 306.000000 394.090000 ;
        RECT 301.000000 397.910000 306.000000 398.090000 ;
        RECT 301.000000 405.910000 306.000000 406.090000 ;
        RECT 301.000000 401.910000 306.000000 402.090000 ;
        RECT 301.000000 413.910000 306.000000 414.090000 ;
        RECT 301.000000 409.910000 306.000000 410.090000 ;
        RECT 351.000000 381.910000 356.000000 382.090000 ;
        RECT 351.000000 385.910000 356.000000 386.090000 ;
        RECT 351.000000 397.910000 356.000000 398.090000 ;
        RECT 351.000000 393.910000 356.000000 394.090000 ;
        RECT 351.000000 389.910000 356.000000 390.090000 ;
        RECT 351.000000 413.910000 356.000000 414.090000 ;
        RECT 351.000000 409.910000 356.000000 410.090000 ;
        RECT 351.000000 405.910000 356.000000 406.090000 ;
        RECT 351.000000 401.910000 356.000000 402.090000 ;
        RECT 401.000000 345.910000 406.000000 346.090000 ;
        RECT 401.000000 349.910000 406.000000 350.090000 ;
        RECT 401.000000 353.910000 406.000000 354.090000 ;
        RECT 401.000000 357.910000 406.000000 358.090000 ;
        RECT 401.000000 369.910000 406.000000 370.090000 ;
        RECT 401.000000 365.910000 406.000000 366.090000 ;
        RECT 401.000000 361.910000 406.000000 362.090000 ;
        RECT 401.000000 373.910000 406.000000 374.090000 ;
        RECT 401.000000 377.910000 406.000000 378.090000 ;
        RECT 401.000000 381.910000 406.000000 382.090000 ;
        RECT 401.000000 385.910000 406.000000 386.090000 ;
        RECT 401.000000 393.910000 406.000000 394.090000 ;
        RECT 401.000000 389.910000 406.000000 390.090000 ;
        RECT 401.000000 397.910000 406.000000 398.090000 ;
        RECT 401.000000 401.910000 406.000000 402.090000 ;
        RECT 401.000000 405.910000 406.000000 406.090000 ;
        RECT 401.000000 413.910000 406.000000 414.090000 ;
        RECT 401.000000 409.910000 406.000000 410.090000 ;
        RECT 301.000000 425.910000 306.000000 426.090000 ;
        RECT 301.000000 417.910000 306.000000 418.090000 ;
        RECT 301.000000 421.910000 306.000000 422.090000 ;
        RECT 301.000000 429.910000 306.000000 430.090000 ;
        RECT 301.000000 433.910000 306.000000 434.090000 ;
        RECT 301.000000 441.910000 306.000000 442.090000 ;
        RECT 301.000000 437.910000 306.000000 438.090000 ;
        RECT 301.000000 453.910000 306.000000 454.090000 ;
        RECT 301.000000 449.910000 306.000000 450.090000 ;
        RECT 301.000000 445.910000 306.000000 446.090000 ;
        RECT 351.000000 425.910000 356.000000 426.090000 ;
        RECT 351.000000 421.910000 356.000000 422.090000 ;
        RECT 351.000000 417.910000 356.000000 418.090000 ;
        RECT 351.000000 433.910000 356.000000 434.090000 ;
        RECT 351.000000 429.910000 356.000000 430.090000 ;
        RECT 351.000000 437.910000 356.000000 438.090000 ;
        RECT 351.000000 441.910000 356.000000 442.090000 ;
        RECT 351.000000 445.910000 356.000000 446.090000 ;
        RECT 351.000000 449.910000 356.000000 450.090000 ;
        RECT 351.000000 453.910000 356.000000 454.090000 ;
        RECT 301.000000 461.910000 306.000000 462.090000 ;
        RECT 301.000000 457.910000 306.000000 458.090000 ;
        RECT 301.000000 465.910000 306.000000 466.090000 ;
        RECT 301.000000 469.910000 306.000000 470.090000 ;
        RECT 301.000000 481.910000 306.000000 482.090000 ;
        RECT 301.000000 477.910000 306.000000 478.090000 ;
        RECT 301.000000 473.910000 306.000000 474.090000 ;
        RECT 301.000000 489.910000 306.000000 490.090000 ;
        RECT 301.000000 485.910000 306.000000 486.090000 ;
        RECT 351.000000 457.910000 356.000000 458.090000 ;
        RECT 351.000000 461.910000 356.000000 462.090000 ;
        RECT 351.000000 469.910000 356.000000 470.090000 ;
        RECT 351.000000 465.910000 356.000000 466.090000 ;
        RECT 351.000000 481.910000 356.000000 482.090000 ;
        RECT 351.000000 473.910000 356.000000 474.090000 ;
        RECT 351.000000 477.910000 356.000000 478.090000 ;
        RECT 351.000000 485.910000 356.000000 486.090000 ;
        RECT 351.000000 489.910000 356.000000 490.090000 ;
        RECT 401.000000 417.910000 406.000000 418.090000 ;
        RECT 401.000000 421.910000 406.000000 422.090000 ;
        RECT 401.000000 425.910000 406.000000 426.090000 ;
        RECT 401.000000 429.910000 406.000000 430.090000 ;
        RECT 401.000000 433.910000 406.000000 434.090000 ;
        RECT 401.000000 437.910000 406.000000 438.090000 ;
        RECT 401.000000 441.910000 406.000000 442.090000 ;
        RECT 401.000000 445.910000 406.000000 446.090000 ;
        RECT 401.000000 453.910000 406.000000 454.090000 ;
        RECT 401.000000 449.910000 406.000000 450.090000 ;
        RECT 401.000000 457.910000 406.000000 458.090000 ;
        RECT 401.000000 461.910000 406.000000 462.090000 ;
        RECT 401.000000 465.910000 406.000000 466.090000 ;
        RECT 401.000000 469.910000 406.000000 470.090000 ;
        RECT 401.000000 481.910000 406.000000 482.090000 ;
        RECT 401.000000 473.910000 406.000000 474.090000 ;
        RECT 401.000000 477.910000 406.000000 478.090000 ;
        RECT 401.000000 485.910000 406.000000 486.090000 ;
        RECT 401.000000 489.910000 406.000000 490.090000 ;
        RECT 451.000000 345.910000 456.000000 346.090000 ;
        RECT 451.000000 366.105000 456.000000 367.105000 ;
        RECT 451.000000 369.910000 456.000000 370.090000 ;
        RECT 451.000000 373.910000 456.000000 374.090000 ;
        RECT 451.000000 377.910000 456.000000 378.090000 ;
        RECT 501.000000 345.910000 506.000000 346.090000 ;
        RECT 501.000000 349.910000 506.000000 350.090000 ;
        RECT 501.000000 353.910000 506.000000 354.090000 ;
        RECT 501.000000 357.910000 506.000000 358.090000 ;
        RECT 501.000000 361.910000 506.000000 362.090000 ;
        RECT 501.000000 365.910000 506.000000 366.090000 ;
        RECT 501.000000 369.910000 506.000000 370.090000 ;
        RECT 501.000000 377.910000 506.000000 378.090000 ;
        RECT 501.000000 373.910000 506.000000 374.090000 ;
        RECT 451.000000 381.910000 456.000000 382.090000 ;
        RECT 451.000000 385.910000 456.000000 386.090000 ;
        RECT 451.000000 397.910000 456.000000 398.090000 ;
        RECT 451.000000 393.910000 456.000000 394.090000 ;
        RECT 451.000000 389.910000 456.000000 390.090000 ;
        RECT 451.000000 416.105000 456.000000 417.105000 ;
        RECT 501.000000 381.910000 506.000000 382.090000 ;
        RECT 501.000000 385.910000 506.000000 386.090000 ;
        RECT 501.000000 393.910000 506.000000 394.090000 ;
        RECT 501.000000 389.910000 506.000000 390.090000 ;
        RECT 501.000000 397.910000 506.000000 398.090000 ;
        RECT 501.000000 401.910000 506.000000 402.090000 ;
        RECT 501.000000 405.910000 506.000000 406.090000 ;
        RECT 501.000000 409.910000 506.000000 410.090000 ;
        RECT 501.000000 413.910000 506.000000 414.090000 ;
        RECT 551.000000 357.910000 556.000000 358.090000 ;
        RECT 551.000000 353.910000 556.000000 354.090000 ;
        RECT 551.000000 349.910000 556.000000 350.090000 ;
        RECT 551.000000 345.910000 556.000000 346.090000 ;
        RECT 551.000000 361.910000 556.000000 362.090000 ;
        RECT 551.000000 365.910000 556.000000 366.090000 ;
        RECT 551.000000 369.910000 556.000000 370.090000 ;
        RECT 551.000000 373.910000 556.000000 374.090000 ;
        RECT 551.000000 377.910000 556.000000 378.090000 ;
        RECT 551.000000 385.910000 556.000000 386.090000 ;
        RECT 551.000000 381.910000 556.000000 382.090000 ;
        RECT 551.000000 397.910000 556.000000 398.090000 ;
        RECT 551.000000 393.910000 556.000000 394.090000 ;
        RECT 551.000000 389.910000 556.000000 390.090000 ;
        RECT 551.000000 401.910000 556.000000 402.090000 ;
        RECT 551.000000 405.910000 556.000000 406.090000 ;
        RECT 551.000000 409.910000 556.000000 410.090000 ;
        RECT 551.000000 413.910000 556.000000 414.090000 ;
        RECT 451.000000 425.910000 456.000000 426.090000 ;
        RECT 451.000000 421.910000 456.000000 422.090000 ;
        RECT 451.000000 429.910000 456.000000 430.090000 ;
        RECT 451.000000 433.910000 456.000000 434.090000 ;
        RECT 451.000000 441.910000 456.000000 442.090000 ;
        RECT 451.000000 437.910000 456.000000 438.090000 ;
        RECT 451.000000 453.910000 456.000000 454.090000 ;
        RECT 451.000000 449.910000 456.000000 450.090000 ;
        RECT 451.000000 445.910000 456.000000 446.090000 ;
        RECT 501.000000 425.910000 506.000000 426.090000 ;
        RECT 501.000000 421.910000 506.000000 422.090000 ;
        RECT 501.000000 417.910000 506.000000 418.090000 ;
        RECT 501.000000 429.910000 506.000000 430.090000 ;
        RECT 501.000000 433.910000 506.000000 434.090000 ;
        RECT 501.000000 437.910000 506.000000 438.090000 ;
        RECT 501.000000 441.910000 506.000000 442.090000 ;
        RECT 501.000000 445.910000 506.000000 446.090000 ;
        RECT 501.000000 449.910000 506.000000 450.090000 ;
        RECT 501.000000 453.910000 506.000000 454.090000 ;
        RECT 451.000000 461.910000 456.000000 462.090000 ;
        RECT 451.000000 457.910000 456.000000 458.090000 ;
        RECT 451.000000 465.910000 456.000000 466.090000 ;
        RECT 451.000000 469.910000 456.000000 470.090000 ;
        RECT 451.000000 481.910000 456.000000 482.090000 ;
        RECT 451.000000 477.910000 456.000000 478.090000 ;
        RECT 451.000000 473.910000 456.000000 474.090000 ;
        RECT 451.000000 489.910000 456.000000 490.090000 ;
        RECT 451.000000 485.910000 456.000000 486.090000 ;
        RECT 501.000000 461.910000 506.000000 462.090000 ;
        RECT 501.000000 457.910000 506.000000 458.090000 ;
        RECT 501.000000 469.910000 506.000000 470.090000 ;
        RECT 501.000000 465.910000 506.000000 466.090000 ;
        RECT 501.000000 481.910000 506.000000 482.090000 ;
        RECT 501.000000 477.910000 506.000000 478.090000 ;
        RECT 501.000000 473.910000 506.000000 474.090000 ;
        RECT 501.000000 489.910000 506.000000 490.090000 ;
        RECT 501.000000 485.910000 506.000000 486.090000 ;
        RECT 551.000000 417.910000 556.000000 418.090000 ;
        RECT 551.000000 425.910000 556.000000 426.090000 ;
        RECT 551.000000 421.910000 556.000000 422.090000 ;
        RECT 551.000000 433.910000 556.000000 434.090000 ;
        RECT 551.000000 429.910000 556.000000 430.090000 ;
        RECT 551.000000 437.910000 556.000000 438.090000 ;
        RECT 551.000000 441.910000 556.000000 442.090000 ;
        RECT 551.000000 445.910000 556.000000 446.090000 ;
        RECT 551.000000 449.910000 556.000000 450.090000 ;
        RECT 551.000000 453.910000 556.000000 454.090000 ;
        RECT 551.000000 461.910000 556.000000 462.090000 ;
        RECT 551.000000 457.910000 556.000000 458.090000 ;
        RECT 551.000000 469.910000 556.000000 470.090000 ;
        RECT 551.000000 465.910000 556.000000 466.090000 ;
        RECT 551.000000 481.910000 556.000000 482.090000 ;
        RECT 551.000000 473.910000 556.000000 474.090000 ;
        RECT 551.000000 477.910000 556.000000 478.090000 ;
        RECT 551.000000 485.910000 556.000000 486.090000 ;
        RECT 551.000000 489.910000 556.000000 490.090000 ;
        RECT 301.000000 497.910000 306.000000 498.090000 ;
        RECT 301.000000 493.910000 306.000000 494.090000 ;
        RECT 301.000000 501.910000 306.000000 502.090000 ;
        RECT 301.000000 505.910000 306.000000 506.090000 ;
        RECT 301.000000 517.910000 306.000000 518.090000 ;
        RECT 301.000000 513.910000 306.000000 514.090000 ;
        RECT 301.000000 509.910000 306.000000 510.090000 ;
        RECT 351.000000 493.910000 356.000000 494.090000 ;
        RECT 351.000000 497.910000 356.000000 498.090000 ;
        RECT 351.000000 505.910000 356.000000 506.090000 ;
        RECT 351.000000 501.910000 356.000000 502.090000 ;
        RECT 351.000000 509.910000 356.000000 510.090000 ;
        RECT 351.000000 513.910000 356.000000 514.090000 ;
        RECT 351.000000 517.910000 356.000000 518.090000 ;
        RECT 351.000000 521.910000 356.000000 522.090000 ;
        RECT 351.000000 525.910000 356.000000 526.090000 ;
        RECT 351.000000 537.910000 356.000000 538.090000 ;
        RECT 351.000000 533.910000 356.000000 534.090000 ;
        RECT 351.000000 529.910000 356.000000 530.090000 ;
        RECT 351.000000 541.910000 356.000000 542.090000 ;
        RECT 351.000000 545.910000 356.000000 546.090000 ;
        RECT 351.000000 549.910000 356.000000 550.090000 ;
        RECT 351.000000 553.910000 356.000000 554.090000 ;
        RECT 351.000000 557.910000 356.000000 558.090000 ;
        RECT 351.000000 561.910000 356.000000 562.090000 ;
        RECT 375.000000 493.910000 385.000000 494.090000 ;
        RECT 375.000000 497.910000 385.000000 498.090000 ;
        RECT 375.000000 501.910000 385.000000 502.090000 ;
        RECT 375.000000 505.910000 385.000000 506.090000 ;
        RECT 401.000000 493.910000 406.000000 494.090000 ;
        RECT 401.000000 497.910000 406.000000 498.090000 ;
        RECT 401.000000 501.910000 406.000000 502.090000 ;
        RECT 375.000000 517.910000 385.000000 518.090000 ;
        RECT 375.000000 513.910000 385.000000 514.090000 ;
        RECT 375.000000 509.910000 385.000000 510.090000 ;
        RECT 375.000000 525.910000 385.000000 526.090000 ;
        RECT 375.000000 521.910000 385.000000 522.090000 ;
        RECT 375.000000 533.910000 385.000000 534.090000 ;
        RECT 375.000000 529.910000 385.000000 530.090000 ;
        RECT 375.000000 545.910000 385.000000 546.090000 ;
        RECT 375.000000 541.910000 385.000000 542.090000 ;
        RECT 375.000000 537.910000 385.000000 538.090000 ;
        RECT 375.000000 553.910000 385.000000 554.090000 ;
        RECT 375.000000 549.910000 385.000000 550.090000 ;
        RECT 375.000000 561.910000 385.000000 562.090000 ;
        RECT 375.000000 557.910000 385.000000 558.090000 ;
        RECT 351.000000 581.910000 356.000000 582.090000 ;
        RECT 351.000000 577.910000 356.000000 578.090000 ;
        RECT 351.000000 573.910000 356.000000 574.090000 ;
        RECT 351.000000 569.910000 356.000000 570.090000 ;
        RECT 351.000000 565.910000 356.000000 566.090000 ;
        RECT 351.000000 601.910000 356.000000 602.090000 ;
        RECT 351.000000 597.910000 356.000000 598.090000 ;
        RECT 351.000000 593.910000 356.000000 594.090000 ;
        RECT 351.000000 589.910000 356.000000 590.090000 ;
        RECT 351.000000 585.910000 356.000000 586.090000 ;
        RECT 351.000000 609.910000 356.000000 610.090000 ;
        RECT 351.000000 605.910000 356.000000 606.090000 ;
        RECT 351.000000 613.910000 356.000000 614.090000 ;
        RECT 351.000000 617.910000 356.000000 618.090000 ;
        RECT 351.000000 637.910000 356.000000 638.090000 ;
        RECT 351.000000 633.910000 356.000000 634.090000 ;
        RECT 351.000000 629.910000 356.000000 630.090000 ;
        RECT 351.000000 625.910000 356.000000 626.090000 ;
        RECT 351.000000 621.910000 356.000000 622.090000 ;
        RECT 375.000000 565.910000 385.000000 566.090000 ;
        RECT 375.000000 569.910000 385.000000 570.090000 ;
        RECT 375.000000 573.910000 385.000000 574.090000 ;
        RECT 375.000000 577.910000 385.000000 578.090000 ;
        RECT 375.000000 581.910000 385.000000 582.090000 ;
        RECT 375.000000 589.910000 385.000000 590.090000 ;
        RECT 375.000000 585.910000 385.000000 586.090000 ;
        RECT 375.000000 601.910000 385.000000 602.090000 ;
        RECT 375.000000 597.910000 385.000000 598.090000 ;
        RECT 375.000000 593.910000 385.000000 594.090000 ;
        RECT 375.000000 609.910000 385.000000 610.090000 ;
        RECT 375.000000 605.910000 385.000000 606.090000 ;
        RECT 375.000000 617.910000 385.000000 618.090000 ;
        RECT 375.000000 613.910000 385.000000 614.090000 ;
        RECT 375.000000 629.910000 385.000000 630.090000 ;
        RECT 375.000000 625.910000 385.000000 626.090000 ;
        RECT 375.000000 621.910000 385.000000 622.090000 ;
        RECT 375.000000 637.910000 385.000000 638.090000 ;
        RECT 375.000000 633.910000 385.000000 634.090000 ;
        RECT 451.000000 493.910000 456.000000 494.090000 ;
        RECT 451.000000 497.910000 456.000000 498.090000 ;
        RECT 451.000000 501.910000 456.000000 502.090000 ;
        RECT 501.000000 493.910000 506.000000 494.090000 ;
        RECT 501.000000 497.910000 506.000000 498.090000 ;
        RECT 501.000000 501.910000 506.000000 502.090000 ;
        RECT 551.000000 493.910000 556.000000 494.090000 ;
        RECT 551.000000 497.910000 556.000000 498.090000 ;
        RECT 551.000000 501.910000 556.000000 502.090000 ;
        RECT 351.000000 657.910000 356.000000 658.090000 ;
        RECT 351.000000 641.910000 356.000000 642.090000 ;
        RECT 351.000000 645.910000 356.000000 646.090000 ;
        RECT 351.000000 649.910000 356.000000 650.090000 ;
        RECT 351.000000 653.910000 356.000000 654.090000 ;
        RECT 351.000000 673.910000 356.000000 674.090000 ;
        RECT 351.000000 669.910000 356.000000 670.090000 ;
        RECT 351.000000 665.910000 356.000000 666.090000 ;
        RECT 351.000000 661.910000 356.000000 662.090000 ;
        RECT 301.000000 677.910000 306.000000 678.090000 ;
        RECT 301.000000 681.910000 306.000000 682.090000 ;
        RECT 351.000000 681.910000 356.000000 682.090000 ;
        RECT 351.000000 677.910000 356.000000 678.090000 ;
        RECT 375.000000 657.910000 385.000000 658.090000 ;
        RECT 401.000000 657.910000 406.000000 658.090000 ;
        RECT 375.000000 641.910000 385.000000 642.090000 ;
        RECT 375.000000 645.910000 385.000000 646.090000 ;
        RECT 375.000000 649.910000 385.000000 650.090000 ;
        RECT 375.000000 653.910000 385.000000 654.090000 ;
        RECT 375.000000 665.910000 385.000000 666.090000 ;
        RECT 375.000000 661.910000 385.000000 662.090000 ;
        RECT 375.000000 669.910000 385.000000 670.090000 ;
        RECT 375.000000 673.910000 385.000000 674.090000 ;
        RECT 401.000000 673.910000 406.000000 674.090000 ;
        RECT 401.000000 661.910000 406.000000 662.090000 ;
        RECT 401.000000 665.910000 406.000000 666.090000 ;
        RECT 401.000000 669.910000 406.000000 670.090000 ;
        RECT 375.000000 681.910000 385.000000 682.090000 ;
        RECT 375.000000 677.910000 385.000000 678.090000 ;
        RECT 401.000000 677.910000 406.000000 678.090000 ;
        RECT 401.000000 681.910000 406.000000 682.090000 ;
        RECT 451.000000 657.910000 456.000000 658.090000 ;
        RECT 451.000000 673.910000 456.000000 674.090000 ;
        RECT 451.000000 669.910000 456.000000 670.090000 ;
        RECT 451.000000 665.910000 456.000000 666.090000 ;
        RECT 451.000000 661.910000 456.000000 662.090000 ;
        RECT 501.000000 657.910000 506.000000 658.090000 ;
        RECT 501.000000 665.910000 506.000000 666.090000 ;
        RECT 501.000000 661.910000 506.000000 662.090000 ;
        RECT 501.000000 673.910000 506.000000 674.090000 ;
        RECT 501.000000 669.910000 506.000000 670.090000 ;
        RECT 451.000000 677.910000 456.000000 678.090000 ;
        RECT 451.000000 681.910000 456.000000 682.090000 ;
        RECT 501.000000 677.910000 506.000000 678.090000 ;
        RECT 501.000000 681.910000 506.000000 682.090000 ;
        RECT 551.000000 657.910000 556.000000 658.090000 ;
        RECT 551.000000 661.910000 556.000000 662.090000 ;
        RECT 551.000000 665.910000 556.000000 666.090000 ;
        RECT 551.000000 669.910000 556.000000 670.090000 ;
        RECT 551.000000 673.910000 556.000000 674.090000 ;
        RECT 551.000000 681.910000 556.000000 682.090000 ;
        RECT 551.000000 677.910000 556.000000 678.090000 ;
        RECT 601.000000 345.910000 606.000000 346.090000 ;
        RECT 601.000000 349.910000 606.000000 350.090000 ;
        RECT 601.000000 353.910000 606.000000 354.090000 ;
        RECT 601.000000 357.910000 606.000000 358.090000 ;
        RECT 601.000000 369.910000 606.000000 370.090000 ;
        RECT 601.000000 365.910000 606.000000 366.090000 ;
        RECT 601.000000 361.910000 606.000000 362.090000 ;
        RECT 601.000000 377.910000 606.000000 378.090000 ;
        RECT 601.000000 373.910000 606.000000 374.090000 ;
        RECT 651.000000 349.910000 656.000000 350.090000 ;
        RECT 651.000000 345.910000 656.000000 346.090000 ;
        RECT 651.000000 357.910000 656.000000 358.090000 ;
        RECT 651.000000 353.910000 656.000000 354.090000 ;
        RECT 651.000000 361.910000 656.000000 362.090000 ;
        RECT 651.000000 365.910000 656.000000 366.090000 ;
        RECT 651.000000 369.910000 656.000000 370.090000 ;
        RECT 651.000000 373.910000 656.000000 374.090000 ;
        RECT 651.000000 377.910000 656.000000 378.090000 ;
        RECT 601.000000 385.910000 606.000000 386.090000 ;
        RECT 601.000000 381.910000 606.000000 382.090000 ;
        RECT 601.000000 389.910000 606.000000 390.090000 ;
        RECT 601.000000 393.910000 606.000000 394.090000 ;
        RECT 601.000000 397.910000 606.000000 398.090000 ;
        RECT 601.000000 405.910000 606.000000 406.090000 ;
        RECT 601.000000 401.910000 606.000000 402.090000 ;
        RECT 601.000000 413.910000 606.000000 414.090000 ;
        RECT 601.000000 409.910000 606.000000 410.090000 ;
        RECT 651.000000 381.910000 656.000000 382.090000 ;
        RECT 651.000000 385.910000 656.000000 386.090000 ;
        RECT 651.000000 393.910000 656.000000 394.090000 ;
        RECT 651.000000 389.910000 656.000000 390.090000 ;
        RECT 651.000000 397.910000 656.000000 398.090000 ;
        RECT 651.000000 405.910000 656.000000 406.090000 ;
        RECT 651.000000 401.910000 656.000000 402.090000 ;
        RECT 651.000000 409.910000 656.000000 410.090000 ;
        RECT 651.000000 413.910000 656.000000 414.090000 ;
        RECT 701.000000 357.910000 706.000000 358.090000 ;
        RECT 701.000000 353.910000 706.000000 354.090000 ;
        RECT 701.000000 349.910000 706.000000 350.090000 ;
        RECT 701.000000 345.910000 706.000000 346.090000 ;
        RECT 701.000000 361.910000 706.000000 362.090000 ;
        RECT 701.000000 365.910000 706.000000 366.090000 ;
        RECT 701.000000 369.910000 706.000000 370.090000 ;
        RECT 701.000000 373.910000 706.000000 374.090000 ;
        RECT 701.000000 377.910000 706.000000 378.090000 ;
        RECT 701.000000 385.910000 706.000000 386.090000 ;
        RECT 701.000000 381.910000 706.000000 382.090000 ;
        RECT 701.000000 397.910000 706.000000 398.090000 ;
        RECT 701.000000 393.910000 706.000000 394.090000 ;
        RECT 701.000000 389.910000 706.000000 390.090000 ;
        RECT 701.000000 413.910000 706.000000 414.090000 ;
        RECT 701.000000 409.910000 706.000000 410.090000 ;
        RECT 701.000000 405.910000 706.000000 406.090000 ;
        RECT 701.000000 401.910000 706.000000 402.090000 ;
        RECT 601.000000 417.910000 606.000000 418.090000 ;
        RECT 601.000000 421.910000 606.000000 422.090000 ;
        RECT 601.000000 425.910000 606.000000 426.090000 ;
        RECT 601.000000 429.910000 606.000000 430.090000 ;
        RECT 601.000000 433.910000 606.000000 434.090000 ;
        RECT 601.000000 441.910000 606.000000 442.090000 ;
        RECT 601.000000 437.910000 606.000000 438.090000 ;
        RECT 601.000000 453.910000 606.000000 454.090000 ;
        RECT 601.000000 449.910000 606.000000 450.090000 ;
        RECT 601.000000 445.910000 606.000000 446.090000 ;
        RECT 651.000000 421.910000 656.000000 422.090000 ;
        RECT 651.000000 417.910000 656.000000 418.090000 ;
        RECT 651.000000 425.910000 656.000000 426.090000 ;
        RECT 651.000000 429.910000 656.000000 430.090000 ;
        RECT 651.000000 433.910000 656.000000 434.090000 ;
        RECT 651.000000 437.910000 656.000000 438.090000 ;
        RECT 651.000000 441.910000 656.000000 442.090000 ;
        RECT 651.000000 445.910000 656.000000 446.090000 ;
        RECT 651.000000 449.910000 656.000000 450.090000 ;
        RECT 651.000000 453.910000 656.000000 454.090000 ;
        RECT 601.000000 461.910000 606.000000 462.090000 ;
        RECT 601.000000 457.910000 606.000000 458.090000 ;
        RECT 601.000000 465.910000 606.000000 466.090000 ;
        RECT 601.000000 469.910000 606.000000 470.090000 ;
        RECT 601.000000 481.910000 606.000000 482.090000 ;
        RECT 601.000000 477.910000 606.000000 478.090000 ;
        RECT 601.000000 473.910000 606.000000 474.090000 ;
        RECT 601.000000 489.910000 606.000000 490.090000 ;
        RECT 601.000000 485.910000 606.000000 486.090000 ;
        RECT 651.000000 461.910000 656.000000 462.090000 ;
        RECT 651.000000 457.910000 656.000000 458.090000 ;
        RECT 651.000000 469.910000 656.000000 470.090000 ;
        RECT 651.000000 465.910000 656.000000 466.090000 ;
        RECT 651.000000 481.910000 656.000000 482.090000 ;
        RECT 651.000000 477.910000 656.000000 478.090000 ;
        RECT 651.000000 473.910000 656.000000 474.090000 ;
        RECT 651.000000 489.910000 656.000000 490.090000 ;
        RECT 651.000000 485.910000 656.000000 486.090000 ;
        RECT 701.000000 417.910000 706.000000 418.090000 ;
        RECT 701.000000 421.910000 706.000000 422.090000 ;
        RECT 701.000000 425.910000 706.000000 426.090000 ;
        RECT 701.000000 433.910000 706.000000 434.090000 ;
        RECT 701.000000 429.910000 706.000000 430.090000 ;
        RECT 701.000000 437.910000 706.000000 438.090000 ;
        RECT 701.000000 441.910000 706.000000 442.090000 ;
        RECT 701.000000 445.910000 706.000000 446.090000 ;
        RECT 701.000000 449.910000 706.000000 450.090000 ;
        RECT 701.000000 453.910000 706.000000 454.090000 ;
        RECT 725.000000 433.910000 735.000000 434.090000 ;
        RECT 725.000000 437.910000 735.000000 438.090000 ;
        RECT 725.000000 441.910000 735.000000 442.090000 ;
        RECT 725.000000 453.910000 735.000000 454.090000 ;
        RECT 725.000000 449.910000 735.000000 450.090000 ;
        RECT 725.000000 445.910000 735.000000 446.090000 ;
        RECT 701.000000 457.910000 706.000000 458.090000 ;
        RECT 701.000000 461.910000 706.000000 462.090000 ;
        RECT 701.000000 465.910000 706.000000 466.090000 ;
        RECT 701.000000 469.910000 706.000000 470.090000 ;
        RECT 701.000000 481.910000 706.000000 482.090000 ;
        RECT 701.000000 473.910000 706.000000 474.090000 ;
        RECT 701.000000 477.910000 706.000000 478.090000 ;
        RECT 701.000000 485.910000 706.000000 486.090000 ;
        RECT 701.000000 489.910000 706.000000 490.090000 ;
        RECT 725.000000 469.910000 735.000000 470.090000 ;
        RECT 725.000000 457.910000 735.000000 458.090000 ;
        RECT 725.000000 461.910000 735.000000 462.090000 ;
        RECT 725.000000 465.910000 735.000000 466.090000 ;
        RECT 725.000000 481.910000 735.000000 482.090000 ;
        RECT 725.000000 477.910000 735.000000 478.090000 ;
        RECT 725.000000 473.910000 735.000000 474.090000 ;
        RECT 725.000000 489.910000 735.000000 490.090000 ;
        RECT 725.000000 485.910000 735.000000 486.090000 ;
        RECT 751.000000 349.910000 756.000000 350.090000 ;
        RECT 751.000000 345.910000 756.000000 346.090000 ;
        RECT 751.000000 353.910000 756.000000 354.090000 ;
        RECT 751.000000 357.910000 756.000000 358.090000 ;
        RECT 751.000000 369.910000 756.000000 370.090000 ;
        RECT 751.000000 365.910000 756.000000 366.090000 ;
        RECT 751.000000 361.910000 756.000000 362.090000 ;
        RECT 751.000000 373.910000 756.000000 374.090000 ;
        RECT 751.000000 377.910000 756.000000 378.090000 ;
        RECT 801.000000 349.910000 806.000000 350.090000 ;
        RECT 801.000000 345.910000 806.000000 346.090000 ;
        RECT 801.000000 353.910000 806.000000 354.090000 ;
        RECT 801.000000 357.910000 806.000000 358.090000 ;
        RECT 801.000000 361.910000 806.000000 362.090000 ;
        RECT 801.000000 365.910000 806.000000 366.090000 ;
        RECT 801.000000 369.910000 806.000000 370.090000 ;
        RECT 801.000000 373.910000 806.000000 374.090000 ;
        RECT 801.000000 377.910000 806.000000 378.090000 ;
        RECT 751.000000 397.910000 756.000000 398.090000 ;
        RECT 751.000000 393.910000 756.000000 394.090000 ;
        RECT 751.000000 389.910000 756.000000 390.090000 ;
        RECT 751.000000 381.910000 756.000000 382.090000 ;
        RECT 751.000000 385.910000 756.000000 386.090000 ;
        RECT 751.000000 401.910000 756.000000 402.090000 ;
        RECT 751.000000 405.910000 756.000000 406.090000 ;
        RECT 751.000000 409.910000 756.000000 410.090000 ;
        RECT 751.000000 413.910000 756.000000 414.090000 ;
        RECT 801.000000 385.910000 806.000000 386.090000 ;
        RECT 801.000000 381.910000 806.000000 382.090000 ;
        RECT 801.000000 397.910000 806.000000 398.090000 ;
        RECT 801.000000 393.910000 806.000000 394.090000 ;
        RECT 801.000000 389.910000 806.000000 390.090000 ;
        RECT 801.000000 405.910000 806.000000 406.090000 ;
        RECT 801.000000 401.910000 806.000000 402.090000 ;
        RECT 801.000000 409.910000 806.000000 410.090000 ;
        RECT 801.000000 413.910000 806.000000 414.090000 ;
        RECT 851.000000 357.910000 856.000000 358.090000 ;
        RECT 851.000000 353.910000 856.000000 354.090000 ;
        RECT 851.000000 349.910000 856.000000 350.090000 ;
        RECT 851.000000 345.910000 856.000000 346.090000 ;
        RECT 851.000000 361.910000 856.000000 362.090000 ;
        RECT 851.000000 365.910000 856.000000 366.090000 ;
        RECT 851.000000 369.910000 856.000000 370.090000 ;
        RECT 851.000000 373.910000 856.000000 374.090000 ;
        RECT 851.000000 377.910000 856.000000 378.090000 ;
        RECT 851.000000 385.910000 856.000000 386.090000 ;
        RECT 851.000000 381.910000 856.000000 382.090000 ;
        RECT 851.000000 397.910000 856.000000 398.090000 ;
        RECT 851.000000 393.910000 856.000000 394.090000 ;
        RECT 851.000000 389.910000 856.000000 390.090000 ;
        RECT 851.000000 413.910000 856.000000 414.090000 ;
        RECT 851.000000 409.910000 856.000000 410.090000 ;
        RECT 851.000000 405.910000 856.000000 406.090000 ;
        RECT 851.000000 401.910000 856.000000 402.090000 ;
        RECT 751.000000 421.910000 756.000000 422.090000 ;
        RECT 751.000000 417.910000 756.000000 418.090000 ;
        RECT 751.000000 425.910000 756.000000 426.090000 ;
        RECT 751.000000 433.910000 756.000000 434.090000 ;
        RECT 751.000000 429.910000 756.000000 430.090000 ;
        RECT 751.000000 437.910000 756.000000 438.090000 ;
        RECT 751.000000 441.910000 756.000000 442.090000 ;
        RECT 801.000000 425.910000 806.000000 426.090000 ;
        RECT 801.000000 421.910000 806.000000 422.090000 ;
        RECT 801.000000 417.910000 806.000000 418.090000 ;
        RECT 801.000000 429.910000 806.000000 430.090000 ;
        RECT 801.000000 433.910000 806.000000 434.090000 ;
        RECT 801.000000 437.910000 806.000000 438.090000 ;
        RECT 801.000000 441.910000 806.000000 442.090000 ;
        RECT 851.000000 417.910000 856.000000 418.090000 ;
        RECT 851.000000 421.910000 856.000000 422.090000 ;
        RECT 851.000000 425.910000 856.000000 426.090000 ;
        RECT 851.000000 429.910000 856.000000 430.090000 ;
        RECT 851.000000 433.910000 856.000000 434.090000 ;
        RECT 851.000000 441.910000 856.000000 442.090000 ;
        RECT 851.000000 437.910000 856.000000 438.090000 ;
        RECT 601.000000 493.910000 606.000000 494.090000 ;
        RECT 601.000000 497.910000 606.000000 498.090000 ;
        RECT 601.000000 501.910000 606.000000 502.090000 ;
        RECT 651.000000 493.910000 656.000000 494.090000 ;
        RECT 651.000000 497.910000 656.000000 498.090000 ;
        RECT 651.000000 501.910000 656.000000 502.090000 ;
        RECT 701.000000 501.910000 706.000000 502.090000 ;
        RECT 701.000000 493.910000 706.000000 494.090000 ;
        RECT 701.000000 497.910000 706.000000 498.090000 ;
        RECT 725.000000 501.910000 735.000000 502.090000 ;
        RECT 725.000000 497.910000 735.000000 498.090000 ;
        RECT 725.000000 493.910000 735.000000 494.090000 ;
        RECT 901.000000 357.910000 906.000000 358.090000 ;
        RECT 901.000000 353.910000 906.000000 354.090000 ;
        RECT 901.000000 349.910000 906.000000 350.090000 ;
        RECT 901.000000 345.910000 906.000000 346.090000 ;
        RECT 901.000000 369.910000 906.000000 370.090000 ;
        RECT 901.000000 365.910000 906.000000 366.090000 ;
        RECT 901.000000 361.910000 906.000000 362.090000 ;
        RECT 901.000000 373.910000 906.000000 374.090000 ;
        RECT 901.000000 377.910000 906.000000 378.090000 ;
        RECT 951.000000 345.910000 956.000000 346.090000 ;
        RECT 951.000000 349.910000 956.000000 350.090000 ;
        RECT 951.000000 353.910000 956.000000 354.090000 ;
        RECT 951.000000 357.910000 956.000000 358.090000 ;
        RECT 951.000000 369.910000 956.000000 370.090000 ;
        RECT 951.000000 365.910000 956.000000 366.090000 ;
        RECT 951.000000 361.910000 956.000000 362.090000 ;
        RECT 951.000000 377.910000 956.000000 378.090000 ;
        RECT 951.000000 373.910000 956.000000 374.090000 ;
        RECT 901.000000 397.910000 906.000000 398.090000 ;
        RECT 901.000000 393.910000 906.000000 394.090000 ;
        RECT 901.000000 389.910000 906.000000 390.090000 ;
        RECT 901.000000 381.910000 906.000000 382.090000 ;
        RECT 901.000000 385.910000 906.000000 386.090000 ;
        RECT 901.000000 401.910000 906.000000 402.090000 ;
        RECT 901.000000 405.910000 906.000000 406.090000 ;
        RECT 901.000000 413.910000 906.000000 414.090000 ;
        RECT 901.000000 409.910000 906.000000 410.090000 ;
        RECT 951.000000 397.910000 956.000000 398.090000 ;
        RECT 951.000000 393.910000 956.000000 394.090000 ;
        RECT 951.000000 389.910000 956.000000 390.090000 ;
        RECT 951.000000 381.910000 956.000000 382.090000 ;
        RECT 951.000000 385.910000 956.000000 386.090000 ;
        RECT 951.000000 405.910000 956.000000 406.090000 ;
        RECT 951.000000 401.910000 956.000000 402.090000 ;
        RECT 951.000000 413.910000 956.000000 414.090000 ;
        RECT 951.000000 409.910000 956.000000 410.090000 ;
        RECT 1001.000000 349.910000 1006.000000 350.090000 ;
        RECT 1001.000000 345.910000 1006.000000 346.090000 ;
        RECT 1001.000000 353.910000 1006.000000 354.090000 ;
        RECT 1001.000000 357.910000 1006.000000 358.090000 ;
        RECT 1001.000000 361.910000 1006.000000 362.090000 ;
        RECT 1001.000000 365.910000 1006.000000 366.090000 ;
        RECT 1001.000000 369.910000 1006.000000 370.090000 ;
        RECT 1001.000000 373.910000 1006.000000 374.090000 ;
        RECT 1001.000000 377.910000 1006.000000 378.090000 ;
        RECT 1001.000000 385.910000 1006.000000 386.090000 ;
        RECT 1001.000000 381.910000 1006.000000 382.090000 ;
        RECT 1001.000000 389.910000 1006.000000 390.090000 ;
        RECT 1001.000000 393.910000 1006.000000 394.090000 ;
        RECT 1001.000000 397.910000 1006.000000 398.090000 ;
        RECT 1001.000000 401.910000 1006.000000 402.090000 ;
        RECT 1001.000000 405.910000 1006.000000 406.090000 ;
        RECT 1001.000000 409.910000 1006.000000 410.090000 ;
        RECT 1001.000000 413.910000 1006.000000 414.090000 ;
        RECT 901.000000 417.910000 906.000000 418.090000 ;
        RECT 901.000000 425.910000 906.000000 426.090000 ;
        RECT 901.000000 421.910000 906.000000 422.090000 ;
        RECT 901.000000 429.910000 906.000000 430.090000 ;
        RECT 901.000000 433.910000 906.000000 434.090000 ;
        RECT 901.000000 437.910000 906.000000 438.090000 ;
        RECT 901.000000 441.910000 906.000000 442.090000 ;
        RECT 951.000000 433.910000 956.000000 434.090000 ;
        RECT 951.000000 429.910000 956.000000 430.090000 ;
        RECT 951.000000 425.910000 956.000000 426.090000 ;
        RECT 951.000000 421.910000 956.000000 422.090000 ;
        RECT 951.000000 417.910000 956.000000 418.090000 ;
        RECT 951.000000 437.910000 956.000000 438.090000 ;
        RECT 951.000000 441.910000 956.000000 442.090000 ;
        RECT 1001.000000 425.910000 1006.000000 426.090000 ;
        RECT 1001.000000 421.910000 1006.000000 422.090000 ;
        RECT 1001.000000 417.910000 1006.000000 418.090000 ;
        RECT 1001.000000 429.910000 1006.000000 430.090000 ;
        RECT 1001.000000 433.910000 1006.000000 434.090000 ;
        RECT 1001.000000 437.910000 1006.000000 438.090000 ;
        RECT 1001.000000 441.910000 1006.000000 442.090000 ;
        RECT 1051.000000 357.910000 1056.000000 358.090000 ;
        RECT 1051.000000 353.910000 1056.000000 354.090000 ;
        RECT 1051.000000 349.910000 1056.000000 350.090000 ;
        RECT 1051.000000 345.910000 1056.000000 346.090000 ;
        RECT 1051.000000 369.910000 1056.000000 370.090000 ;
        RECT 1051.000000 365.910000 1056.000000 366.090000 ;
        RECT 1051.000000 361.910000 1056.000000 362.090000 ;
        RECT 1051.000000 373.910000 1056.000000 374.090000 ;
        RECT 1051.000000 377.910000 1056.000000 378.090000 ;
        RECT 1101.000000 345.910000 1106.000000 346.090000 ;
        RECT 1101.000000 349.910000 1106.000000 350.090000 ;
        RECT 1101.000000 353.910000 1106.000000 354.090000 ;
        RECT 1101.000000 357.910000 1106.000000 358.090000 ;
        RECT 1101.000000 369.910000 1106.000000 370.090000 ;
        RECT 1101.000000 365.910000 1106.000000 366.090000 ;
        RECT 1101.000000 361.910000 1106.000000 362.090000 ;
        RECT 1101.000000 377.910000 1106.000000 378.090000 ;
        RECT 1101.000000 373.910000 1106.000000 374.090000 ;
        RECT 1051.000000 397.910000 1056.000000 398.090000 ;
        RECT 1051.000000 393.910000 1056.000000 394.090000 ;
        RECT 1051.000000 389.910000 1056.000000 390.090000 ;
        RECT 1051.000000 381.910000 1056.000000 382.090000 ;
        RECT 1051.000000 385.910000 1056.000000 386.090000 ;
        RECT 1051.000000 405.910000 1056.000000 406.090000 ;
        RECT 1051.000000 401.910000 1056.000000 402.090000 ;
        RECT 1051.000000 413.910000 1056.000000 414.090000 ;
        RECT 1051.000000 409.910000 1056.000000 410.090000 ;
        RECT 1101.000000 397.910000 1106.000000 398.090000 ;
        RECT 1101.000000 393.910000 1106.000000 394.090000 ;
        RECT 1101.000000 389.910000 1106.000000 390.090000 ;
        RECT 1101.000000 381.910000 1106.000000 382.090000 ;
        RECT 1101.000000 385.910000 1106.000000 386.090000 ;
        RECT 1101.000000 405.910000 1106.000000 406.090000 ;
        RECT 1101.000000 401.910000 1106.000000 402.090000 ;
        RECT 1101.000000 413.910000 1106.000000 414.090000 ;
        RECT 1101.000000 409.910000 1106.000000 410.090000 ;
        RECT 1151.000000 357.910000 1156.000000 358.090000 ;
        RECT 1151.000000 353.910000 1156.000000 354.090000 ;
        RECT 1151.000000 349.910000 1156.000000 350.090000 ;
        RECT 1151.000000 345.910000 1156.000000 346.090000 ;
        RECT 1172.000000 357.910000 1182.000000 358.090000 ;
        RECT 1172.000000 353.910000 1182.000000 354.090000 ;
        RECT 1172.000000 349.910000 1182.000000 350.090000 ;
        RECT 1172.000000 345.910000 1182.000000 346.090000 ;
        RECT 1151.000000 365.910000 1156.000000 366.090000 ;
        RECT 1151.000000 361.910000 1156.000000 362.090000 ;
        RECT 1151.000000 369.910000 1156.000000 370.090000 ;
        RECT 1151.000000 377.910000 1156.000000 378.090000 ;
        RECT 1151.000000 373.910000 1156.000000 374.090000 ;
        RECT 1172.000000 369.910000 1182.000000 370.090000 ;
        RECT 1172.000000 365.910000 1182.000000 366.090000 ;
        RECT 1172.000000 361.910000 1182.000000 362.090000 ;
        RECT 1172.000000 373.910000 1182.000000 374.090000 ;
        RECT 1172.000000 377.910000 1182.000000 378.090000 ;
        RECT 1151.000000 385.910000 1156.000000 386.090000 ;
        RECT 1151.000000 381.910000 1156.000000 382.090000 ;
        RECT 1151.000000 389.910000 1156.000000 390.090000 ;
        RECT 1151.000000 393.910000 1156.000000 394.090000 ;
        RECT 1151.000000 397.910000 1156.000000 398.090000 ;
        RECT 1172.000000 385.910000 1182.000000 386.090000 ;
        RECT 1172.000000 381.910000 1182.000000 382.090000 ;
        RECT 1172.000000 389.910000 1182.000000 390.090000 ;
        RECT 1172.000000 393.910000 1182.000000 394.090000 ;
        RECT 1172.000000 397.910000 1182.000000 398.090000 ;
        RECT 1151.000000 405.910000 1156.000000 406.090000 ;
        RECT 1151.000000 401.910000 1156.000000 402.090000 ;
        RECT 1151.000000 409.910000 1156.000000 410.090000 ;
        RECT 1151.000000 413.910000 1156.000000 414.090000 ;
        RECT 1172.000000 405.910000 1182.000000 406.090000 ;
        RECT 1172.000000 401.910000 1182.000000 402.090000 ;
        RECT 1172.000000 409.910000 1182.000000 410.090000 ;
        RECT 1172.000000 413.910000 1182.000000 414.090000 ;
        RECT 1051.000000 425.910000 1056.000000 426.090000 ;
        RECT 1051.000000 417.910000 1056.000000 418.090000 ;
        RECT 1051.000000 421.910000 1056.000000 422.090000 ;
        RECT 1051.000000 429.910000 1056.000000 430.090000 ;
        RECT 1051.000000 433.910000 1056.000000 434.090000 ;
        RECT 1051.000000 437.910000 1056.000000 438.090000 ;
        RECT 1051.000000 441.910000 1056.000000 442.090000 ;
        RECT 1101.000000 433.910000 1106.000000 434.090000 ;
        RECT 1101.000000 429.910000 1106.000000 430.090000 ;
        RECT 1101.000000 425.910000 1106.000000 426.090000 ;
        RECT 1101.000000 421.910000 1106.000000 422.090000 ;
        RECT 1101.000000 417.910000 1106.000000 418.090000 ;
        RECT 1101.000000 441.910000 1106.000000 442.090000 ;
        RECT 1101.000000 437.910000 1106.000000 438.090000 ;
        RECT 1151.000000 417.910000 1156.000000 418.090000 ;
        RECT 1151.000000 421.910000 1156.000000 422.090000 ;
        RECT 1151.000000 425.910000 1156.000000 426.090000 ;
        RECT 1151.000000 429.910000 1156.000000 430.090000 ;
        RECT 1151.000000 433.910000 1156.000000 434.090000 ;
        RECT 1172.000000 425.910000 1182.000000 426.090000 ;
        RECT 1172.000000 417.910000 1182.000000 418.090000 ;
        RECT 1172.000000 421.910000 1182.000000 422.090000 ;
        RECT 1172.000000 429.910000 1182.000000 430.090000 ;
        RECT 1172.000000 433.910000 1182.000000 434.090000 ;
        RECT 1151.000000 437.910000 1156.000000 438.090000 ;
        RECT 1151.000000 441.910000 1156.000000 442.090000 ;
        RECT 1151.000000 453.910000 1156.000000 454.090000 ;
        RECT 1151.000000 449.910000 1156.000000 450.090000 ;
        RECT 1151.000000 445.910000 1156.000000 446.090000 ;
        RECT 1172.000000 437.910000 1182.000000 438.090000 ;
        RECT 1172.000000 441.910000 1182.000000 442.090000 ;
        RECT 1151.000000 461.910000 1156.000000 462.090000 ;
        RECT 1151.000000 457.910000 1156.000000 458.090000 ;
        RECT 1151.000000 465.910000 1156.000000 466.090000 ;
        RECT 1151.000000 469.910000 1156.000000 470.090000 ;
        RECT 1151.000000 481.910000 1156.000000 482.090000 ;
        RECT 1151.000000 477.910000 1156.000000 478.090000 ;
        RECT 1151.000000 473.910000 1156.000000 474.090000 ;
        RECT 1151.000000 489.910000 1156.000000 490.090000 ;
        RECT 1151.000000 485.910000 1156.000000 486.090000 ;
        RECT 1151.000000 493.910000 1156.000000 494.090000 ;
        RECT 1151.000000 497.910000 1156.000000 498.090000 ;
        RECT 1151.000000 505.910000 1156.000000 506.090000 ;
        RECT 1151.000000 501.910000 1156.000000 502.090000 ;
        RECT 1151.000000 509.910000 1156.000000 510.090000 ;
        RECT 1151.000000 513.910000 1156.000000 514.090000 ;
        RECT 1151.000000 517.910000 1156.000000 518.090000 ;
        RECT 1151.000000 521.910000 1156.000000 522.090000 ;
        RECT 1151.000000 525.910000 1156.000000 526.090000 ;
        RECT 1151.000000 533.910000 1156.000000 534.090000 ;
        RECT 1151.000000 529.910000 1156.000000 530.090000 ;
        RECT 1151.000000 545.910000 1156.000000 546.090000 ;
        RECT 1151.000000 537.910000 1156.000000 538.090000 ;
        RECT 1151.000000 541.910000 1156.000000 542.090000 ;
        RECT 1151.000000 549.910000 1156.000000 550.090000 ;
        RECT 1151.000000 553.910000 1156.000000 554.090000 ;
        RECT 1151.000000 561.910000 1156.000000 562.090000 ;
        RECT 1151.000000 557.910000 1156.000000 558.090000 ;
        RECT 1151.000000 565.910000 1156.000000 566.090000 ;
        RECT 1151.000000 569.910000 1156.000000 570.090000 ;
        RECT 1151.000000 573.910000 1156.000000 574.090000 ;
        RECT 1151.000000 577.910000 1156.000000 578.090000 ;
        RECT 1151.000000 581.910000 1156.000000 582.090000 ;
        RECT 1151.000000 585.910000 1156.000000 586.090000 ;
        RECT 1151.000000 589.910000 1156.000000 590.090000 ;
        RECT 1151.000000 593.910000 1156.000000 594.090000 ;
        RECT 1151.000000 597.910000 1156.000000 598.090000 ;
        RECT 1151.000000 601.910000 1156.000000 602.090000 ;
        RECT 1151.000000 609.910000 1156.000000 610.090000 ;
        RECT 1151.000000 605.910000 1156.000000 606.090000 ;
        RECT 1151.000000 613.910000 1156.000000 614.090000 ;
        RECT 1151.000000 617.910000 1156.000000 618.090000 ;
        RECT 1151.000000 621.910000 1156.000000 622.090000 ;
        RECT 1151.000000 625.910000 1156.000000 626.090000 ;
        RECT 1151.000000 629.910000 1156.000000 630.090000 ;
        RECT 1151.000000 637.910000 1156.000000 638.090000 ;
        RECT 1151.000000 633.910000 1156.000000 634.090000 ;
        RECT 601.000000 657.910000 606.000000 658.090000 ;
        RECT 601.000000 673.910000 606.000000 674.090000 ;
        RECT 601.000000 669.910000 606.000000 670.090000 ;
        RECT 601.000000 665.910000 606.000000 666.090000 ;
        RECT 601.000000 661.910000 606.000000 662.090000 ;
        RECT 651.000000 657.910000 656.000000 658.090000 ;
        RECT 651.000000 661.910000 656.000000 662.090000 ;
        RECT 651.000000 665.910000 656.000000 666.090000 ;
        RECT 651.000000 673.910000 656.000000 674.090000 ;
        RECT 651.000000 669.910000 656.000000 670.090000 ;
        RECT 601.000000 677.910000 606.000000 678.090000 ;
        RECT 601.000000 681.910000 606.000000 682.090000 ;
        RECT 651.000000 677.910000 656.000000 678.090000 ;
        RECT 651.000000 681.910000 656.000000 682.090000 ;
        RECT 1151.000000 657.910000 1156.000000 658.090000 ;
        RECT 1151.000000 641.910000 1156.000000 642.090000 ;
        RECT 1151.000000 645.910000 1156.000000 646.090000 ;
        RECT 1151.000000 653.910000 1156.000000 654.090000 ;
        RECT 1151.000000 649.910000 1156.000000 650.090000 ;
        RECT 1151.000000 665.910000 1156.000000 666.090000 ;
        RECT 1151.000000 661.910000 1156.000000 662.090000 ;
        RECT 1151.000000 669.910000 1156.000000 670.090000 ;
        RECT 1151.000000 673.910000 1156.000000 674.090000 ;
        RECT 1151.000000 681.910000 1156.000000 682.090000 ;
        RECT 1151.000000 677.910000 1156.000000 678.090000 ;
    END
# end of P/G power stripe data as pin

  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M7 ;
        RECT 60.000000 0.000000 65.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 60.000000 681.000000 65.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 110.000000 0.000000 115.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 110.000000 681.000000 115.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 160.000000 0.000000 165.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 210.000000 0.000000 215.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 260.000000 0.000000 265.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 260.000000 681.000000 265.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 310.000000 0.000000 315.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 310.000000 681.000000 315.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 360.000000 0.000000 365.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 360.000000 681.000000 365.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 410.000000 0.000000 415.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 410.000000 501.000000 415.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 410.000000 656.000000 415.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 410.000000 681.000000 415.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 460.000000 0.000000 465.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 460.000000 501.000000 465.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 460.000000 656.000000 465.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 460.000000 681.000000 465.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 510.000000 0.000000 515.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 510.000000 501.000000 515.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 510.000000 656.000000 515.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 510.000000 681.000000 515.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 560.000000 0.000000 565.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 560.000000 501.000000 565.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 560.000000 656.000000 565.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 560.000000 681.000000 565.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 610.000000 0.000000 615.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 610.000000 501.000000 615.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 610.000000 656.000000 615.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 610.000000 681.000000 615.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 660.000000 0.000000 665.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 660.000000 501.000000 665.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 660.000000 656.000000 665.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 660.000000 681.000000 665.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 710.000000 0.000000 715.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 710.000000 501.000000 715.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 760.000000 0.000000 765.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 760.000000 441.000000 765.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 810.000000 0.000000 815.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 810.000000 441.000000 815.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 860.000000 0.000000 865.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 860.000000 441.000000 865.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 910.000000 0.000000 915.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 910.000000 441.000000 915.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 960.000000 0.000000 965.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 960.000000 441.000000 965.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1010.000000 0.000000 1015.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1010.000000 441.000000 1015.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1060.000000 0.000000 1065.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1060.000000 441.000000 1065.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1110.000000 0.000000 1115.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1110.000000 441.000000 1115.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1160.000000 0.000000 1165.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1160.000000 681.000000 1165.000000 686.000000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER M2 ;
        RECT 60.000000 3.910000 65.000000 4.090000 ;
        RECT 60.000000 7.910000 65.000000 8.090000 ;
        RECT 110.000000 7.910000 115.000000 8.090000 ;
        RECT 110.000000 3.910000 115.000000 4.090000 ;
        RECT 160.000000 7.910000 165.000000 8.090000 ;
        RECT 160.000000 3.910000 165.000000 4.090000 ;
        RECT 210.000000 7.910000 215.000000 8.090000 ;
        RECT 210.000000 3.910000 215.000000 4.090000 ;
        RECT 260.000000 7.910000 265.000000 8.090000 ;
        RECT 260.000000 3.910000 265.000000 4.090000 ;
        RECT 310.000000 7.910000 315.000000 8.090000 ;
        RECT 310.000000 3.910000 315.000000 4.090000 ;
        RECT 360.000000 7.910000 365.000000 8.090000 ;
        RECT 360.000000 3.910000 365.000000 4.090000 ;
        RECT 410.000000 7.910000 415.000000 8.090000 ;
        RECT 410.000000 3.910000 415.000000 4.090000 ;
        RECT 460.000000 7.910000 465.000000 8.090000 ;
        RECT 460.000000 3.910000 465.000000 4.090000 ;
        RECT 510.000000 7.910000 515.000000 8.090000 ;
        RECT 510.000000 3.910000 515.000000 4.090000 ;
        RECT 560.000000 7.910000 565.000000 8.090000 ;
        RECT 560.000000 3.910000 565.000000 4.090000 ;
        RECT 18.000000 267.910000 28.000000 268.090000 ;
        RECT 18.000000 259.910000 28.000000 260.090000 ;
        RECT 18.000000 263.910000 28.000000 264.090000 ;
        RECT 60.000000 267.910000 65.000000 268.090000 ;
        RECT 60.000000 263.910000 65.000000 264.090000 ;
        RECT 60.000000 259.910000 65.000000 260.090000 ;
        RECT 110.000000 267.910000 115.000000 268.090000 ;
        RECT 110.000000 259.910000 115.000000 260.090000 ;
        RECT 110.000000 263.910000 115.000000 264.090000 ;
        RECT 18.000000 283.910000 28.000000 284.090000 ;
        RECT 18.000000 279.910000 28.000000 280.090000 ;
        RECT 18.000000 275.910000 28.000000 276.090000 ;
        RECT 18.000000 271.910000 28.000000 272.090000 ;
        RECT 18.000000 287.910000 28.000000 288.090000 ;
        RECT 18.000000 291.910000 28.000000 292.090000 ;
        RECT 18.000000 295.910000 28.000000 296.090000 ;
        RECT 18.000000 299.910000 28.000000 300.090000 ;
        RECT 18.000000 303.910000 28.000000 304.090000 ;
        RECT 60.000000 283.910000 65.000000 284.090000 ;
        RECT 60.000000 279.910000 65.000000 280.090000 ;
        RECT 60.000000 275.910000 65.000000 276.090000 ;
        RECT 60.000000 271.910000 65.000000 272.090000 ;
        RECT 60.000000 287.910000 65.000000 288.090000 ;
        RECT 60.000000 291.910000 65.000000 292.090000 ;
        RECT 60.000000 295.910000 65.000000 296.090000 ;
        RECT 60.000000 299.910000 65.000000 300.090000 ;
        RECT 60.000000 303.910000 65.000000 304.090000 ;
        RECT 18.000000 307.910000 28.000000 308.090000 ;
        RECT 18.000000 311.910000 28.000000 312.090000 ;
        RECT 18.000000 315.910000 28.000000 316.090000 ;
        RECT 18.000000 319.910000 28.000000 320.090000 ;
        RECT 18.000000 323.910000 28.000000 324.090000 ;
        RECT 18.000000 339.910000 28.000000 340.090000 ;
        RECT 18.000000 335.910000 28.000000 336.090000 ;
        RECT 18.000000 331.910000 28.000000 332.090000 ;
        RECT 18.000000 327.910000 28.000000 328.090000 ;
        RECT 60.000000 307.910000 65.000000 308.090000 ;
        RECT 60.000000 311.910000 65.000000 312.090000 ;
        RECT 60.000000 315.910000 65.000000 316.090000 ;
        RECT 60.000000 319.910000 65.000000 320.090000 ;
        RECT 60.000000 323.910000 65.000000 324.090000 ;
        RECT 60.000000 339.910000 65.000000 340.090000 ;
        RECT 60.000000 335.910000 65.000000 336.090000 ;
        RECT 60.000000 331.910000 65.000000 332.090000 ;
        RECT 60.000000 327.910000 65.000000 328.090000 ;
        RECT 110.000000 271.910000 115.000000 272.090000 ;
        RECT 110.000000 275.910000 115.000000 276.090000 ;
        RECT 110.000000 279.910000 115.000000 280.090000 ;
        RECT 110.000000 283.910000 115.000000 284.090000 ;
        RECT 110.000000 287.910000 115.000000 288.090000 ;
        RECT 110.000000 291.910000 115.000000 292.090000 ;
        RECT 110.000000 295.910000 115.000000 296.090000 ;
        RECT 110.000000 299.910000 115.000000 300.090000 ;
        RECT 110.000000 303.910000 115.000000 304.090000 ;
        RECT 110.000000 311.910000 115.000000 312.090000 ;
        RECT 110.000000 307.910000 115.000000 308.090000 ;
        RECT 110.000000 323.910000 115.000000 324.090000 ;
        RECT 110.000000 319.910000 115.000000 320.090000 ;
        RECT 110.000000 315.910000 115.000000 316.090000 ;
        RECT 110.000000 339.910000 115.000000 340.090000 ;
        RECT 110.000000 335.910000 115.000000 336.090000 ;
        RECT 110.000000 331.910000 115.000000 332.090000 ;
        RECT 110.000000 327.910000 115.000000 328.090000 ;
        RECT 160.000000 259.910000 165.000000 260.090000 ;
        RECT 160.000000 263.910000 165.000000 264.090000 ;
        RECT 160.000000 267.910000 165.000000 268.090000 ;
        RECT 210.000000 267.910000 215.000000 268.090000 ;
        RECT 210.000000 263.910000 215.000000 264.090000 ;
        RECT 210.000000 259.910000 215.000000 260.090000 ;
        RECT 260.000000 267.910000 265.000000 268.090000 ;
        RECT 260.000000 259.910000 265.000000 260.090000 ;
        RECT 260.000000 263.910000 265.000000 264.090000 ;
        RECT 160.000000 271.910000 165.000000 272.090000 ;
        RECT 160.000000 275.910000 165.000000 276.090000 ;
        RECT 160.000000 283.910000 165.000000 284.090000 ;
        RECT 160.000000 279.910000 165.000000 280.090000 ;
        RECT 160.000000 287.910000 165.000000 288.090000 ;
        RECT 160.000000 291.910000 165.000000 292.090000 ;
        RECT 160.000000 295.910000 165.000000 296.090000 ;
        RECT 160.000000 303.910000 165.000000 304.090000 ;
        RECT 160.000000 299.910000 165.000000 300.090000 ;
        RECT 210.000000 283.910000 215.000000 284.090000 ;
        RECT 210.000000 279.910000 215.000000 280.090000 ;
        RECT 210.000000 275.910000 215.000000 276.090000 ;
        RECT 210.000000 271.910000 215.000000 272.090000 ;
        RECT 210.000000 287.910000 215.000000 288.090000 ;
        RECT 210.000000 291.910000 215.000000 292.090000 ;
        RECT 210.000000 295.910000 215.000000 296.090000 ;
        RECT 210.000000 299.910000 215.000000 300.090000 ;
        RECT 210.000000 303.910000 215.000000 304.090000 ;
        RECT 160.000000 311.910000 165.000000 312.090000 ;
        RECT 160.000000 307.910000 165.000000 308.090000 ;
        RECT 160.000000 315.910000 165.000000 316.090000 ;
        RECT 160.000000 319.910000 165.000000 320.090000 ;
        RECT 160.000000 323.910000 165.000000 324.090000 ;
        RECT 160.000000 331.910000 165.000000 332.090000 ;
        RECT 160.000000 327.910000 165.000000 328.090000 ;
        RECT 160.000000 335.910000 165.000000 336.090000 ;
        RECT 160.000000 339.910000 165.000000 340.090000 ;
        RECT 210.000000 307.910000 215.000000 308.090000 ;
        RECT 210.000000 311.910000 215.000000 312.090000 ;
        RECT 210.000000 315.910000 215.000000 316.090000 ;
        RECT 210.000000 319.910000 215.000000 320.090000 ;
        RECT 210.000000 323.910000 215.000000 324.090000 ;
        RECT 210.000000 327.910000 215.000000 328.090000 ;
        RECT 210.000000 331.910000 215.000000 332.090000 ;
        RECT 210.000000 335.910000 215.000000 336.090000 ;
        RECT 210.000000 339.910000 215.000000 340.090000 ;
        RECT 260.000000 271.910000 265.000000 272.090000 ;
        RECT 260.000000 275.910000 265.000000 276.090000 ;
        RECT 260.000000 279.910000 265.000000 280.090000 ;
        RECT 260.000000 283.910000 265.000000 284.090000 ;
        RECT 260.000000 291.910000 265.000000 292.090000 ;
        RECT 260.000000 287.910000 265.000000 288.090000 ;
        RECT 260.000000 295.910000 265.000000 296.090000 ;
        RECT 260.000000 299.910000 265.000000 300.090000 ;
        RECT 260.000000 303.910000 265.000000 304.090000 ;
        RECT 260.000000 311.910000 265.000000 312.090000 ;
        RECT 260.000000 307.910000 265.000000 308.090000 ;
        RECT 260.000000 323.910000 265.000000 324.090000 ;
        RECT 260.000000 319.910000 265.000000 320.090000 ;
        RECT 260.000000 315.910000 265.000000 316.090000 ;
        RECT 260.000000 331.910000 265.000000 332.090000 ;
        RECT 260.000000 327.910000 265.000000 328.090000 ;
        RECT 260.000000 339.910000 265.000000 340.090000 ;
        RECT 260.000000 335.910000 265.000000 336.090000 ;
        RECT 310.000000 259.910000 315.000000 260.090000 ;
        RECT 310.000000 263.910000 315.000000 264.090000 ;
        RECT 310.000000 267.910000 315.000000 268.090000 ;
        RECT 360.000000 267.910000 365.000000 268.090000 ;
        RECT 360.000000 263.910000 365.000000 264.090000 ;
        RECT 360.000000 259.910000 365.000000 260.090000 ;
        RECT 410.000000 267.910000 415.000000 268.090000 ;
        RECT 410.000000 259.910000 415.000000 260.090000 ;
        RECT 410.000000 263.910000 415.000000 264.090000 ;
        RECT 310.000000 271.910000 315.000000 272.090000 ;
        RECT 310.000000 275.910000 315.000000 276.090000 ;
        RECT 310.000000 279.910000 315.000000 280.090000 ;
        RECT 310.000000 283.910000 315.000000 284.090000 ;
        RECT 310.000000 291.910000 315.000000 292.090000 ;
        RECT 310.000000 287.910000 315.000000 288.090000 ;
        RECT 310.000000 295.910000 315.000000 296.090000 ;
        RECT 310.000000 299.910000 315.000000 300.090000 ;
        RECT 310.000000 303.910000 315.000000 304.090000 ;
        RECT 360.000000 283.910000 365.000000 284.090000 ;
        RECT 360.000000 279.910000 365.000000 280.090000 ;
        RECT 360.000000 275.910000 365.000000 276.090000 ;
        RECT 360.000000 271.910000 365.000000 272.090000 ;
        RECT 360.000000 287.910000 365.000000 288.090000 ;
        RECT 360.000000 291.910000 365.000000 292.090000 ;
        RECT 360.000000 295.910000 365.000000 296.090000 ;
        RECT 360.000000 299.910000 365.000000 300.090000 ;
        RECT 360.000000 303.910000 365.000000 304.090000 ;
        RECT 310.000000 307.910000 315.000000 308.090000 ;
        RECT 310.000000 311.910000 315.000000 312.090000 ;
        RECT 310.000000 315.910000 315.000000 316.090000 ;
        RECT 310.000000 323.910000 315.000000 324.090000 ;
        RECT 310.000000 319.910000 315.000000 320.090000 ;
        RECT 310.000000 327.910000 315.000000 328.090000 ;
        RECT 310.000000 331.910000 315.000000 332.090000 ;
        RECT 310.000000 335.910000 315.000000 336.090000 ;
        RECT 310.000000 339.910000 315.000000 340.090000 ;
        RECT 360.000000 307.910000 365.000000 308.090000 ;
        RECT 360.000000 311.910000 365.000000 312.090000 ;
        RECT 360.000000 315.910000 365.000000 316.090000 ;
        RECT 360.000000 319.910000 365.000000 320.090000 ;
        RECT 360.000000 323.910000 365.000000 324.090000 ;
        RECT 360.000000 339.910000 365.000000 340.090000 ;
        RECT 360.000000 335.910000 365.000000 336.090000 ;
        RECT 360.000000 331.910000 365.000000 332.090000 ;
        RECT 360.000000 327.910000 365.000000 328.090000 ;
        RECT 410.000000 271.910000 415.000000 272.090000 ;
        RECT 410.000000 275.910000 415.000000 276.090000 ;
        RECT 410.000000 279.910000 415.000000 280.090000 ;
        RECT 410.000000 283.910000 415.000000 284.090000 ;
        RECT 410.000000 295.910000 415.000000 296.090000 ;
        RECT 410.000000 291.910000 415.000000 292.090000 ;
        RECT 410.000000 287.910000 415.000000 288.090000 ;
        RECT 410.000000 299.910000 415.000000 300.090000 ;
        RECT 410.000000 303.910000 415.000000 304.090000 ;
        RECT 410.000000 307.910000 415.000000 308.090000 ;
        RECT 410.000000 311.910000 415.000000 312.090000 ;
        RECT 410.000000 315.910000 415.000000 316.090000 ;
        RECT 410.000000 319.910000 415.000000 320.090000 ;
        RECT 410.000000 323.910000 415.000000 324.090000 ;
        RECT 410.000000 327.910000 415.000000 328.090000 ;
        RECT 410.000000 331.910000 415.000000 332.090000 ;
        RECT 410.000000 335.910000 415.000000 336.090000 ;
        RECT 410.000000 339.910000 415.000000 340.090000 ;
        RECT 460.000000 267.910000 465.000000 268.090000 ;
        RECT 460.000000 263.910000 465.000000 264.090000 ;
        RECT 460.000000 259.910000 465.000000 260.090000 ;
        RECT 510.000000 259.910000 515.000000 260.090000 ;
        RECT 510.000000 263.910000 515.000000 264.090000 ;
        RECT 510.000000 267.910000 515.000000 268.090000 ;
        RECT 560.000000 267.910000 565.000000 268.090000 ;
        RECT 560.000000 259.910000 565.000000 260.090000 ;
        RECT 560.000000 263.910000 565.000000 264.090000 ;
        RECT 460.000000 283.910000 465.000000 284.090000 ;
        RECT 460.000000 279.910000 465.000000 280.090000 ;
        RECT 460.000000 275.910000 465.000000 276.090000 ;
        RECT 460.000000 271.910000 465.000000 272.090000 ;
        RECT 460.000000 295.910000 465.000000 296.090000 ;
        RECT 460.000000 291.910000 465.000000 292.090000 ;
        RECT 460.000000 287.910000 465.000000 288.090000 ;
        RECT 510.000000 271.910000 515.000000 272.090000 ;
        RECT 510.000000 275.910000 515.000000 276.090000 ;
        RECT 510.000000 283.910000 515.000000 284.090000 ;
        RECT 510.000000 279.910000 515.000000 280.090000 ;
        RECT 510.000000 287.910000 515.000000 288.090000 ;
        RECT 510.000000 291.910000 515.000000 292.090000 ;
        RECT 510.000000 295.910000 515.000000 296.090000 ;
        RECT 510.000000 303.910000 515.000000 304.090000 ;
        RECT 510.000000 299.910000 515.000000 300.090000 ;
        RECT 460.000000 319.910000 465.000000 320.090000 ;
        RECT 460.000000 323.910000 465.000000 324.090000 ;
        RECT 460.000000 339.910000 465.000000 340.090000 ;
        RECT 460.000000 335.910000 465.000000 336.090000 ;
        RECT 460.000000 331.910000 465.000000 332.090000 ;
        RECT 460.000000 327.910000 465.000000 328.090000 ;
        RECT 510.000000 311.910000 515.000000 312.090000 ;
        RECT 510.000000 307.910000 515.000000 308.090000 ;
        RECT 510.000000 315.910000 515.000000 316.090000 ;
        RECT 510.000000 319.910000 515.000000 320.090000 ;
        RECT 510.000000 323.910000 515.000000 324.090000 ;
        RECT 510.000000 331.910000 515.000000 332.090000 ;
        RECT 510.000000 327.910000 515.000000 328.090000 ;
        RECT 510.000000 335.910000 515.000000 336.090000 ;
        RECT 510.000000 339.910000 515.000000 340.090000 ;
        RECT 560.000000 275.910000 565.000000 276.090000 ;
        RECT 560.000000 271.910000 565.000000 272.090000 ;
        RECT 560.000000 283.910000 565.000000 284.090000 ;
        RECT 560.000000 279.910000 565.000000 280.090000 ;
        RECT 560.000000 295.910000 565.000000 296.090000 ;
        RECT 560.000000 291.910000 565.000000 292.090000 ;
        RECT 560.000000 287.910000 565.000000 288.090000 ;
        RECT 560.000000 303.910000 565.000000 304.090000 ;
        RECT 560.000000 299.910000 565.000000 300.090000 ;
        RECT 560.000000 307.910000 565.000000 308.090000 ;
        RECT 560.000000 311.910000 565.000000 312.090000 ;
        RECT 560.000000 315.910000 565.000000 316.090000 ;
        RECT 560.000000 319.910000 565.000000 320.090000 ;
        RECT 560.000000 323.910000 565.000000 324.090000 ;
        RECT 560.000000 327.910000 565.000000 328.090000 ;
        RECT 560.000000 331.910000 565.000000 332.090000 ;
        RECT 560.000000 339.910000 565.000000 340.090000 ;
        RECT 560.000000 335.910000 565.000000 336.090000 ;
        RECT 610.000000 3.910000 615.000000 4.090000 ;
        RECT 610.000000 7.910000 615.000000 8.090000 ;
        RECT 660.000000 7.910000 665.000000 8.090000 ;
        RECT 660.000000 3.910000 665.000000 4.090000 ;
        RECT 710.000000 7.910000 715.000000 8.090000 ;
        RECT 710.000000 3.910000 715.000000 4.090000 ;
        RECT 760.000000 7.910000 765.000000 8.090000 ;
        RECT 760.000000 3.910000 765.000000 4.090000 ;
        RECT 810.000000 7.910000 815.000000 8.090000 ;
        RECT 810.000000 3.910000 815.000000 4.090000 ;
        RECT 860.000000 7.910000 865.000000 8.090000 ;
        RECT 860.000000 3.910000 865.000000 4.090000 ;
        RECT 960.000000 7.910000 965.000000 8.090000 ;
        RECT 960.000000 3.910000 965.000000 4.090000 ;
        RECT 910.000000 7.910000 915.000000 8.090000 ;
        RECT 910.000000 3.910000 915.000000 4.090000 ;
        RECT 1010.000000 7.910000 1015.000000 8.090000 ;
        RECT 1010.000000 3.910000 1015.000000 4.090000 ;
        RECT 1110.000000 7.910000 1115.000000 8.090000 ;
        RECT 1110.000000 3.910000 1115.000000 4.090000 ;
        RECT 1060.000000 7.910000 1065.000000 8.090000 ;
        RECT 1060.000000 3.910000 1065.000000 4.090000 ;
        RECT 1160.000000 3.910000 1165.000000 4.090000 ;
        RECT 1160.000000 7.910000 1165.000000 8.090000 ;
        RECT 1158.000000 27.910000 1168.000000 28.090000 ;
        RECT 1158.000000 23.910000 1168.000000 24.090000 ;
        RECT 1158.000000 19.910000 1168.000000 20.090000 ;
        RECT 1160.000000 15.910000 1165.000000 16.090000 ;
        RECT 1160.000000 11.910000 1165.000000 12.090000 ;
        RECT 1158.000000 31.910000 1168.000000 32.090000 ;
        RECT 1158.000000 35.910000 1168.000000 36.090000 ;
        RECT 1158.000000 43.910000 1168.000000 44.090000 ;
        RECT 1158.000000 39.910000 1168.000000 40.090000 ;
        RECT 610.000000 263.910000 615.000000 264.090000 ;
        RECT 610.000000 259.910000 615.000000 260.090000 ;
        RECT 610.000000 267.910000 615.000000 268.090000 ;
        RECT 660.000000 259.910000 665.000000 260.090000 ;
        RECT 660.000000 263.910000 665.000000 264.090000 ;
        RECT 660.000000 267.910000 665.000000 268.090000 ;
        RECT 710.000000 267.910000 715.000000 268.090000 ;
        RECT 710.000000 259.910000 715.000000 260.090000 ;
        RECT 710.000000 263.910000 715.000000 264.090000 ;
        RECT 610.000000 271.910000 615.000000 272.090000 ;
        RECT 610.000000 275.910000 615.000000 276.090000 ;
        RECT 610.000000 279.910000 615.000000 280.090000 ;
        RECT 610.000000 283.910000 615.000000 284.090000 ;
        RECT 610.000000 287.910000 615.000000 288.090000 ;
        RECT 610.000000 291.910000 615.000000 292.090000 ;
        RECT 610.000000 295.910000 615.000000 296.090000 ;
        RECT 610.000000 299.910000 615.000000 300.090000 ;
        RECT 610.000000 303.910000 615.000000 304.090000 ;
        RECT 660.000000 271.910000 665.000000 272.090000 ;
        RECT 660.000000 275.910000 665.000000 276.090000 ;
        RECT 660.000000 283.910000 665.000000 284.090000 ;
        RECT 660.000000 279.910000 665.000000 280.090000 ;
        RECT 660.000000 287.910000 665.000000 288.090000 ;
        RECT 660.000000 291.910000 665.000000 292.090000 ;
        RECT 660.000000 295.910000 665.000000 296.090000 ;
        RECT 660.000000 299.910000 665.000000 300.090000 ;
        RECT 660.000000 303.910000 665.000000 304.090000 ;
        RECT 610.000000 307.910000 615.000000 308.090000 ;
        RECT 610.000000 311.910000 615.000000 312.090000 ;
        RECT 610.000000 315.910000 615.000000 316.090000 ;
        RECT 610.000000 319.910000 615.000000 320.090000 ;
        RECT 610.000000 323.910000 615.000000 324.090000 ;
        RECT 610.000000 339.910000 615.000000 340.090000 ;
        RECT 610.000000 335.910000 615.000000 336.090000 ;
        RECT 610.000000 331.910000 615.000000 332.090000 ;
        RECT 610.000000 327.910000 615.000000 328.090000 ;
        RECT 660.000000 311.910000 665.000000 312.090000 ;
        RECT 660.000000 307.910000 665.000000 308.090000 ;
        RECT 660.000000 315.910000 665.000000 316.090000 ;
        RECT 660.000000 319.910000 665.000000 320.090000 ;
        RECT 660.000000 323.910000 665.000000 324.090000 ;
        RECT 660.000000 331.910000 665.000000 332.090000 ;
        RECT 660.000000 327.910000 665.000000 328.090000 ;
        RECT 660.000000 335.910000 665.000000 336.090000 ;
        RECT 660.000000 339.910000 665.000000 340.090000 ;
        RECT 710.000000 271.910000 715.000000 272.090000 ;
        RECT 710.000000 275.910000 715.000000 276.090000 ;
        RECT 710.000000 279.910000 715.000000 280.090000 ;
        RECT 710.000000 283.910000 715.000000 284.090000 ;
        RECT 710.000000 295.910000 715.000000 296.090000 ;
        RECT 710.000000 291.910000 715.000000 292.090000 ;
        RECT 710.000000 287.910000 715.000000 288.090000 ;
        RECT 710.000000 303.910000 715.000000 304.090000 ;
        RECT 710.000000 299.910000 715.000000 300.090000 ;
        RECT 710.000000 323.910000 715.000000 324.090000 ;
        RECT 710.000000 319.910000 715.000000 320.090000 ;
        RECT 710.000000 315.910000 715.000000 316.090000 ;
        RECT 710.000000 311.910000 715.000000 312.090000 ;
        RECT 710.000000 307.910000 715.000000 308.090000 ;
        RECT 710.000000 331.910000 715.000000 332.090000 ;
        RECT 710.000000 327.910000 715.000000 328.090000 ;
        RECT 710.000000 339.910000 715.000000 340.090000 ;
        RECT 710.000000 335.910000 715.000000 336.090000 ;
        RECT 760.000000 267.910000 765.000000 268.090000 ;
        RECT 760.000000 263.910000 765.000000 264.090000 ;
        RECT 760.000000 259.910000 765.000000 260.090000 ;
        RECT 810.000000 259.910000 815.000000 260.090000 ;
        RECT 810.000000 263.910000 815.000000 264.090000 ;
        RECT 810.000000 267.910000 815.000000 268.090000 ;
        RECT 860.000000 267.910000 865.000000 268.090000 ;
        RECT 860.000000 259.910000 865.000000 260.090000 ;
        RECT 860.000000 263.910000 865.000000 264.090000 ;
        RECT 760.000000 283.910000 765.000000 284.090000 ;
        RECT 760.000000 279.910000 765.000000 280.090000 ;
        RECT 760.000000 275.910000 765.000000 276.090000 ;
        RECT 760.000000 271.910000 765.000000 272.090000 ;
        RECT 760.000000 287.910000 765.000000 288.090000 ;
        RECT 760.000000 291.910000 765.000000 292.090000 ;
        RECT 760.000000 295.910000 765.000000 296.090000 ;
        RECT 760.000000 299.910000 765.000000 300.090000 ;
        RECT 760.000000 303.910000 765.000000 304.090000 ;
        RECT 810.000000 271.910000 815.000000 272.090000 ;
        RECT 810.000000 275.910000 815.000000 276.090000 ;
        RECT 810.000000 283.910000 815.000000 284.090000 ;
        RECT 810.000000 279.910000 815.000000 280.090000 ;
        RECT 810.000000 287.910000 815.000000 288.090000 ;
        RECT 810.000000 291.910000 815.000000 292.090000 ;
        RECT 810.000000 295.910000 815.000000 296.090000 ;
        RECT 810.000000 303.910000 815.000000 304.090000 ;
        RECT 810.000000 299.910000 815.000000 300.090000 ;
        RECT 760.000000 307.910000 765.000000 308.090000 ;
        RECT 760.000000 311.910000 765.000000 312.090000 ;
        RECT 760.000000 315.910000 765.000000 316.090000 ;
        RECT 760.000000 319.910000 765.000000 320.090000 ;
        RECT 760.000000 323.910000 765.000000 324.090000 ;
        RECT 760.000000 339.910000 765.000000 340.090000 ;
        RECT 760.000000 335.910000 765.000000 336.090000 ;
        RECT 760.000000 331.910000 765.000000 332.090000 ;
        RECT 760.000000 327.910000 765.000000 328.090000 ;
        RECT 810.000000 307.910000 815.000000 308.090000 ;
        RECT 810.000000 311.910000 815.000000 312.090000 ;
        RECT 810.000000 315.910000 815.000000 316.090000 ;
        RECT 810.000000 323.910000 815.000000 324.090000 ;
        RECT 810.000000 319.910000 815.000000 320.090000 ;
        RECT 810.000000 327.910000 815.000000 328.090000 ;
        RECT 810.000000 331.910000 815.000000 332.090000 ;
        RECT 810.000000 335.910000 815.000000 336.090000 ;
        RECT 810.000000 339.910000 815.000000 340.090000 ;
        RECT 860.000000 271.910000 865.000000 272.090000 ;
        RECT 860.000000 275.910000 865.000000 276.090000 ;
        RECT 860.000000 279.910000 865.000000 280.090000 ;
        RECT 860.000000 283.910000 865.000000 284.090000 ;
        RECT 860.000000 295.910000 865.000000 296.090000 ;
        RECT 860.000000 291.910000 865.000000 292.090000 ;
        RECT 860.000000 287.910000 865.000000 288.090000 ;
        RECT 860.000000 303.910000 865.000000 304.090000 ;
        RECT 860.000000 299.910000 865.000000 300.090000 ;
        RECT 860.000000 307.910000 865.000000 308.090000 ;
        RECT 860.000000 311.910000 865.000000 312.090000 ;
        RECT 860.000000 315.910000 865.000000 316.090000 ;
        RECT 860.000000 319.910000 865.000000 320.090000 ;
        RECT 860.000000 323.910000 865.000000 324.090000 ;
        RECT 860.000000 339.910000 865.000000 340.090000 ;
        RECT 860.000000 335.910000 865.000000 336.090000 ;
        RECT 860.000000 331.910000 865.000000 332.090000 ;
        RECT 860.000000 327.910000 865.000000 328.090000 ;
        RECT 1158.000000 47.910000 1168.000000 48.090000 ;
        RECT 1158.000000 51.910000 1168.000000 52.090000 ;
        RECT 1158.000000 63.910000 1168.000000 64.090000 ;
        RECT 1158.000000 59.910000 1168.000000 60.090000 ;
        RECT 1158.000000 55.910000 1168.000000 56.090000 ;
        RECT 1158.000000 67.910000 1168.000000 68.090000 ;
        RECT 1158.000000 71.910000 1168.000000 72.090000 ;
        RECT 1158.000000 79.910000 1168.000000 80.090000 ;
        RECT 1158.000000 75.910000 1168.000000 76.090000 ;
        RECT 1158.000000 83.910000 1168.000000 84.090000 ;
        RECT 1158.000000 87.910000 1168.000000 88.090000 ;
        RECT 1158.000000 91.910000 1168.000000 92.090000 ;
        RECT 1158.000000 99.910000 1168.000000 100.090000 ;
        RECT 1158.000000 95.910000 1168.000000 96.090000 ;
        RECT 1158.000000 103.910000 1168.000000 104.090000 ;
        RECT 1158.000000 107.910000 1168.000000 108.090000 ;
        RECT 1158.000000 119.910000 1168.000000 120.090000 ;
        RECT 1158.000000 115.910000 1168.000000 116.090000 ;
        RECT 1158.000000 111.910000 1168.000000 112.090000 ;
        RECT 1158.000000 123.910000 1168.000000 124.090000 ;
        RECT 1158.000000 127.910000 1168.000000 128.090000 ;
        RECT 1158.000000 135.910000 1168.000000 136.090000 ;
        RECT 1158.000000 131.910000 1168.000000 132.090000 ;
        RECT 1158.000000 139.910000 1168.000000 140.090000 ;
        RECT 1158.000000 143.910000 1168.000000 144.090000 ;
        RECT 1158.000000 147.910000 1168.000000 148.090000 ;
        RECT 1158.000000 155.910000 1168.000000 156.090000 ;
        RECT 1158.000000 151.910000 1168.000000 152.090000 ;
        RECT 1158.000000 159.910000 1168.000000 160.090000 ;
        RECT 1158.000000 163.910000 1168.000000 164.090000 ;
        RECT 1158.000000 175.910000 1168.000000 176.090000 ;
        RECT 1158.000000 171.910000 1168.000000 172.090000 ;
        RECT 1158.000000 167.910000 1168.000000 168.090000 ;
        RECT 1158.000000 179.910000 1168.000000 180.090000 ;
        RECT 1158.000000 183.910000 1168.000000 184.090000 ;
        RECT 1158.000000 191.910000 1168.000000 192.090000 ;
        RECT 1158.000000 187.910000 1168.000000 188.090000 ;
        RECT 960.000000 267.910000 965.000000 268.090000 ;
        RECT 960.000000 263.910000 965.000000 264.090000 ;
        RECT 960.000000 259.910000 965.000000 260.090000 ;
        RECT 910.000000 267.910000 915.000000 268.090000 ;
        RECT 910.000000 263.910000 915.000000 264.090000 ;
        RECT 910.000000 259.910000 915.000000 260.090000 ;
        RECT 1010.000000 259.910000 1015.000000 260.090000 ;
        RECT 1010.000000 263.910000 1015.000000 264.090000 ;
        RECT 1010.000000 267.910000 1015.000000 268.090000 ;
        RECT 960.000000 283.910000 965.000000 284.090000 ;
        RECT 960.000000 279.910000 965.000000 280.090000 ;
        RECT 960.000000 275.910000 965.000000 276.090000 ;
        RECT 960.000000 271.910000 965.000000 272.090000 ;
        RECT 960.000000 287.910000 965.000000 288.090000 ;
        RECT 960.000000 291.910000 965.000000 292.090000 ;
        RECT 960.000000 295.910000 965.000000 296.090000 ;
        RECT 960.000000 299.910000 965.000000 300.090000 ;
        RECT 960.000000 303.910000 965.000000 304.090000 ;
        RECT 960.000000 311.910000 965.000000 312.090000 ;
        RECT 960.000000 307.910000 965.000000 308.090000 ;
        RECT 960.000000 323.910000 965.000000 324.090000 ;
        RECT 960.000000 319.910000 965.000000 320.090000 ;
        RECT 960.000000 315.910000 965.000000 316.090000 ;
        RECT 960.000000 339.910000 965.000000 340.090000 ;
        RECT 960.000000 335.910000 965.000000 336.090000 ;
        RECT 960.000000 331.910000 965.000000 332.090000 ;
        RECT 960.000000 327.910000 965.000000 328.090000 ;
        RECT 910.000000 283.910000 915.000000 284.090000 ;
        RECT 910.000000 279.910000 915.000000 280.090000 ;
        RECT 910.000000 275.910000 915.000000 276.090000 ;
        RECT 910.000000 271.910000 915.000000 272.090000 ;
        RECT 910.000000 287.910000 915.000000 288.090000 ;
        RECT 910.000000 291.910000 915.000000 292.090000 ;
        RECT 910.000000 295.910000 915.000000 296.090000 ;
        RECT 910.000000 299.910000 915.000000 300.090000 ;
        RECT 910.000000 303.910000 915.000000 304.090000 ;
        RECT 910.000000 307.910000 915.000000 308.090000 ;
        RECT 910.000000 311.910000 915.000000 312.090000 ;
        RECT 910.000000 315.910000 915.000000 316.090000 ;
        RECT 910.000000 319.910000 915.000000 320.090000 ;
        RECT 910.000000 323.910000 915.000000 324.090000 ;
        RECT 910.000000 339.910000 915.000000 340.090000 ;
        RECT 910.000000 335.910000 915.000000 336.090000 ;
        RECT 910.000000 331.910000 915.000000 332.090000 ;
        RECT 910.000000 327.910000 915.000000 328.090000 ;
        RECT 1010.000000 271.910000 1015.000000 272.090000 ;
        RECT 1010.000000 275.910000 1015.000000 276.090000 ;
        RECT 1010.000000 283.910000 1015.000000 284.090000 ;
        RECT 1010.000000 279.910000 1015.000000 280.090000 ;
        RECT 1010.000000 287.910000 1015.000000 288.090000 ;
        RECT 1010.000000 291.910000 1015.000000 292.090000 ;
        RECT 1010.000000 295.910000 1015.000000 296.090000 ;
        RECT 1010.000000 303.910000 1015.000000 304.090000 ;
        RECT 1010.000000 299.910000 1015.000000 300.090000 ;
        RECT 1010.000000 311.910000 1015.000000 312.090000 ;
        RECT 1010.000000 307.910000 1015.000000 308.090000 ;
        RECT 1010.000000 315.910000 1015.000000 316.090000 ;
        RECT 1010.000000 319.910000 1015.000000 320.090000 ;
        RECT 1010.000000 323.910000 1015.000000 324.090000 ;
        RECT 1010.000000 331.910000 1015.000000 332.090000 ;
        RECT 1010.000000 327.910000 1015.000000 328.090000 ;
        RECT 1010.000000 335.910000 1015.000000 336.090000 ;
        RECT 1010.000000 339.910000 1015.000000 340.090000 ;
        RECT 1110.000000 267.910000 1115.000000 268.090000 ;
        RECT 1110.000000 263.910000 1115.000000 264.090000 ;
        RECT 1110.000000 259.910000 1115.000000 260.090000 ;
        RECT 1060.000000 267.910000 1065.000000 268.090000 ;
        RECT 1060.000000 263.910000 1065.000000 264.090000 ;
        RECT 1060.000000 259.910000 1065.000000 260.090000 ;
        RECT 1158.000000 203.910000 1168.000000 204.090000 ;
        RECT 1158.000000 195.910000 1168.000000 196.090000 ;
        RECT 1158.000000 199.910000 1168.000000 200.090000 ;
        RECT 1158.000000 211.910000 1168.000000 212.090000 ;
        RECT 1158.000000 207.910000 1168.000000 208.090000 ;
        RECT 1158.000000 215.910000 1168.000000 216.090000 ;
        RECT 1158.000000 219.910000 1168.000000 220.090000 ;
        RECT 1158.000000 227.910000 1168.000000 228.090000 ;
        RECT 1158.000000 223.910000 1168.000000 224.090000 ;
        RECT 1158.000000 231.910000 1168.000000 232.090000 ;
        RECT 1158.000000 235.910000 1168.000000 236.090000 ;
        RECT 1158.000000 239.910000 1168.000000 240.090000 ;
        RECT 1158.000000 247.910000 1168.000000 248.090000 ;
        RECT 1158.000000 243.910000 1168.000000 244.090000 ;
        RECT 1158.000000 251.910000 1168.000000 252.090000 ;
        RECT 1158.000000 255.910000 1168.000000 256.090000 ;
        RECT 1158.000000 267.910000 1168.000000 268.090000 ;
        RECT 1158.000000 259.910000 1168.000000 260.090000 ;
        RECT 1158.000000 263.910000 1168.000000 264.090000 ;
        RECT 1110.000000 283.910000 1115.000000 284.090000 ;
        RECT 1110.000000 279.910000 1115.000000 280.090000 ;
        RECT 1110.000000 275.910000 1115.000000 276.090000 ;
        RECT 1110.000000 271.910000 1115.000000 272.090000 ;
        RECT 1110.000000 287.910000 1115.000000 288.090000 ;
        RECT 1110.000000 291.910000 1115.000000 292.090000 ;
        RECT 1110.000000 295.910000 1115.000000 296.090000 ;
        RECT 1110.000000 299.910000 1115.000000 300.090000 ;
        RECT 1110.000000 303.910000 1115.000000 304.090000 ;
        RECT 1110.000000 311.910000 1115.000000 312.090000 ;
        RECT 1110.000000 307.910000 1115.000000 308.090000 ;
        RECT 1110.000000 323.910000 1115.000000 324.090000 ;
        RECT 1110.000000 319.910000 1115.000000 320.090000 ;
        RECT 1110.000000 315.910000 1115.000000 316.090000 ;
        RECT 1110.000000 339.910000 1115.000000 340.090000 ;
        RECT 1110.000000 335.910000 1115.000000 336.090000 ;
        RECT 1110.000000 331.910000 1115.000000 332.090000 ;
        RECT 1110.000000 327.910000 1115.000000 328.090000 ;
        RECT 1060.000000 283.910000 1065.000000 284.090000 ;
        RECT 1060.000000 279.910000 1065.000000 280.090000 ;
        RECT 1060.000000 275.910000 1065.000000 276.090000 ;
        RECT 1060.000000 271.910000 1065.000000 272.090000 ;
        RECT 1060.000000 287.910000 1065.000000 288.090000 ;
        RECT 1060.000000 291.910000 1065.000000 292.090000 ;
        RECT 1060.000000 295.910000 1065.000000 296.090000 ;
        RECT 1060.000000 299.910000 1065.000000 300.090000 ;
        RECT 1060.000000 303.910000 1065.000000 304.090000 ;
        RECT 1060.000000 307.910000 1065.000000 308.090000 ;
        RECT 1060.000000 311.910000 1065.000000 312.090000 ;
        RECT 1060.000000 315.910000 1065.000000 316.090000 ;
        RECT 1060.000000 319.910000 1065.000000 320.090000 ;
        RECT 1060.000000 323.910000 1065.000000 324.090000 ;
        RECT 1060.000000 339.910000 1065.000000 340.090000 ;
        RECT 1060.000000 335.910000 1065.000000 336.090000 ;
        RECT 1060.000000 331.910000 1065.000000 332.090000 ;
        RECT 1060.000000 327.910000 1065.000000 328.090000 ;
        RECT 1158.000000 283.910000 1168.000000 284.090000 ;
        RECT 1158.000000 279.910000 1168.000000 280.090000 ;
        RECT 1158.000000 275.910000 1168.000000 276.090000 ;
        RECT 1158.000000 271.910000 1168.000000 272.090000 ;
        RECT 1158.000000 287.910000 1168.000000 288.090000 ;
        RECT 1158.000000 291.910000 1168.000000 292.090000 ;
        RECT 1158.000000 295.910000 1168.000000 296.090000 ;
        RECT 1158.000000 299.910000 1168.000000 300.090000 ;
        RECT 1158.000000 303.910000 1168.000000 304.090000 ;
        RECT 1158.000000 307.910000 1168.000000 308.090000 ;
        RECT 1158.000000 311.910000 1168.000000 312.090000 ;
        RECT 1158.000000 315.910000 1168.000000 316.090000 ;
        RECT 1158.000000 319.910000 1168.000000 320.090000 ;
        RECT 1158.000000 323.910000 1168.000000 324.090000 ;
        RECT 1158.000000 339.910000 1168.000000 340.090000 ;
        RECT 1158.000000 335.910000 1168.000000 336.090000 ;
        RECT 1158.000000 331.910000 1168.000000 332.090000 ;
        RECT 1158.000000 327.910000 1168.000000 328.090000 ;
        RECT 60.000000 379.910000 65.000000 380.090000 ;
        RECT 18.000000 379.910000 28.000000 380.090000 ;
        RECT 18.000000 343.910000 28.000000 344.090000 ;
        RECT 18.000000 347.910000 28.000000 348.090000 ;
        RECT 18.000000 351.910000 28.000000 352.090000 ;
        RECT 18.000000 359.910000 28.000000 360.090000 ;
        RECT 18.000000 355.910000 28.000000 356.090000 ;
        RECT 18.000000 375.910000 28.000000 376.090000 ;
        RECT 18.000000 371.910000 28.000000 372.090000 ;
        RECT 18.000000 367.910000 28.000000 368.090000 ;
        RECT 18.000000 363.910000 28.000000 364.090000 ;
        RECT 60.000000 347.910000 65.000000 348.090000 ;
        RECT 60.000000 343.910000 65.000000 344.090000 ;
        RECT 60.000000 375.910000 65.000000 376.090000 ;
        RECT 60.000000 371.910000 65.000000 372.090000 ;
        RECT 60.000000 367.910000 65.000000 368.090000 ;
        RECT 60.000000 363.910000 65.000000 364.090000 ;
        RECT 18.000000 395.910000 28.000000 396.090000 ;
        RECT 18.000000 391.910000 28.000000 392.090000 ;
        RECT 18.000000 387.910000 28.000000 388.090000 ;
        RECT 18.000000 383.910000 28.000000 384.090000 ;
        RECT 18.000000 399.910000 28.000000 400.090000 ;
        RECT 18.000000 403.910000 28.000000 404.090000 ;
        RECT 18.000000 407.910000 28.000000 408.090000 ;
        RECT 18.000000 411.910000 28.000000 412.090000 ;
        RECT 18.000000 415.910000 28.000000 416.090000 ;
        RECT 60.000000 395.910000 65.000000 396.090000 ;
        RECT 60.000000 391.910000 65.000000 392.090000 ;
        RECT 60.000000 387.910000 65.000000 388.090000 ;
        RECT 60.000000 383.910000 65.000000 384.090000 ;
        RECT 60.000000 399.910000 65.000000 400.090000 ;
        RECT 60.000000 403.910000 65.000000 404.090000 ;
        RECT 60.000000 407.910000 65.000000 408.090000 ;
        RECT 60.000000 411.910000 65.000000 412.090000 ;
        RECT 60.000000 415.910000 65.000000 416.090000 ;
        RECT 110.000000 379.910000 115.000000 380.090000 ;
        RECT 110.000000 351.910000 115.000000 352.090000 ;
        RECT 110.000000 347.910000 115.000000 348.090000 ;
        RECT 110.000000 343.910000 115.000000 344.090000 ;
        RECT 110.000000 359.910000 115.000000 360.090000 ;
        RECT 110.000000 355.910000 115.000000 356.090000 ;
        RECT 110.000000 375.910000 115.000000 376.090000 ;
        RECT 110.000000 371.910000 115.000000 372.090000 ;
        RECT 110.000000 367.910000 115.000000 368.090000 ;
        RECT 110.000000 363.910000 115.000000 364.090000 ;
        RECT 110.000000 383.910000 115.000000 384.090000 ;
        RECT 110.000000 387.910000 115.000000 388.090000 ;
        RECT 110.000000 391.910000 115.000000 392.090000 ;
        RECT 110.000000 395.910000 115.000000 396.090000 ;
        RECT 110.000000 399.910000 115.000000 400.090000 ;
        RECT 110.000000 403.910000 115.000000 404.090000 ;
        RECT 110.000000 407.910000 115.000000 408.090000 ;
        RECT 110.000000 411.910000 115.000000 412.090000 ;
        RECT 110.000000 415.910000 115.000000 416.090000 ;
        RECT 18.000000 431.910000 28.000000 432.090000 ;
        RECT 18.000000 427.910000 28.000000 428.090000 ;
        RECT 18.000000 423.910000 28.000000 424.090000 ;
        RECT 18.000000 419.910000 28.000000 420.090000 ;
        RECT 18.000000 435.910000 28.000000 436.090000 ;
        RECT 18.000000 439.910000 28.000000 440.090000 ;
        RECT 18.000000 443.910000 28.000000 444.090000 ;
        RECT 18.000000 447.910000 28.000000 448.090000 ;
        RECT 18.000000 451.910000 28.000000 452.090000 ;
        RECT 60.000000 431.910000 65.000000 432.090000 ;
        RECT 60.000000 427.910000 65.000000 428.090000 ;
        RECT 60.000000 423.910000 65.000000 424.090000 ;
        RECT 60.000000 419.910000 65.000000 420.090000 ;
        RECT 60.000000 435.910000 65.000000 436.090000 ;
        RECT 60.000000 439.910000 65.000000 440.090000 ;
        RECT 60.000000 443.910000 65.000000 444.090000 ;
        RECT 60.000000 447.910000 65.000000 448.090000 ;
        RECT 60.000000 451.910000 65.000000 452.090000 ;
        RECT 18.000000 455.910000 28.000000 456.090000 ;
        RECT 18.000000 459.910000 28.000000 460.090000 ;
        RECT 18.000000 463.910000 28.000000 464.090000 ;
        RECT 18.000000 467.910000 28.000000 468.090000 ;
        RECT 18.000000 471.910000 28.000000 472.090000 ;
        RECT 18.000000 487.910000 28.000000 488.090000 ;
        RECT 18.000000 483.910000 28.000000 484.090000 ;
        RECT 18.000000 479.910000 28.000000 480.090000 ;
        RECT 18.000000 475.910000 28.000000 476.090000 ;
        RECT 60.000000 455.910000 65.000000 456.090000 ;
        RECT 60.000000 459.910000 65.000000 460.090000 ;
        RECT 60.000000 463.910000 65.000000 464.090000 ;
        RECT 60.000000 467.910000 65.000000 468.090000 ;
        RECT 60.000000 471.910000 65.000000 472.090000 ;
        RECT 60.000000 487.910000 65.000000 488.090000 ;
        RECT 60.000000 483.910000 65.000000 484.090000 ;
        RECT 60.000000 479.910000 65.000000 480.090000 ;
        RECT 60.000000 475.910000 65.000000 476.090000 ;
        RECT 110.000000 419.910000 115.000000 420.090000 ;
        RECT 110.000000 423.910000 115.000000 424.090000 ;
        RECT 110.000000 427.910000 115.000000 428.090000 ;
        RECT 110.000000 431.910000 115.000000 432.090000 ;
        RECT 110.000000 435.910000 115.000000 436.090000 ;
        RECT 110.000000 439.910000 115.000000 440.090000 ;
        RECT 110.000000 443.910000 115.000000 444.090000 ;
        RECT 110.000000 447.910000 115.000000 448.090000 ;
        RECT 110.000000 451.910000 115.000000 452.090000 ;
        RECT 110.000000 459.910000 115.000000 460.090000 ;
        RECT 110.000000 455.910000 115.000000 456.090000 ;
        RECT 110.000000 471.910000 115.000000 472.090000 ;
        RECT 110.000000 467.910000 115.000000 468.090000 ;
        RECT 110.000000 463.910000 115.000000 464.090000 ;
        RECT 110.000000 487.910000 115.000000 488.090000 ;
        RECT 110.000000 483.910000 115.000000 484.090000 ;
        RECT 110.000000 479.910000 115.000000 480.090000 ;
        RECT 110.000000 475.910000 115.000000 476.090000 ;
        RECT 210.000000 379.910000 215.000000 380.090000 ;
        RECT 160.000000 379.910000 165.000000 380.090000 ;
        RECT 160.000000 343.910000 165.000000 344.090000 ;
        RECT 160.000000 347.910000 165.000000 348.090000 ;
        RECT 160.000000 351.910000 165.000000 352.090000 ;
        RECT 160.000000 359.910000 165.000000 360.090000 ;
        RECT 160.000000 355.910000 165.000000 356.090000 ;
        RECT 160.000000 363.910000 165.000000 364.090000 ;
        RECT 160.000000 367.910000 165.000000 368.090000 ;
        RECT 160.000000 371.910000 165.000000 372.090000 ;
        RECT 160.000000 375.910000 165.000000 376.090000 ;
        RECT 210.000000 343.910000 215.000000 344.090000 ;
        RECT 210.000000 347.910000 215.000000 348.090000 ;
        RECT 210.000000 351.910000 215.000000 352.090000 ;
        RECT 210.000000 355.910000 215.000000 356.090000 ;
        RECT 210.000000 359.910000 215.000000 360.090000 ;
        RECT 210.000000 375.910000 215.000000 376.090000 ;
        RECT 210.000000 371.910000 215.000000 372.090000 ;
        RECT 210.000000 367.910000 215.000000 368.090000 ;
        RECT 210.000000 363.910000 215.000000 364.090000 ;
        RECT 160.000000 383.910000 165.000000 384.090000 ;
        RECT 160.000000 387.910000 165.000000 388.090000 ;
        RECT 160.000000 391.910000 165.000000 392.090000 ;
        RECT 160.000000 395.910000 165.000000 396.090000 ;
        RECT 160.000000 403.910000 165.000000 404.090000 ;
        RECT 160.000000 399.910000 165.000000 400.090000 ;
        RECT 160.000000 407.910000 165.000000 408.090000 ;
        RECT 210.000000 383.910000 215.000000 384.090000 ;
        RECT 210.000000 387.910000 215.000000 388.090000 ;
        RECT 210.000000 391.910000 215.000000 392.090000 ;
        RECT 210.000000 395.910000 215.000000 396.090000 ;
        RECT 210.000000 399.910000 215.000000 400.090000 ;
        RECT 210.000000 403.910000 215.000000 404.090000 ;
        RECT 210.000000 407.910000 215.000000 408.090000 ;
        RECT 210.000000 411.910000 215.000000 412.090000 ;
        RECT 210.000000 415.910000 215.000000 416.090000 ;
        RECT 260.000000 379.910000 265.000000 380.090000 ;
        RECT 260.000000 351.910000 265.000000 352.090000 ;
        RECT 260.000000 347.910000 265.000000 348.090000 ;
        RECT 260.000000 343.910000 265.000000 344.090000 ;
        RECT 260.000000 359.910000 265.000000 360.090000 ;
        RECT 260.000000 355.910000 265.000000 356.090000 ;
        RECT 260.000000 367.910000 265.000000 368.090000 ;
        RECT 260.000000 363.910000 265.000000 364.090000 ;
        RECT 260.000000 375.910000 265.000000 376.090000 ;
        RECT 260.000000 371.910000 265.000000 372.090000 ;
        RECT 260.000000 383.910000 265.000000 384.090000 ;
        RECT 260.000000 387.910000 265.000000 388.090000 ;
        RECT 260.000000 391.910000 265.000000 392.090000 ;
        RECT 260.000000 395.910000 265.000000 396.090000 ;
        RECT 260.000000 399.910000 265.000000 400.090000 ;
        RECT 260.000000 403.910000 265.000000 404.090000 ;
        RECT 260.000000 407.910000 265.000000 408.090000 ;
        RECT 210.000000 431.910000 215.000000 432.090000 ;
        RECT 210.000000 427.910000 215.000000 428.090000 ;
        RECT 210.000000 423.910000 215.000000 424.090000 ;
        RECT 210.000000 419.910000 215.000000 420.090000 ;
        RECT 210.000000 435.910000 215.000000 436.090000 ;
        RECT 210.000000 439.910000 215.000000 440.090000 ;
        RECT 210.000000 443.910000 215.000000 444.090000 ;
        RECT 210.000000 447.910000 215.000000 448.090000 ;
        RECT 210.000000 451.910000 215.000000 452.090000 ;
        RECT 160.000000 463.910000 165.000000 464.090000 ;
        RECT 160.000000 467.910000 165.000000 468.090000 ;
        RECT 160.000000 471.910000 165.000000 472.090000 ;
        RECT 160.000000 479.910000 165.000000 480.090000 ;
        RECT 160.000000 475.910000 165.000000 476.090000 ;
        RECT 160.000000 487.910000 165.000000 488.090000 ;
        RECT 160.000000 483.910000 165.000000 484.090000 ;
        RECT 210.000000 455.910000 215.000000 456.090000 ;
        RECT 210.000000 459.910000 215.000000 460.090000 ;
        RECT 210.000000 467.910000 215.000000 468.090000 ;
        RECT 210.000000 463.910000 215.000000 464.090000 ;
        RECT 210.000000 471.910000 215.000000 472.090000 ;
        RECT 210.000000 487.910000 215.000000 488.090000 ;
        RECT 210.000000 483.910000 215.000000 484.090000 ;
        RECT 210.000000 479.910000 215.000000 480.090000 ;
        RECT 210.000000 475.910000 215.000000 476.090000 ;
        RECT 260.000000 471.910000 265.000000 472.090000 ;
        RECT 260.000000 467.910000 265.000000 468.090000 ;
        RECT 260.000000 463.910000 265.000000 464.090000 ;
        RECT 260.000000 479.910000 265.000000 480.090000 ;
        RECT 260.000000 475.910000 265.000000 476.090000 ;
        RECT 260.000000 483.910000 265.000000 484.090000 ;
        RECT 260.000000 487.910000 265.000000 488.090000 ;
        RECT 18.000000 491.910000 28.000000 492.090000 ;
        RECT 18.000000 495.910000 28.000000 496.090000 ;
        RECT 18.000000 499.910000 28.000000 500.090000 ;
        RECT 18.000000 503.910000 28.000000 504.090000 ;
        RECT 18.000000 507.910000 28.000000 508.090000 ;
        RECT 18.000000 515.910000 28.000000 516.090000 ;
        RECT 18.000000 511.910000 28.000000 512.090000 ;
        RECT 60.000000 491.910000 65.000000 492.090000 ;
        RECT 60.000000 495.910000 65.000000 496.090000 ;
        RECT 60.000000 499.910000 65.000000 500.090000 ;
        RECT 60.000000 503.910000 65.000000 504.090000 ;
        RECT 60.000000 507.910000 65.000000 508.090000 ;
        RECT 60.000000 515.910000 65.000000 516.090000 ;
        RECT 60.000000 511.910000 65.000000 512.090000 ;
        RECT 110.000000 499.910000 115.000000 500.090000 ;
        RECT 110.000000 495.910000 115.000000 496.090000 ;
        RECT 110.000000 491.910000 115.000000 492.090000 ;
        RECT 110.000000 507.910000 115.000000 508.090000 ;
        RECT 110.000000 503.910000 115.000000 504.090000 ;
        RECT 110.000000 515.910000 115.000000 516.090000 ;
        RECT 110.000000 511.910000 115.000000 512.090000 ;
        RECT 160.000000 491.910000 165.000000 492.090000 ;
        RECT 160.000000 495.910000 165.000000 496.090000 ;
        RECT 160.000000 499.910000 165.000000 500.090000 ;
        RECT 160.000000 507.910000 165.000000 508.090000 ;
        RECT 160.000000 503.910000 165.000000 504.090000 ;
        RECT 160.000000 511.910000 165.000000 512.090000 ;
        RECT 160.000000 515.910000 165.000000 516.090000 ;
        RECT 210.000000 491.910000 215.000000 492.090000 ;
        RECT 210.000000 495.910000 215.000000 496.090000 ;
        RECT 210.000000 499.910000 215.000000 500.090000 ;
        RECT 210.000000 503.910000 215.000000 504.090000 ;
        RECT 210.000000 507.910000 215.000000 508.090000 ;
        RECT 210.000000 515.910000 215.000000 516.090000 ;
        RECT 210.000000 511.910000 215.000000 512.090000 ;
        RECT 260.000000 491.910000 265.000000 492.090000 ;
        RECT 260.000000 495.910000 265.000000 496.090000 ;
        RECT 260.000000 499.910000 265.000000 500.090000 ;
        RECT 260.000000 503.910000 265.000000 504.090000 ;
        RECT 260.000000 507.910000 265.000000 508.090000 ;
        RECT 260.000000 511.910000 265.000000 512.090000 ;
        RECT 260.000000 515.910000 265.000000 516.090000 ;
        RECT 310.000000 379.910000 315.000000 380.090000 ;
        RECT 360.000000 379.910000 365.000000 380.090000 ;
        RECT 310.000000 343.910000 315.000000 344.090000 ;
        RECT 310.000000 351.910000 315.000000 352.090000 ;
        RECT 310.000000 347.910000 315.000000 348.090000 ;
        RECT 310.000000 355.910000 315.000000 356.090000 ;
        RECT 310.000000 359.910000 315.000000 360.090000 ;
        RECT 310.000000 363.910000 315.000000 364.090000 ;
        RECT 310.000000 367.910000 315.000000 368.090000 ;
        RECT 310.000000 371.910000 315.000000 372.090000 ;
        RECT 310.000000 375.910000 315.000000 376.090000 ;
        RECT 360.000000 343.910000 365.000000 344.090000 ;
        RECT 360.000000 347.910000 365.000000 348.090000 ;
        RECT 360.000000 351.910000 365.000000 352.090000 ;
        RECT 360.000000 355.910000 365.000000 356.090000 ;
        RECT 360.000000 359.910000 365.000000 360.090000 ;
        RECT 360.000000 363.910000 365.000000 364.090000 ;
        RECT 360.000000 367.910000 365.000000 368.090000 ;
        RECT 360.000000 371.910000 365.000000 372.090000 ;
        RECT 360.000000 375.910000 365.000000 376.090000 ;
        RECT 310.000000 383.910000 315.000000 384.090000 ;
        RECT 310.000000 387.910000 315.000000 388.090000 ;
        RECT 310.000000 391.910000 315.000000 392.090000 ;
        RECT 310.000000 395.910000 315.000000 396.090000 ;
        RECT 310.000000 399.910000 315.000000 400.090000 ;
        RECT 310.000000 403.910000 315.000000 404.090000 ;
        RECT 310.000000 411.910000 315.000000 412.090000 ;
        RECT 310.000000 407.910000 315.000000 408.090000 ;
        RECT 310.000000 415.910000 315.000000 416.090000 ;
        RECT 360.000000 383.910000 365.000000 384.090000 ;
        RECT 360.000000 387.910000 365.000000 388.090000 ;
        RECT 360.000000 391.910000 365.000000 392.090000 ;
        RECT 360.000000 395.910000 365.000000 396.090000 ;
        RECT 360.000000 399.910000 365.000000 400.090000 ;
        RECT 360.000000 403.910000 365.000000 404.090000 ;
        RECT 360.000000 407.910000 365.000000 408.090000 ;
        RECT 360.000000 411.910000 365.000000 412.090000 ;
        RECT 360.000000 415.910000 365.000000 416.090000 ;
        RECT 410.000000 379.910000 415.000000 380.090000 ;
        RECT 410.000000 343.910000 415.000000 344.090000 ;
        RECT 410.000000 347.910000 415.000000 348.090000 ;
        RECT 410.000000 351.910000 415.000000 352.090000 ;
        RECT 410.000000 355.910000 415.000000 356.090000 ;
        RECT 410.000000 359.910000 415.000000 360.090000 ;
        RECT 410.000000 363.910000 415.000000 364.090000 ;
        RECT 410.000000 367.910000 415.000000 368.090000 ;
        RECT 410.000000 371.910000 415.000000 372.090000 ;
        RECT 410.000000 375.910000 415.000000 376.090000 ;
        RECT 410.000000 383.910000 415.000000 384.090000 ;
        RECT 410.000000 387.910000 415.000000 388.090000 ;
        RECT 410.000000 391.910000 415.000000 392.090000 ;
        RECT 410.000000 395.910000 415.000000 396.090000 ;
        RECT 410.000000 399.910000 415.000000 400.090000 ;
        RECT 410.000000 403.910000 415.000000 404.090000 ;
        RECT 410.000000 411.910000 415.000000 412.090000 ;
        RECT 410.000000 407.910000 415.000000 408.090000 ;
        RECT 410.000000 415.910000 415.000000 416.090000 ;
        RECT 361.000000 479.910000 371.000000 480.090000 ;
        RECT 361.000000 483.910000 371.000000 484.090000 ;
        RECT 361.000000 487.910000 371.000000 488.090000 ;
        RECT 310.000000 419.910000 315.000000 420.090000 ;
        RECT 310.000000 423.910000 315.000000 424.090000 ;
        RECT 310.000000 427.910000 315.000000 428.090000 ;
        RECT 310.000000 431.910000 315.000000 432.090000 ;
        RECT 310.000000 439.910000 315.000000 440.090000 ;
        RECT 310.000000 435.910000 315.000000 436.090000 ;
        RECT 310.000000 443.910000 315.000000 444.090000 ;
        RECT 310.000000 447.910000 315.000000 448.090000 ;
        RECT 310.000000 451.910000 315.000000 452.090000 ;
        RECT 360.000000 419.910000 365.000000 420.090000 ;
        RECT 360.000000 423.910000 365.000000 424.090000 ;
        RECT 360.000000 427.910000 365.000000 428.090000 ;
        RECT 360.000000 431.910000 365.000000 432.090000 ;
        RECT 360.000000 435.910000 365.000000 436.090000 ;
        RECT 360.000000 439.910000 365.000000 440.090000 ;
        RECT 360.000000 443.910000 365.000000 444.090000 ;
        RECT 360.000000 447.910000 365.000000 448.090000 ;
        RECT 360.000000 451.910000 365.000000 452.090000 ;
        RECT 310.000000 455.910000 315.000000 456.090000 ;
        RECT 310.000000 459.910000 315.000000 460.090000 ;
        RECT 310.000000 467.910000 315.000000 468.090000 ;
        RECT 310.000000 463.910000 315.000000 464.090000 ;
        RECT 310.000000 471.910000 315.000000 472.090000 ;
        RECT 310.000000 475.910000 315.000000 476.090000 ;
        RECT 310.000000 479.910000 315.000000 480.090000 ;
        RECT 310.000000 487.910000 315.000000 488.090000 ;
        RECT 310.000000 483.910000 315.000000 484.090000 ;
        RECT 360.000000 455.910000 365.000000 456.090000 ;
        RECT 360.000000 459.910000 365.000000 460.090000 ;
        RECT 360.000000 471.910000 368.500000 472.090000 ;
        RECT 360.000000 463.910000 365.000000 464.090000 ;
        RECT 360.000000 467.910000 365.000000 468.090000 ;
        RECT 363.500000 475.910000 368.500000 476.090000 ;
        RECT 410.000000 419.910000 415.000000 420.090000 ;
        RECT 410.000000 423.910000 415.000000 424.090000 ;
        RECT 410.000000 427.910000 415.000000 428.090000 ;
        RECT 410.000000 431.910000 415.000000 432.090000 ;
        RECT 410.000000 439.910000 415.000000 440.090000 ;
        RECT 410.000000 435.910000 415.000000 436.090000 ;
        RECT 410.000000 443.910000 415.000000 444.090000 ;
        RECT 410.000000 451.910000 415.000000 452.090000 ;
        RECT 410.000000 447.910000 415.000000 448.090000 ;
        RECT 410.000000 455.910000 415.000000 456.090000 ;
        RECT 410.000000 459.910000 415.000000 460.090000 ;
        RECT 410.000000 467.910000 415.000000 468.090000 ;
        RECT 410.000000 463.910000 415.000000 464.090000 ;
        RECT 410.000000 471.910000 415.000000 472.090000 ;
        RECT 410.000000 475.910000 415.000000 476.090000 ;
        RECT 410.000000 479.910000 415.000000 480.090000 ;
        RECT 410.000000 483.910000 415.000000 484.090000 ;
        RECT 410.000000 487.910000 415.000000 488.090000 ;
        RECT 460.000000 379.910000 465.000000 380.090000 ;
        RECT 510.000000 379.910000 515.000000 380.090000 ;
        RECT 460.000000 347.910000 465.000000 348.090000 ;
        RECT 460.000000 343.910000 465.000000 344.090000 ;
        RECT 460.000000 375.910000 465.000000 376.090000 ;
        RECT 460.000000 371.910000 465.000000 372.090000 ;
        RECT 510.000000 343.910000 515.000000 344.090000 ;
        RECT 510.000000 351.910000 515.000000 352.090000 ;
        RECT 510.000000 347.910000 515.000000 348.090000 ;
        RECT 510.000000 359.910000 515.000000 360.090000 ;
        RECT 510.000000 355.910000 515.000000 356.090000 ;
        RECT 510.000000 363.910000 515.000000 364.090000 ;
        RECT 510.000000 367.910000 515.000000 368.090000 ;
        RECT 510.000000 375.910000 515.000000 376.090000 ;
        RECT 510.000000 371.910000 515.000000 372.090000 ;
        RECT 460.000000 383.910000 465.000000 384.090000 ;
        RECT 460.000000 387.910000 465.000000 388.090000 ;
        RECT 460.000000 391.910000 465.000000 392.090000 ;
        RECT 460.000000 395.910000 465.000000 396.090000 ;
        RECT 510.000000 383.910000 515.000000 384.090000 ;
        RECT 510.000000 387.910000 515.000000 388.090000 ;
        RECT 510.000000 391.910000 515.000000 392.090000 ;
        RECT 510.000000 395.910000 515.000000 396.090000 ;
        RECT 510.000000 399.910000 515.000000 400.090000 ;
        RECT 510.000000 403.910000 515.000000 404.090000 ;
        RECT 510.000000 407.910000 515.000000 408.090000 ;
        RECT 510.000000 411.910000 515.000000 412.090000 ;
        RECT 510.000000 415.910000 515.000000 416.090000 ;
        RECT 560.000000 379.910000 565.000000 380.090000 ;
        RECT 560.000000 343.910000 565.000000 344.090000 ;
        RECT 560.000000 347.910000 565.000000 348.090000 ;
        RECT 560.000000 351.910000 565.000000 352.090000 ;
        RECT 560.000000 355.910000 565.000000 356.090000 ;
        RECT 560.000000 359.910000 565.000000 360.090000 ;
        RECT 560.000000 363.910000 565.000000 364.090000 ;
        RECT 560.000000 367.910000 565.000000 368.090000 ;
        RECT 560.000000 371.910000 565.000000 372.090000 ;
        RECT 560.000000 375.910000 565.000000 376.090000 ;
        RECT 560.000000 383.910000 565.000000 384.090000 ;
        RECT 560.000000 387.910000 565.000000 388.090000 ;
        RECT 560.000000 391.910000 565.000000 392.090000 ;
        RECT 560.000000 395.910000 565.000000 396.090000 ;
        RECT 560.000000 403.910000 565.000000 404.090000 ;
        RECT 560.000000 399.910000 565.000000 400.090000 ;
        RECT 560.000000 411.910000 565.000000 412.090000 ;
        RECT 560.000000 407.910000 565.000000 408.090000 ;
        RECT 560.000000 415.910000 565.000000 416.090000 ;
        RECT 460.000000 423.910000 465.000000 424.090000 ;
        RECT 460.000000 419.910000 465.000000 420.090000 ;
        RECT 460.000000 427.910000 465.000000 428.090000 ;
        RECT 460.000000 431.910000 465.000000 432.090000 ;
        RECT 460.000000 435.910000 465.000000 436.090000 ;
        RECT 460.000000 439.910000 465.000000 440.090000 ;
        RECT 460.000000 443.910000 465.000000 444.090000 ;
        RECT 460.000000 447.910000 465.000000 448.090000 ;
        RECT 460.000000 451.910000 465.000000 452.090000 ;
        RECT 510.000000 419.910000 515.000000 420.090000 ;
        RECT 510.000000 423.910000 515.000000 424.090000 ;
        RECT 510.000000 431.910000 515.000000 432.090000 ;
        RECT 510.000000 427.910000 515.000000 428.090000 ;
        RECT 510.000000 435.910000 515.000000 436.090000 ;
        RECT 510.000000 439.910000 515.000000 440.090000 ;
        RECT 510.000000 443.910000 515.000000 444.090000 ;
        RECT 510.000000 447.910000 515.000000 448.090000 ;
        RECT 510.000000 451.910000 515.000000 452.090000 ;
        RECT 460.000000 455.910000 465.000000 456.090000 ;
        RECT 460.000000 459.910000 465.000000 460.090000 ;
        RECT 460.000000 463.910000 465.000000 464.090000 ;
        RECT 460.000000 467.910000 465.000000 468.090000 ;
        RECT 460.000000 471.910000 465.000000 472.090000 ;
        RECT 460.000000 475.910000 465.000000 476.090000 ;
        RECT 460.000000 479.910000 465.000000 480.090000 ;
        RECT 460.000000 483.910000 465.000000 484.090000 ;
        RECT 460.000000 487.910000 465.000000 488.090000 ;
        RECT 510.000000 459.910000 515.000000 460.090000 ;
        RECT 510.000000 455.910000 515.000000 456.090000 ;
        RECT 510.000000 463.910000 515.000000 464.090000 ;
        RECT 510.000000 467.910000 515.000000 468.090000 ;
        RECT 510.000000 471.910000 515.000000 472.090000 ;
        RECT 510.000000 479.910000 515.000000 480.090000 ;
        RECT 510.000000 475.910000 515.000000 476.090000 ;
        RECT 510.000000 487.910000 515.000000 488.090000 ;
        RECT 510.000000 483.910000 515.000000 484.090000 ;
        RECT 560.000000 419.910000 565.000000 420.090000 ;
        RECT 560.000000 423.910000 565.000000 424.090000 ;
        RECT 560.000000 427.910000 565.000000 428.090000 ;
        RECT 560.000000 431.910000 565.000000 432.090000 ;
        RECT 560.000000 443.910000 565.000000 444.090000 ;
        RECT 560.000000 439.910000 565.000000 440.090000 ;
        RECT 560.000000 435.910000 565.000000 436.090000 ;
        RECT 560.000000 451.910000 565.000000 452.090000 ;
        RECT 560.000000 447.910000 565.000000 448.090000 ;
        RECT 560.000000 455.910000 565.000000 456.090000 ;
        RECT 560.000000 459.910000 565.000000 460.090000 ;
        RECT 560.000000 471.910000 565.000000 472.090000 ;
        RECT 560.000000 463.910000 565.000000 464.090000 ;
        RECT 560.000000 467.910000 565.000000 468.090000 ;
        RECT 560.000000 475.910000 565.000000 476.090000 ;
        RECT 560.000000 479.910000 565.000000 480.090000 ;
        RECT 560.000000 483.910000 565.000000 484.090000 ;
        RECT 560.000000 487.910000 565.000000 488.090000 ;
        RECT 360.000000 499.910000 371.000000 500.090000 ;
        RECT 360.000000 491.910000 371.000000 492.090000 ;
        RECT 360.000000 495.910000 371.000000 496.090000 ;
        RECT 360.000000 507.910000 371.000000 508.090000 ;
        RECT 360.000000 503.910000 371.000000 504.090000 ;
        RECT 360.000000 511.910000 371.000000 512.090000 ;
        RECT 360.000000 515.910000 371.000000 516.090000 ;
        RECT 360.000000 519.910000 371.000000 520.090000 ;
        RECT 360.000000 523.910000 371.000000 524.090000 ;
        RECT 360.000000 527.910000 371.000000 528.090000 ;
        RECT 360.000000 535.910000 371.000000 536.090000 ;
        RECT 360.000000 531.910000 371.000000 532.090000 ;
        RECT 360.000000 543.910000 371.000000 544.090000 ;
        RECT 360.000000 539.910000 371.000000 540.090000 ;
        RECT 360.000000 547.910000 371.000000 548.090000 ;
        RECT 360.000000 551.910000 371.000000 552.090000 ;
        RECT 360.000000 555.910000 371.000000 556.090000 ;
        RECT 360.000000 563.910000 371.000000 564.090000 ;
        RECT 360.000000 559.910000 371.000000 560.090000 ;
        RECT 310.000000 491.910000 315.000000 492.090000 ;
        RECT 310.000000 495.910000 315.000000 496.090000 ;
        RECT 310.000000 499.910000 315.000000 500.090000 ;
        RECT 310.000000 507.910000 315.000000 508.090000 ;
        RECT 310.000000 503.910000 315.000000 504.090000 ;
        RECT 310.000000 511.910000 315.000000 512.090000 ;
        RECT 310.000000 515.910000 315.000000 516.090000 ;
        RECT 410.000000 491.910000 415.000000 492.090000 ;
        RECT 410.000000 495.910000 415.000000 496.090000 ;
        RECT 410.000000 499.910000 415.000000 500.090000 ;
        RECT 410.000000 503.910000 415.000000 504.090000 ;
        RECT 360.000000 571.910000 371.000000 572.090000 ;
        RECT 360.000000 567.910000 371.000000 568.090000 ;
        RECT 360.000000 579.910000 371.000000 580.090000 ;
        RECT 360.000000 575.910000 371.000000 576.090000 ;
        RECT 360.000000 583.910000 371.000000 584.090000 ;
        RECT 360.000000 587.910000 371.000000 588.090000 ;
        RECT 360.000000 591.910000 371.000000 592.090000 ;
        RECT 360.000000 599.910000 371.000000 600.090000 ;
        RECT 360.000000 595.910000 371.000000 596.090000 ;
        RECT 360.000000 607.910000 371.000000 608.090000 ;
        RECT 360.000000 603.910000 371.000000 604.090000 ;
        RECT 360.000000 619.910000 371.000000 620.090000 ;
        RECT 360.000000 615.910000 371.000000 616.090000 ;
        RECT 360.000000 611.910000 371.000000 612.090000 ;
        RECT 360.000000 623.910000 371.000000 624.090000 ;
        RECT 360.000000 627.910000 371.000000 628.090000 ;
        RECT 360.000000 635.910000 371.000000 636.090000 ;
        RECT 360.000000 631.910000 371.000000 632.090000 ;
        RECT 460.000000 503.910000 465.000000 504.090000 ;
        RECT 460.000000 499.910000 465.000000 500.090000 ;
        RECT 460.000000 491.910000 465.000000 492.090000 ;
        RECT 460.000000 495.910000 465.000000 496.090000 ;
        RECT 510.000000 495.910000 515.000000 496.090000 ;
        RECT 510.000000 491.910000 515.000000 492.090000 ;
        RECT 510.000000 499.910000 515.000000 500.090000 ;
        RECT 510.000000 503.910000 515.000000 504.090000 ;
        RECT 560.000000 499.910000 565.000000 500.090000 ;
        RECT 560.000000 495.910000 565.000000 496.090000 ;
        RECT 560.000000 491.910000 565.000000 492.090000 ;
        RECT 560.000000 503.910000 565.000000 504.090000 ;
        RECT 360.000000 647.910000 371.000000 648.090000 ;
        RECT 360.000000 639.910000 371.000000 640.090000 ;
        RECT 360.000000 643.910000 371.000000 644.090000 ;
        RECT 360.000000 655.910000 371.000000 656.090000 ;
        RECT 360.000000 651.910000 371.000000 652.090000 ;
        RECT 360.000000 667.910000 371.000000 668.090000 ;
        RECT 360.000000 663.910000 371.000000 664.090000 ;
        RECT 360.000000 659.910000 371.000000 660.090000 ;
        RECT 360.000000 675.910000 365.000000 676.090000 ;
        RECT 360.000000 671.910000 365.000000 672.090000 ;
        RECT 310.000000 679.910000 315.000000 680.090000 ;
        RECT 310.000000 683.910000 315.000000 684.090000 ;
        RECT 360.000000 679.910000 365.000000 680.090000 ;
        RECT 360.000000 683.910000 365.000000 684.090000 ;
        RECT 410.000000 659.910000 415.000000 660.090000 ;
        RECT 410.000000 663.910000 415.000000 664.090000 ;
        RECT 410.000000 667.910000 415.000000 668.090000 ;
        RECT 410.000000 671.910000 415.000000 672.090000 ;
        RECT 410.000000 675.910000 415.000000 676.090000 ;
        RECT 410.000000 683.910000 415.000000 684.090000 ;
        RECT 410.000000 679.910000 415.000000 680.090000 ;
        RECT 460.000000 659.910000 465.000000 660.090000 ;
        RECT 460.000000 663.910000 465.000000 664.090000 ;
        RECT 460.000000 667.910000 465.000000 668.090000 ;
        RECT 460.000000 671.910000 465.000000 672.090000 ;
        RECT 460.000000 675.910000 465.000000 676.090000 ;
        RECT 510.000000 663.910000 515.000000 664.090000 ;
        RECT 510.000000 659.910000 515.000000 660.090000 ;
        RECT 510.000000 667.910000 515.000000 668.090000 ;
        RECT 510.000000 671.910000 515.000000 672.090000 ;
        RECT 510.000000 675.910000 515.000000 676.090000 ;
        RECT 460.000000 683.910000 465.000000 684.090000 ;
        RECT 460.000000 679.910000 465.000000 680.090000 ;
        RECT 510.000000 683.910000 515.000000 684.090000 ;
        RECT 510.000000 679.910000 515.000000 680.090000 ;
        RECT 560.000000 659.910000 565.000000 660.090000 ;
        RECT 560.000000 663.910000 565.000000 664.090000 ;
        RECT 560.000000 667.910000 565.000000 668.090000 ;
        RECT 560.000000 671.910000 565.000000 672.090000 ;
        RECT 560.000000 675.910000 565.000000 676.090000 ;
        RECT 560.000000 683.910000 565.000000 684.090000 ;
        RECT 560.000000 679.910000 565.000000 680.090000 ;
        RECT 610.000000 379.910000 615.000000 380.090000 ;
        RECT 660.000000 379.910000 665.000000 380.090000 ;
        RECT 610.000000 343.910000 615.000000 344.090000 ;
        RECT 610.000000 347.910000 615.000000 348.090000 ;
        RECT 610.000000 351.910000 615.000000 352.090000 ;
        RECT 610.000000 355.910000 615.000000 356.090000 ;
        RECT 610.000000 359.910000 615.000000 360.090000 ;
        RECT 610.000000 363.910000 615.000000 364.090000 ;
        RECT 610.000000 367.910000 615.000000 368.090000 ;
        RECT 610.000000 371.910000 615.000000 372.090000 ;
        RECT 610.000000 375.910000 615.000000 376.090000 ;
        RECT 660.000000 343.910000 665.000000 344.090000 ;
        RECT 660.000000 351.910000 665.000000 352.090000 ;
        RECT 660.000000 347.910000 665.000000 348.090000 ;
        RECT 660.000000 355.910000 665.000000 356.090000 ;
        RECT 660.000000 359.910000 665.000000 360.090000 ;
        RECT 660.000000 363.910000 665.000000 364.090000 ;
        RECT 660.000000 367.910000 665.000000 368.090000 ;
        RECT 660.000000 371.910000 665.000000 372.090000 ;
        RECT 660.000000 375.910000 665.000000 376.090000 ;
        RECT 610.000000 395.910000 615.000000 396.090000 ;
        RECT 610.000000 391.910000 615.000000 392.090000 ;
        RECT 610.000000 387.910000 615.000000 388.090000 ;
        RECT 610.000000 383.910000 615.000000 384.090000 ;
        RECT 610.000000 399.910000 615.000000 400.090000 ;
        RECT 610.000000 403.910000 615.000000 404.090000 ;
        RECT 610.000000 407.910000 615.000000 408.090000 ;
        RECT 610.000000 411.910000 615.000000 412.090000 ;
        RECT 610.000000 415.910000 615.000000 416.090000 ;
        RECT 660.000000 383.910000 665.000000 384.090000 ;
        RECT 660.000000 387.910000 665.000000 388.090000 ;
        RECT 660.000000 391.910000 665.000000 392.090000 ;
        RECT 660.000000 395.910000 665.000000 396.090000 ;
        RECT 660.000000 403.910000 665.000000 404.090000 ;
        RECT 660.000000 399.910000 665.000000 400.090000 ;
        RECT 660.000000 407.910000 665.000000 408.090000 ;
        RECT 660.000000 411.910000 665.000000 412.090000 ;
        RECT 660.000000 415.910000 665.000000 416.090000 ;
        RECT 710.000000 379.910000 715.000000 380.090000 ;
        RECT 710.000000 343.910000 715.000000 344.090000 ;
        RECT 710.000000 347.910000 715.000000 348.090000 ;
        RECT 710.000000 351.910000 715.000000 352.090000 ;
        RECT 710.000000 355.910000 715.000000 356.090000 ;
        RECT 710.000000 359.910000 715.000000 360.090000 ;
        RECT 710.000000 367.910000 715.000000 368.090000 ;
        RECT 710.000000 363.910000 715.000000 364.090000 ;
        RECT 710.000000 375.910000 715.000000 376.090000 ;
        RECT 710.000000 371.910000 715.000000 372.090000 ;
        RECT 710.000000 383.910000 715.000000 384.090000 ;
        RECT 710.000000 387.910000 715.000000 388.090000 ;
        RECT 710.000000 391.910000 715.000000 392.090000 ;
        RECT 710.000000 395.910000 715.000000 396.090000 ;
        RECT 710.000000 403.910000 715.000000 404.090000 ;
        RECT 710.000000 399.910000 715.000000 400.090000 ;
        RECT 713.500000 415.910000 718.500000 416.090000 ;
        RECT 710.000000 411.910000 718.500000 412.090000 ;
        RECT 710.000000 407.910000 715.000000 408.090000 ;
        RECT 610.000000 431.910000 615.000000 432.090000 ;
        RECT 610.000000 427.910000 615.000000 428.090000 ;
        RECT 610.000000 423.910000 615.000000 424.090000 ;
        RECT 610.000000 419.910000 615.000000 420.090000 ;
        RECT 610.000000 435.910000 615.000000 436.090000 ;
        RECT 610.000000 439.910000 615.000000 440.090000 ;
        RECT 610.000000 443.910000 615.000000 444.090000 ;
        RECT 610.000000 447.910000 615.000000 448.090000 ;
        RECT 610.000000 451.910000 615.000000 452.090000 ;
        RECT 660.000000 419.910000 665.000000 420.090000 ;
        RECT 660.000000 423.910000 665.000000 424.090000 ;
        RECT 660.000000 427.910000 665.000000 428.090000 ;
        RECT 660.000000 431.910000 665.000000 432.090000 ;
        RECT 660.000000 439.910000 665.000000 440.090000 ;
        RECT 660.000000 435.910000 665.000000 436.090000 ;
        RECT 660.000000 443.910000 665.000000 444.090000 ;
        RECT 660.000000 447.910000 665.000000 448.090000 ;
        RECT 660.000000 451.910000 665.000000 452.090000 ;
        RECT 610.000000 455.910000 615.000000 456.090000 ;
        RECT 610.000000 459.910000 615.000000 460.090000 ;
        RECT 610.000000 463.910000 615.000000 464.090000 ;
        RECT 610.000000 467.910000 615.000000 468.090000 ;
        RECT 610.000000 471.910000 615.000000 472.090000 ;
        RECT 610.000000 475.910000 615.000000 476.090000 ;
        RECT 610.000000 479.910000 615.000000 480.090000 ;
        RECT 610.000000 483.910000 615.000000 484.090000 ;
        RECT 610.000000 487.910000 615.000000 488.090000 ;
        RECT 660.000000 459.910000 665.000000 460.090000 ;
        RECT 660.000000 455.910000 665.000000 456.090000 ;
        RECT 660.000000 463.910000 665.000000 464.090000 ;
        RECT 660.000000 467.910000 665.000000 468.090000 ;
        RECT 660.000000 471.910000 665.000000 472.090000 ;
        RECT 660.000000 479.910000 665.000000 480.090000 ;
        RECT 660.000000 475.910000 665.000000 476.090000 ;
        RECT 660.000000 487.910000 665.000000 488.090000 ;
        RECT 660.000000 483.910000 665.000000 484.090000 ;
        RECT 711.000000 423.910000 721.000000 424.090000 ;
        RECT 711.000000 419.910000 721.000000 420.090000 ;
        RECT 710.000000 431.910000 721.000000 432.090000 ;
        RECT 711.000000 427.910000 721.000000 428.090000 ;
        RECT 710.000000 435.910000 721.000000 436.090000 ;
        RECT 710.000000 439.910000 721.000000 440.090000 ;
        RECT 710.000000 443.910000 721.000000 444.090000 ;
        RECT 710.000000 451.910000 721.000000 452.090000 ;
        RECT 710.000000 447.910000 721.000000 448.090000 ;
        RECT 710.000000 455.910000 721.000000 456.090000 ;
        RECT 710.000000 459.910000 721.000000 460.090000 ;
        RECT 710.000000 471.910000 721.000000 472.090000 ;
        RECT 710.000000 463.910000 721.000000 464.090000 ;
        RECT 710.000000 467.910000 721.000000 468.090000 ;
        RECT 710.000000 475.910000 721.000000 476.090000 ;
        RECT 710.000000 479.910000 721.000000 480.090000 ;
        RECT 710.000000 483.910000 721.000000 484.090000 ;
        RECT 710.000000 487.910000 721.000000 488.090000 ;
        RECT 810.000000 379.910000 815.000000 380.090000 ;
        RECT 760.000000 379.910000 765.000000 380.090000 ;
        RECT 760.000000 343.910000 765.000000 344.090000 ;
        RECT 760.000000 347.910000 765.000000 348.090000 ;
        RECT 760.000000 351.910000 765.000000 352.090000 ;
        RECT 760.000000 355.910000 765.000000 356.090000 ;
        RECT 760.000000 359.910000 765.000000 360.090000 ;
        RECT 760.000000 363.910000 765.000000 364.090000 ;
        RECT 760.000000 367.910000 765.000000 368.090000 ;
        RECT 760.000000 375.910000 765.000000 376.090000 ;
        RECT 760.000000 371.910000 765.000000 372.090000 ;
        RECT 810.000000 343.910000 815.000000 344.090000 ;
        RECT 810.000000 347.910000 815.000000 348.090000 ;
        RECT 810.000000 351.910000 815.000000 352.090000 ;
        RECT 810.000000 359.910000 815.000000 360.090000 ;
        RECT 810.000000 355.910000 815.000000 356.090000 ;
        RECT 810.000000 363.910000 815.000000 364.090000 ;
        RECT 810.000000 367.910000 815.000000 368.090000 ;
        RECT 810.000000 371.910000 815.000000 372.090000 ;
        RECT 810.000000 375.910000 815.000000 376.090000 ;
        RECT 760.000000 395.910000 765.000000 396.090000 ;
        RECT 760.000000 391.910000 765.000000 392.090000 ;
        RECT 760.000000 387.910000 765.000000 388.090000 ;
        RECT 760.000000 383.910000 765.000000 384.090000 ;
        RECT 760.000000 399.910000 765.000000 400.090000 ;
        RECT 760.000000 403.910000 765.000000 404.090000 ;
        RECT 760.000000 407.910000 765.000000 408.090000 ;
        RECT 760.000000 411.910000 765.000000 412.090000 ;
        RECT 760.000000 415.910000 765.000000 416.090000 ;
        RECT 810.000000 387.910000 815.000000 388.090000 ;
        RECT 810.000000 383.910000 815.000000 384.090000 ;
        RECT 810.000000 391.910000 815.000000 392.090000 ;
        RECT 810.000000 395.910000 815.000000 396.090000 ;
        RECT 810.000000 403.910000 815.000000 404.090000 ;
        RECT 810.000000 399.910000 815.000000 400.090000 ;
        RECT 810.000000 407.910000 815.000000 408.090000 ;
        RECT 810.000000 411.910000 815.000000 412.090000 ;
        RECT 810.000000 415.910000 815.000000 416.090000 ;
        RECT 860.000000 379.910000 865.000000 380.090000 ;
        RECT 860.000000 359.910000 865.000000 360.090000 ;
        RECT 860.000000 355.910000 865.000000 356.090000 ;
        RECT 860.000000 351.910000 865.000000 352.090000 ;
        RECT 860.000000 347.910000 865.000000 348.090000 ;
        RECT 860.000000 343.910000 865.000000 344.090000 ;
        RECT 860.000000 363.910000 865.000000 364.090000 ;
        RECT 860.000000 367.910000 865.000000 368.090000 ;
        RECT 860.000000 371.910000 865.000000 372.090000 ;
        RECT 860.000000 375.910000 865.000000 376.090000 ;
        RECT 860.000000 383.910000 865.000000 384.090000 ;
        RECT 860.000000 387.910000 865.000000 388.090000 ;
        RECT 860.000000 391.910000 865.000000 392.090000 ;
        RECT 860.000000 395.910000 865.000000 396.090000 ;
        RECT 860.000000 403.910000 865.000000 404.090000 ;
        RECT 860.000000 399.910000 865.000000 400.090000 ;
        RECT 860.000000 415.910000 865.000000 416.090000 ;
        RECT 860.000000 411.910000 865.000000 412.090000 ;
        RECT 860.000000 407.910000 865.000000 408.090000 ;
        RECT 760.000000 419.910000 765.000000 420.090000 ;
        RECT 760.000000 423.910000 765.000000 424.090000 ;
        RECT 760.000000 427.910000 765.000000 428.090000 ;
        RECT 760.000000 431.910000 765.000000 432.090000 ;
        RECT 760.000000 435.910000 765.000000 436.090000 ;
        RECT 760.000000 439.910000 765.000000 440.090000 ;
        RECT 760.000000 443.910000 765.000000 444.090000 ;
        RECT 810.000000 419.910000 815.000000 420.090000 ;
        RECT 810.000000 423.910000 815.000000 424.090000 ;
        RECT 810.000000 431.910000 815.000000 432.090000 ;
        RECT 810.000000 427.910000 815.000000 428.090000 ;
        RECT 810.000000 435.910000 815.000000 436.090000 ;
        RECT 810.000000 439.910000 815.000000 440.090000 ;
        RECT 810.000000 443.910000 815.000000 444.090000 ;
        RECT 860.000000 419.910000 865.000000 420.090000 ;
        RECT 860.000000 423.910000 865.000000 424.090000 ;
        RECT 860.000000 427.910000 865.000000 428.090000 ;
        RECT 860.000000 431.910000 865.000000 432.090000 ;
        RECT 860.000000 443.910000 865.000000 444.090000 ;
        RECT 860.000000 439.910000 865.000000 440.090000 ;
        RECT 860.000000 435.910000 865.000000 436.090000 ;
        RECT 610.000000 491.910000 615.000000 492.090000 ;
        RECT 610.000000 499.910000 615.000000 500.090000 ;
        RECT 610.000000 495.910000 615.000000 496.090000 ;
        RECT 610.000000 503.910000 615.000000 504.090000 ;
        RECT 660.000000 495.910000 665.000000 496.090000 ;
        RECT 660.000000 491.910000 665.000000 492.090000 ;
        RECT 660.000000 499.910000 665.000000 500.090000 ;
        RECT 660.000000 503.910000 665.000000 504.090000 ;
        RECT 710.000000 503.910000 715.000000 504.090000 ;
        RECT 710.000000 499.910000 715.000000 500.090000 ;
        RECT 710.000000 495.910000 715.000000 496.090000 ;
        RECT 710.000000 491.910000 715.000000 492.090000 ;
        RECT 960.000000 379.910000 965.000000 380.090000 ;
        RECT 960.000000 343.910000 965.000000 344.090000 ;
        RECT 960.000000 347.910000 965.000000 348.090000 ;
        RECT 960.000000 351.910000 965.000000 352.090000 ;
        RECT 960.000000 359.910000 965.000000 360.090000 ;
        RECT 960.000000 355.910000 965.000000 356.090000 ;
        RECT 960.000000 375.910000 965.000000 376.090000 ;
        RECT 960.000000 371.910000 965.000000 372.090000 ;
        RECT 960.000000 367.910000 965.000000 368.090000 ;
        RECT 960.000000 363.910000 965.000000 364.090000 ;
        RECT 960.000000 383.910000 965.000000 384.090000 ;
        RECT 960.000000 387.910000 965.000000 388.090000 ;
        RECT 960.000000 391.910000 965.000000 392.090000 ;
        RECT 960.000000 395.910000 965.000000 396.090000 ;
        RECT 960.000000 399.910000 965.000000 400.090000 ;
        RECT 960.000000 403.910000 965.000000 404.090000 ;
        RECT 960.000000 407.910000 965.000000 408.090000 ;
        RECT 960.000000 411.910000 965.000000 412.090000 ;
        RECT 960.000000 415.910000 965.000000 416.090000 ;
        RECT 910.000000 379.910000 915.000000 380.090000 ;
        RECT 910.000000 343.910000 915.000000 344.090000 ;
        RECT 910.000000 347.910000 915.000000 348.090000 ;
        RECT 910.000000 351.910000 915.000000 352.090000 ;
        RECT 910.000000 355.910000 915.000000 356.090000 ;
        RECT 910.000000 359.910000 915.000000 360.090000 ;
        RECT 910.000000 363.910000 915.000000 364.090000 ;
        RECT 910.000000 367.910000 915.000000 368.090000 ;
        RECT 910.000000 371.910000 915.000000 372.090000 ;
        RECT 910.000000 375.910000 915.000000 376.090000 ;
        RECT 910.000000 395.910000 915.000000 396.090000 ;
        RECT 910.000000 391.910000 915.000000 392.090000 ;
        RECT 910.000000 387.910000 915.000000 388.090000 ;
        RECT 910.000000 383.910000 915.000000 384.090000 ;
        RECT 910.000000 399.910000 915.000000 400.090000 ;
        RECT 910.000000 403.910000 915.000000 404.090000 ;
        RECT 910.000000 407.910000 915.000000 408.090000 ;
        RECT 910.000000 411.910000 915.000000 412.090000 ;
        RECT 910.000000 415.910000 915.000000 416.090000 ;
        RECT 1010.000000 379.910000 1015.000000 380.090000 ;
        RECT 1010.000000 343.910000 1015.000000 344.090000 ;
        RECT 1010.000000 347.910000 1015.000000 348.090000 ;
        RECT 1010.000000 351.910000 1015.000000 352.090000 ;
        RECT 1010.000000 359.910000 1015.000000 360.090000 ;
        RECT 1010.000000 355.910000 1015.000000 356.090000 ;
        RECT 1010.000000 363.910000 1015.000000 364.090000 ;
        RECT 1010.000000 367.910000 1015.000000 368.090000 ;
        RECT 1010.000000 371.910000 1015.000000 372.090000 ;
        RECT 1010.000000 375.910000 1015.000000 376.090000 ;
        RECT 1010.000000 387.910000 1015.000000 388.090000 ;
        RECT 1010.000000 383.910000 1015.000000 384.090000 ;
        RECT 1010.000000 391.910000 1015.000000 392.090000 ;
        RECT 1010.000000 395.910000 1015.000000 396.090000 ;
        RECT 1010.000000 399.910000 1015.000000 400.090000 ;
        RECT 1010.000000 403.910000 1015.000000 404.090000 ;
        RECT 1010.000000 407.910000 1015.000000 408.090000 ;
        RECT 1010.000000 411.910000 1015.000000 412.090000 ;
        RECT 1010.000000 415.910000 1015.000000 416.090000 ;
        RECT 960.000000 431.910000 965.000000 432.090000 ;
        RECT 960.000000 427.910000 965.000000 428.090000 ;
        RECT 960.000000 423.910000 965.000000 424.090000 ;
        RECT 960.000000 419.910000 965.000000 420.090000 ;
        RECT 960.000000 443.910000 965.000000 444.090000 ;
        RECT 960.000000 439.910000 965.000000 440.090000 ;
        RECT 960.000000 435.910000 965.000000 436.090000 ;
        RECT 910.000000 431.910000 915.000000 432.090000 ;
        RECT 910.000000 427.910000 915.000000 428.090000 ;
        RECT 910.000000 423.910000 915.000000 424.090000 ;
        RECT 910.000000 419.910000 915.000000 420.090000 ;
        RECT 910.000000 435.910000 915.000000 436.090000 ;
        RECT 910.000000 439.910000 915.000000 440.090000 ;
        RECT 910.000000 443.910000 915.000000 444.090000 ;
        RECT 1010.000000 419.910000 1015.000000 420.090000 ;
        RECT 1010.000000 423.910000 1015.000000 424.090000 ;
        RECT 1010.000000 427.910000 1015.000000 428.090000 ;
        RECT 1010.000000 431.910000 1015.000000 432.090000 ;
        RECT 1010.000000 435.910000 1015.000000 436.090000 ;
        RECT 1010.000000 439.910000 1015.000000 440.090000 ;
        RECT 1010.000000 443.910000 1015.000000 444.090000 ;
        RECT 1110.000000 379.910000 1115.000000 380.090000 ;
        RECT 1110.000000 343.910000 1115.000000 344.090000 ;
        RECT 1110.000000 347.910000 1115.000000 348.090000 ;
        RECT 1110.000000 351.910000 1115.000000 352.090000 ;
        RECT 1110.000000 359.910000 1115.000000 360.090000 ;
        RECT 1110.000000 355.910000 1115.000000 356.090000 ;
        RECT 1110.000000 375.910000 1115.000000 376.090000 ;
        RECT 1110.000000 371.910000 1115.000000 372.090000 ;
        RECT 1110.000000 367.910000 1115.000000 368.090000 ;
        RECT 1110.000000 363.910000 1115.000000 364.090000 ;
        RECT 1110.000000 383.910000 1115.000000 384.090000 ;
        RECT 1110.000000 387.910000 1115.000000 388.090000 ;
        RECT 1110.000000 391.910000 1115.000000 392.090000 ;
        RECT 1110.000000 395.910000 1115.000000 396.090000 ;
        RECT 1110.000000 399.910000 1115.000000 400.090000 ;
        RECT 1110.000000 403.910000 1115.000000 404.090000 ;
        RECT 1110.000000 407.910000 1115.000000 408.090000 ;
        RECT 1110.000000 411.910000 1115.000000 412.090000 ;
        RECT 1110.000000 415.910000 1115.000000 416.090000 ;
        RECT 1060.000000 379.910000 1065.000000 380.090000 ;
        RECT 1060.000000 343.910000 1065.000000 344.090000 ;
        RECT 1060.000000 347.910000 1065.000000 348.090000 ;
        RECT 1060.000000 351.910000 1065.000000 352.090000 ;
        RECT 1060.000000 355.910000 1065.000000 356.090000 ;
        RECT 1060.000000 359.910000 1065.000000 360.090000 ;
        RECT 1060.000000 375.910000 1065.000000 376.090000 ;
        RECT 1060.000000 371.910000 1065.000000 372.090000 ;
        RECT 1060.000000 367.910000 1065.000000 368.090000 ;
        RECT 1060.000000 363.910000 1065.000000 364.090000 ;
        RECT 1060.000000 395.910000 1065.000000 396.090000 ;
        RECT 1060.000000 391.910000 1065.000000 392.090000 ;
        RECT 1060.000000 387.910000 1065.000000 388.090000 ;
        RECT 1060.000000 383.910000 1065.000000 384.090000 ;
        RECT 1060.000000 399.910000 1065.000000 400.090000 ;
        RECT 1060.000000 403.910000 1065.000000 404.090000 ;
        RECT 1060.000000 407.910000 1065.000000 408.090000 ;
        RECT 1060.000000 411.910000 1065.000000 412.090000 ;
        RECT 1060.000000 415.910000 1065.000000 416.090000 ;
        RECT 1158.000000 379.910000 1168.000000 380.090000 ;
        RECT 1158.000000 343.910000 1168.000000 344.090000 ;
        RECT 1158.000000 347.910000 1168.000000 348.090000 ;
        RECT 1158.000000 351.910000 1168.000000 352.090000 ;
        RECT 1158.000000 355.910000 1168.000000 356.090000 ;
        RECT 1158.000000 359.910000 1168.000000 360.090000 ;
        RECT 1158.000000 375.910000 1168.000000 376.090000 ;
        RECT 1158.000000 371.910000 1168.000000 372.090000 ;
        RECT 1158.000000 367.910000 1168.000000 368.090000 ;
        RECT 1158.000000 363.910000 1168.000000 364.090000 ;
        RECT 1158.000000 395.910000 1168.000000 396.090000 ;
        RECT 1158.000000 391.910000 1168.000000 392.090000 ;
        RECT 1158.000000 387.910000 1168.000000 388.090000 ;
        RECT 1158.000000 383.910000 1168.000000 384.090000 ;
        RECT 1158.000000 399.910000 1168.000000 400.090000 ;
        RECT 1158.000000 403.910000 1168.000000 404.090000 ;
        RECT 1158.000000 407.910000 1168.000000 408.090000 ;
        RECT 1158.000000 411.910000 1168.000000 412.090000 ;
        RECT 1158.000000 415.910000 1168.000000 416.090000 ;
        RECT 1110.000000 431.910000 1115.000000 432.090000 ;
        RECT 1110.000000 427.910000 1115.000000 428.090000 ;
        RECT 1110.000000 423.910000 1115.000000 424.090000 ;
        RECT 1110.000000 419.910000 1115.000000 420.090000 ;
        RECT 1110.000000 443.910000 1115.000000 444.090000 ;
        RECT 1110.000000 439.910000 1115.000000 440.090000 ;
        RECT 1110.000000 435.910000 1115.000000 436.090000 ;
        RECT 1060.000000 419.910000 1065.000000 420.090000 ;
        RECT 1060.000000 423.910000 1065.000000 424.090000 ;
        RECT 1060.000000 427.910000 1065.000000 428.090000 ;
        RECT 1060.000000 431.910000 1065.000000 432.090000 ;
        RECT 1060.000000 435.910000 1065.000000 436.090000 ;
        RECT 1060.000000 439.910000 1065.000000 440.090000 ;
        RECT 1060.000000 443.910000 1065.000000 444.090000 ;
        RECT 1158.000000 427.910000 1168.000000 428.090000 ;
        RECT 1158.000000 423.910000 1168.000000 424.090000 ;
        RECT 1158.000000 419.910000 1168.000000 420.090000 ;
        RECT 1160.000000 431.910000 1165.000000 432.090000 ;
        RECT 1160.000000 435.910000 1165.000000 436.090000 ;
        RECT 1160.000000 439.910000 1165.000000 440.090000 ;
        RECT 1160.000000 443.910000 1165.000000 444.090000 ;
        RECT 1160.000000 447.910000 1165.000000 448.090000 ;
        RECT 1160.000000 451.910000 1165.000000 452.090000 ;
        RECT 1160.000000 459.910000 1165.000000 460.090000 ;
        RECT 1160.000000 455.910000 1165.000000 456.090000 ;
        RECT 1160.000000 463.910000 1165.000000 464.090000 ;
        RECT 1160.000000 467.910000 1165.000000 468.090000 ;
        RECT 1160.000000 471.910000 1165.000000 472.090000 ;
        RECT 1160.000000 479.910000 1165.000000 480.090000 ;
        RECT 1160.000000 475.910000 1165.000000 476.090000 ;
        RECT 1160.000000 487.910000 1165.000000 488.090000 ;
        RECT 1160.000000 483.910000 1165.000000 484.090000 ;
        RECT 1160.000000 491.910000 1165.000000 492.090000 ;
        RECT 1160.000000 495.910000 1165.000000 496.090000 ;
        RECT 1160.000000 499.910000 1165.000000 500.090000 ;
        RECT 1160.000000 507.910000 1165.000000 508.090000 ;
        RECT 1160.000000 503.910000 1165.000000 504.090000 ;
        RECT 1160.000000 511.910000 1165.000000 512.090000 ;
        RECT 1160.000000 515.910000 1165.000000 516.090000 ;
        RECT 1160.000000 519.910000 1165.000000 520.090000 ;
        RECT 1160.000000 523.910000 1165.000000 524.090000 ;
        RECT 1160.000000 527.910000 1165.000000 528.090000 ;
        RECT 1160.000000 535.910000 1165.000000 536.090000 ;
        RECT 1160.000000 531.910000 1165.000000 532.090000 ;
        RECT 1160.000000 539.910000 1165.000000 540.090000 ;
        RECT 1160.000000 543.910000 1165.000000 544.090000 ;
        RECT 1160.000000 547.910000 1165.000000 548.090000 ;
        RECT 1160.000000 551.910000 1165.000000 552.090000 ;
        RECT 1160.000000 555.910000 1165.000000 556.090000 ;
        RECT 1160.000000 563.910000 1165.000000 564.090000 ;
        RECT 1160.000000 559.910000 1165.000000 560.090000 ;
        RECT 1160.000000 567.910000 1165.000000 568.090000 ;
        RECT 1160.000000 571.910000 1165.000000 572.090000 ;
        RECT 1160.000000 579.910000 1165.000000 580.090000 ;
        RECT 1160.000000 575.910000 1165.000000 576.090000 ;
        RECT 1160.000000 583.910000 1165.000000 584.090000 ;
        RECT 1160.000000 587.910000 1165.000000 588.090000 ;
        RECT 1160.000000 591.910000 1165.000000 592.090000 ;
        RECT 1160.000000 595.910000 1165.000000 596.090000 ;
        RECT 1160.000000 599.910000 1165.000000 600.090000 ;
        RECT 1160.000000 607.910000 1165.000000 608.090000 ;
        RECT 1160.000000 603.910000 1165.000000 604.090000 ;
        RECT 1160.000000 611.910000 1165.000000 612.090000 ;
        RECT 1160.000000 615.910000 1165.000000 616.090000 ;
        RECT 1160.000000 619.910000 1165.000000 620.090000 ;
        RECT 1160.000000 623.910000 1165.000000 624.090000 ;
        RECT 1160.000000 627.910000 1165.000000 628.090000 ;
        RECT 1160.000000 635.910000 1165.000000 636.090000 ;
        RECT 1160.000000 631.910000 1165.000000 632.090000 ;
        RECT 610.000000 659.910000 615.000000 660.090000 ;
        RECT 610.000000 663.910000 615.000000 664.090000 ;
        RECT 610.000000 667.910000 615.000000 668.090000 ;
        RECT 610.000000 671.910000 615.000000 672.090000 ;
        RECT 610.000000 675.910000 615.000000 676.090000 ;
        RECT 660.000000 663.910000 665.000000 664.090000 ;
        RECT 660.000000 659.910000 665.000000 660.090000 ;
        RECT 660.000000 667.910000 665.000000 668.090000 ;
        RECT 660.000000 671.910000 665.000000 672.090000 ;
        RECT 660.000000 675.910000 665.000000 676.090000 ;
        RECT 610.000000 683.910000 615.000000 684.090000 ;
        RECT 610.000000 679.910000 615.000000 680.090000 ;
        RECT 660.000000 683.910000 665.000000 684.090000 ;
        RECT 660.000000 679.910000 665.000000 680.090000 ;
        RECT 1160.000000 639.910000 1165.000000 640.090000 ;
        RECT 1160.000000 643.910000 1165.000000 644.090000 ;
        RECT 1160.000000 647.910000 1165.000000 648.090000 ;
        RECT 1160.000000 655.910000 1165.000000 656.090000 ;
        RECT 1160.000000 651.910000 1165.000000 652.090000 ;
        RECT 1160.000000 663.910000 1165.000000 664.090000 ;
        RECT 1160.000000 659.910000 1165.000000 660.090000 ;
        RECT 1160.000000 667.910000 1165.000000 668.090000 ;
        RECT 1160.000000 671.910000 1165.000000 672.090000 ;
        RECT 1160.000000 675.910000 1165.000000 676.090000 ;
        RECT 1160.000000 683.910000 1165.000000 684.090000 ;
        RECT 1160.000000 679.910000 1165.000000 680.090000 ;
      LAYER M3 ;
        RECT 60.000000 3.910000 65.000000 4.090000 ;
        RECT 60.000000 7.910000 65.000000 8.090000 ;
        RECT 110.000000 7.910000 115.000000 8.090000 ;
        RECT 110.000000 3.910000 115.000000 4.090000 ;
        RECT 160.000000 7.910000 165.000000 8.090000 ;
        RECT 160.000000 3.910000 165.000000 4.090000 ;
        RECT 210.000000 7.910000 215.000000 8.090000 ;
        RECT 210.000000 3.910000 215.000000 4.090000 ;
        RECT 260.000000 7.910000 265.000000 8.090000 ;
        RECT 260.000000 3.910000 265.000000 4.090000 ;
        RECT 310.000000 7.910000 315.000000 8.090000 ;
        RECT 310.000000 3.910000 315.000000 4.090000 ;
        RECT 360.000000 7.910000 365.000000 8.090000 ;
        RECT 360.000000 3.910000 365.000000 4.090000 ;
        RECT 410.000000 7.910000 415.000000 8.090000 ;
        RECT 410.000000 3.910000 415.000000 4.090000 ;
        RECT 460.000000 7.910000 465.000000 8.090000 ;
        RECT 460.000000 3.910000 465.000000 4.090000 ;
        RECT 510.000000 7.910000 515.000000 8.090000 ;
        RECT 510.000000 3.910000 515.000000 4.090000 ;
        RECT 560.000000 7.910000 565.000000 8.090000 ;
        RECT 560.000000 3.910000 565.000000 4.090000 ;
        RECT 18.000000 259.910000 28.000000 260.090000 ;
        RECT 18.000000 263.910000 28.000000 264.090000 ;
        RECT 18.000000 267.910000 28.000000 268.090000 ;
        RECT 60.000000 267.910000 65.000000 268.090000 ;
        RECT 60.000000 263.910000 65.000000 264.090000 ;
        RECT 60.000000 259.910000 65.000000 260.090000 ;
        RECT 110.000000 267.910000 115.000000 268.090000 ;
        RECT 110.000000 259.910000 115.000000 260.090000 ;
        RECT 110.000000 263.910000 115.000000 264.090000 ;
        RECT 18.000000 283.910000 28.000000 284.090000 ;
        RECT 18.000000 279.910000 28.000000 280.090000 ;
        RECT 18.000000 275.910000 28.000000 276.090000 ;
        RECT 18.000000 271.910000 28.000000 272.090000 ;
        RECT 18.000000 287.910000 28.000000 288.090000 ;
        RECT 18.000000 291.910000 28.000000 292.090000 ;
        RECT 18.000000 295.910000 28.000000 296.090000 ;
        RECT 18.000000 299.910000 28.000000 300.090000 ;
        RECT 18.000000 303.910000 28.000000 304.090000 ;
        RECT 60.000000 283.910000 65.000000 284.090000 ;
        RECT 60.000000 279.910000 65.000000 280.090000 ;
        RECT 60.000000 275.910000 65.000000 276.090000 ;
        RECT 60.000000 271.910000 65.000000 272.090000 ;
        RECT 60.000000 287.910000 65.000000 288.090000 ;
        RECT 60.000000 291.910000 65.000000 292.090000 ;
        RECT 60.000000 295.910000 65.000000 296.090000 ;
        RECT 60.000000 299.910000 65.000000 300.090000 ;
        RECT 60.000000 303.910000 65.000000 304.090000 ;
        RECT 18.000000 307.910000 28.000000 308.090000 ;
        RECT 18.000000 311.910000 28.000000 312.090000 ;
        RECT 18.000000 315.910000 28.000000 316.090000 ;
        RECT 18.000000 319.910000 28.000000 320.090000 ;
        RECT 18.000000 323.910000 28.000000 324.090000 ;
        RECT 18.000000 339.910000 28.000000 340.090000 ;
        RECT 18.000000 335.910000 28.000000 336.090000 ;
        RECT 18.000000 331.910000 28.000000 332.090000 ;
        RECT 18.000000 327.910000 28.000000 328.090000 ;
        RECT 60.000000 307.910000 65.000000 308.090000 ;
        RECT 60.000000 311.910000 65.000000 312.090000 ;
        RECT 60.000000 315.910000 65.000000 316.090000 ;
        RECT 60.000000 319.910000 65.000000 320.090000 ;
        RECT 60.000000 323.910000 65.000000 324.090000 ;
        RECT 60.000000 339.910000 65.000000 340.090000 ;
        RECT 60.000000 335.910000 65.000000 336.090000 ;
        RECT 60.000000 331.910000 65.000000 332.090000 ;
        RECT 60.000000 327.910000 65.000000 328.090000 ;
        RECT 110.000000 271.910000 115.000000 272.090000 ;
        RECT 110.000000 275.910000 115.000000 276.090000 ;
        RECT 110.000000 279.910000 115.000000 280.090000 ;
        RECT 110.000000 283.910000 115.000000 284.090000 ;
        RECT 110.000000 287.910000 115.000000 288.090000 ;
        RECT 110.000000 291.910000 115.000000 292.090000 ;
        RECT 110.000000 295.910000 115.000000 296.090000 ;
        RECT 110.000000 299.910000 115.000000 300.090000 ;
        RECT 110.000000 303.910000 115.000000 304.090000 ;
        RECT 110.000000 311.910000 115.000000 312.090000 ;
        RECT 110.000000 307.910000 115.000000 308.090000 ;
        RECT 110.000000 323.910000 115.000000 324.090000 ;
        RECT 110.000000 319.910000 115.000000 320.090000 ;
        RECT 110.000000 315.910000 115.000000 316.090000 ;
        RECT 110.000000 339.910000 115.000000 340.090000 ;
        RECT 110.000000 335.910000 115.000000 336.090000 ;
        RECT 110.000000 331.910000 115.000000 332.090000 ;
        RECT 110.000000 327.910000 115.000000 328.090000 ;
        RECT 160.000000 259.910000 165.000000 260.090000 ;
        RECT 160.000000 263.910000 165.000000 264.090000 ;
        RECT 160.000000 267.910000 165.000000 268.090000 ;
        RECT 210.000000 267.910000 215.000000 268.090000 ;
        RECT 210.000000 263.910000 215.000000 264.090000 ;
        RECT 210.000000 259.910000 215.000000 260.090000 ;
        RECT 260.000000 267.910000 265.000000 268.090000 ;
        RECT 260.000000 259.910000 265.000000 260.090000 ;
        RECT 260.000000 263.910000 265.000000 264.090000 ;
        RECT 160.000000 271.910000 165.000000 272.090000 ;
        RECT 160.000000 275.910000 165.000000 276.090000 ;
        RECT 160.000000 283.910000 165.000000 284.090000 ;
        RECT 160.000000 279.910000 165.000000 280.090000 ;
        RECT 160.000000 287.910000 165.000000 288.090000 ;
        RECT 160.000000 291.910000 165.000000 292.090000 ;
        RECT 160.000000 295.910000 165.000000 296.090000 ;
        RECT 160.000000 303.910000 165.000000 304.090000 ;
        RECT 160.000000 299.910000 165.000000 300.090000 ;
        RECT 210.000000 283.910000 215.000000 284.090000 ;
        RECT 210.000000 279.910000 215.000000 280.090000 ;
        RECT 210.000000 275.910000 215.000000 276.090000 ;
        RECT 210.000000 271.910000 215.000000 272.090000 ;
        RECT 210.000000 287.910000 215.000000 288.090000 ;
        RECT 210.000000 291.910000 215.000000 292.090000 ;
        RECT 210.000000 295.910000 215.000000 296.090000 ;
        RECT 210.000000 299.910000 215.000000 300.090000 ;
        RECT 210.000000 303.910000 215.000000 304.090000 ;
        RECT 160.000000 311.910000 165.000000 312.090000 ;
        RECT 160.000000 307.910000 165.000000 308.090000 ;
        RECT 160.000000 315.910000 165.000000 316.090000 ;
        RECT 160.000000 319.910000 165.000000 320.090000 ;
        RECT 160.000000 323.910000 165.000000 324.090000 ;
        RECT 160.000000 331.910000 165.000000 332.090000 ;
        RECT 160.000000 327.910000 165.000000 328.090000 ;
        RECT 160.000000 335.910000 165.000000 336.090000 ;
        RECT 160.000000 339.910000 165.000000 340.090000 ;
        RECT 210.000000 307.910000 215.000000 308.090000 ;
        RECT 210.000000 311.910000 215.000000 312.090000 ;
        RECT 210.000000 315.910000 215.000000 316.090000 ;
        RECT 210.000000 319.910000 215.000000 320.090000 ;
        RECT 210.000000 323.910000 215.000000 324.090000 ;
        RECT 210.000000 327.910000 215.000000 328.090000 ;
        RECT 210.000000 331.910000 215.000000 332.090000 ;
        RECT 210.000000 335.910000 215.000000 336.090000 ;
        RECT 210.000000 339.910000 215.000000 340.090000 ;
        RECT 260.000000 271.910000 265.000000 272.090000 ;
        RECT 260.000000 275.910000 265.000000 276.090000 ;
        RECT 260.000000 279.910000 265.000000 280.090000 ;
        RECT 260.000000 283.910000 265.000000 284.090000 ;
        RECT 260.000000 291.910000 265.000000 292.090000 ;
        RECT 260.000000 287.910000 265.000000 288.090000 ;
        RECT 260.000000 295.910000 265.000000 296.090000 ;
        RECT 260.000000 299.910000 265.000000 300.090000 ;
        RECT 260.000000 303.910000 265.000000 304.090000 ;
        RECT 260.000000 311.910000 265.000000 312.090000 ;
        RECT 260.000000 307.910000 265.000000 308.090000 ;
        RECT 260.000000 323.910000 265.000000 324.090000 ;
        RECT 260.000000 319.910000 265.000000 320.090000 ;
        RECT 260.000000 315.910000 265.000000 316.090000 ;
        RECT 260.000000 331.910000 265.000000 332.090000 ;
        RECT 260.000000 327.910000 265.000000 328.090000 ;
        RECT 260.000000 339.910000 265.000000 340.090000 ;
        RECT 260.000000 335.910000 265.000000 336.090000 ;
        RECT 310.000000 259.910000 315.000000 260.090000 ;
        RECT 310.000000 263.910000 315.000000 264.090000 ;
        RECT 310.000000 267.910000 315.000000 268.090000 ;
        RECT 360.000000 267.910000 365.000000 268.090000 ;
        RECT 360.000000 263.910000 365.000000 264.090000 ;
        RECT 360.000000 259.910000 365.000000 260.090000 ;
        RECT 410.000000 267.910000 415.000000 268.090000 ;
        RECT 410.000000 259.910000 415.000000 260.090000 ;
        RECT 410.000000 263.910000 415.000000 264.090000 ;
        RECT 310.000000 271.910000 315.000000 272.090000 ;
        RECT 310.000000 275.910000 315.000000 276.090000 ;
        RECT 310.000000 279.910000 315.000000 280.090000 ;
        RECT 310.000000 283.910000 315.000000 284.090000 ;
        RECT 310.000000 291.910000 315.000000 292.090000 ;
        RECT 310.000000 287.910000 315.000000 288.090000 ;
        RECT 310.000000 295.910000 315.000000 296.090000 ;
        RECT 310.000000 299.910000 315.000000 300.090000 ;
        RECT 310.000000 303.910000 315.000000 304.090000 ;
        RECT 360.000000 283.910000 365.000000 284.090000 ;
        RECT 360.000000 279.910000 365.000000 280.090000 ;
        RECT 360.000000 275.910000 365.000000 276.090000 ;
        RECT 360.000000 271.910000 365.000000 272.090000 ;
        RECT 360.000000 287.910000 365.000000 288.090000 ;
        RECT 360.000000 291.910000 365.000000 292.090000 ;
        RECT 360.000000 295.910000 365.000000 296.090000 ;
        RECT 360.000000 299.910000 365.000000 300.090000 ;
        RECT 360.000000 303.910000 365.000000 304.090000 ;
        RECT 310.000000 307.910000 315.000000 308.090000 ;
        RECT 310.000000 311.910000 315.000000 312.090000 ;
        RECT 310.000000 315.910000 315.000000 316.090000 ;
        RECT 310.000000 323.910000 315.000000 324.090000 ;
        RECT 310.000000 319.910000 315.000000 320.090000 ;
        RECT 310.000000 327.910000 315.000000 328.090000 ;
        RECT 310.000000 331.910000 315.000000 332.090000 ;
        RECT 310.000000 335.910000 315.000000 336.090000 ;
        RECT 310.000000 339.910000 315.000000 340.090000 ;
        RECT 360.000000 307.910000 365.000000 308.090000 ;
        RECT 360.000000 311.910000 365.000000 312.090000 ;
        RECT 360.000000 315.910000 365.000000 316.090000 ;
        RECT 360.000000 319.910000 365.000000 320.090000 ;
        RECT 360.000000 323.910000 365.000000 324.090000 ;
        RECT 360.000000 339.910000 365.000000 340.090000 ;
        RECT 360.000000 335.910000 365.000000 336.090000 ;
        RECT 360.000000 331.910000 365.000000 332.090000 ;
        RECT 360.000000 327.910000 365.000000 328.090000 ;
        RECT 410.000000 271.910000 415.000000 272.090000 ;
        RECT 410.000000 275.910000 415.000000 276.090000 ;
        RECT 410.000000 279.910000 415.000000 280.090000 ;
        RECT 410.000000 283.910000 415.000000 284.090000 ;
        RECT 410.000000 295.910000 415.000000 296.090000 ;
        RECT 410.000000 291.910000 415.000000 292.090000 ;
        RECT 410.000000 287.910000 415.000000 288.090000 ;
        RECT 410.000000 299.910000 415.000000 300.090000 ;
        RECT 410.000000 303.910000 415.000000 304.090000 ;
        RECT 410.000000 307.910000 415.000000 308.090000 ;
        RECT 410.000000 311.910000 415.000000 312.090000 ;
        RECT 410.000000 315.910000 415.000000 316.090000 ;
        RECT 410.000000 319.910000 415.000000 320.090000 ;
        RECT 410.000000 323.910000 415.000000 324.090000 ;
        RECT 410.000000 327.910000 415.000000 328.090000 ;
        RECT 410.000000 331.910000 415.000000 332.090000 ;
        RECT 410.000000 335.910000 415.000000 336.090000 ;
        RECT 410.000000 339.910000 415.000000 340.090000 ;
        RECT 460.000000 267.910000 465.000000 268.090000 ;
        RECT 460.000000 263.910000 465.000000 264.090000 ;
        RECT 460.000000 259.910000 465.000000 260.090000 ;
        RECT 510.000000 259.910000 515.000000 260.090000 ;
        RECT 510.000000 263.910000 515.000000 264.090000 ;
        RECT 510.000000 267.910000 515.000000 268.090000 ;
        RECT 560.000000 267.910000 565.000000 268.090000 ;
        RECT 560.000000 259.910000 565.000000 260.090000 ;
        RECT 560.000000 263.910000 565.000000 264.090000 ;
        RECT 460.000000 283.910000 465.000000 284.090000 ;
        RECT 460.000000 279.910000 465.000000 280.090000 ;
        RECT 460.000000 275.910000 465.000000 276.090000 ;
        RECT 460.000000 271.910000 465.000000 272.090000 ;
        RECT 460.000000 295.910000 465.000000 296.090000 ;
        RECT 460.000000 291.910000 465.000000 292.090000 ;
        RECT 460.000000 287.910000 465.000000 288.090000 ;
        RECT 460.000000 301.230000 465.000000 302.230000 ;
        RECT 510.000000 271.910000 515.000000 272.090000 ;
        RECT 510.000000 275.910000 515.000000 276.090000 ;
        RECT 510.000000 283.910000 515.000000 284.090000 ;
        RECT 510.000000 279.910000 515.000000 280.090000 ;
        RECT 510.000000 287.910000 515.000000 288.090000 ;
        RECT 510.000000 291.910000 515.000000 292.090000 ;
        RECT 510.000000 295.910000 515.000000 296.090000 ;
        RECT 510.000000 303.910000 515.000000 304.090000 ;
        RECT 510.000000 299.910000 515.000000 300.090000 ;
        RECT 460.000000 319.910000 465.000000 320.090000 ;
        RECT 460.000000 323.910000 465.000000 324.090000 ;
        RECT 460.000000 339.910000 465.000000 340.090000 ;
        RECT 460.000000 335.910000 465.000000 336.090000 ;
        RECT 460.000000 331.910000 465.000000 332.090000 ;
        RECT 460.000000 327.910000 465.000000 328.090000 ;
        RECT 510.000000 311.910000 515.000000 312.090000 ;
        RECT 510.000000 307.910000 515.000000 308.090000 ;
        RECT 510.000000 315.910000 515.000000 316.090000 ;
        RECT 510.000000 319.910000 515.000000 320.090000 ;
        RECT 510.000000 323.910000 515.000000 324.090000 ;
        RECT 510.000000 331.910000 515.000000 332.090000 ;
        RECT 510.000000 327.910000 515.000000 328.090000 ;
        RECT 510.000000 335.910000 515.000000 336.090000 ;
        RECT 510.000000 339.910000 515.000000 340.090000 ;
        RECT 560.000000 275.910000 565.000000 276.090000 ;
        RECT 560.000000 271.910000 565.000000 272.090000 ;
        RECT 560.000000 283.910000 565.000000 284.090000 ;
        RECT 560.000000 279.910000 565.000000 280.090000 ;
        RECT 560.000000 295.910000 565.000000 296.090000 ;
        RECT 560.000000 291.910000 565.000000 292.090000 ;
        RECT 560.000000 287.910000 565.000000 288.090000 ;
        RECT 560.000000 303.910000 565.000000 304.090000 ;
        RECT 560.000000 299.910000 565.000000 300.090000 ;
        RECT 560.000000 307.910000 565.000000 308.090000 ;
        RECT 560.000000 311.910000 565.000000 312.090000 ;
        RECT 560.000000 315.910000 565.000000 316.090000 ;
        RECT 560.000000 319.910000 565.000000 320.090000 ;
        RECT 560.000000 323.910000 565.000000 324.090000 ;
        RECT 560.000000 327.910000 565.000000 328.090000 ;
        RECT 560.000000 331.910000 565.000000 332.090000 ;
        RECT 560.000000 339.910000 565.000000 340.090000 ;
        RECT 560.000000 335.910000 565.000000 336.090000 ;
        RECT 610.000000 3.910000 615.000000 4.090000 ;
        RECT 610.000000 7.910000 615.000000 8.090000 ;
        RECT 660.000000 7.910000 665.000000 8.090000 ;
        RECT 660.000000 3.910000 665.000000 4.090000 ;
        RECT 710.000000 7.910000 715.000000 8.090000 ;
        RECT 710.000000 3.910000 715.000000 4.090000 ;
        RECT 760.000000 7.910000 765.000000 8.090000 ;
        RECT 760.000000 3.910000 765.000000 4.090000 ;
        RECT 810.000000 7.910000 815.000000 8.090000 ;
        RECT 810.000000 3.910000 815.000000 4.090000 ;
        RECT 860.000000 7.910000 865.000000 8.090000 ;
        RECT 860.000000 3.910000 865.000000 4.090000 ;
        RECT 960.000000 7.910000 965.000000 8.090000 ;
        RECT 960.000000 3.910000 965.000000 4.090000 ;
        RECT 910.000000 7.910000 915.000000 8.090000 ;
        RECT 910.000000 3.910000 915.000000 4.090000 ;
        RECT 1010.000000 7.910000 1015.000000 8.090000 ;
        RECT 1010.000000 3.910000 1015.000000 4.090000 ;
        RECT 1110.000000 7.910000 1115.000000 8.090000 ;
        RECT 1110.000000 3.910000 1115.000000 4.090000 ;
        RECT 1060.000000 7.910000 1065.000000 8.090000 ;
        RECT 1060.000000 3.910000 1065.000000 4.090000 ;
        RECT 1160.000000 3.910000 1165.000000 4.090000 ;
        RECT 1160.000000 7.910000 1165.000000 8.090000 ;
        RECT 1158.000000 27.910000 1168.000000 28.090000 ;
        RECT 1158.000000 23.910000 1168.000000 24.090000 ;
        RECT 1158.000000 19.910000 1168.000000 20.090000 ;
        RECT 1160.000000 15.910000 1165.000000 16.090000 ;
        RECT 1160.000000 11.910000 1165.000000 12.090000 ;
        RECT 1158.000000 31.910000 1168.000000 32.090000 ;
        RECT 1158.000000 35.910000 1168.000000 36.090000 ;
        RECT 1158.000000 43.910000 1168.000000 44.090000 ;
        RECT 1158.000000 39.910000 1168.000000 40.090000 ;
        RECT 610.000000 263.910000 615.000000 264.090000 ;
        RECT 610.000000 259.910000 615.000000 260.090000 ;
        RECT 610.000000 267.910000 615.000000 268.090000 ;
        RECT 660.000000 259.910000 665.000000 260.090000 ;
        RECT 660.000000 263.910000 665.000000 264.090000 ;
        RECT 660.000000 267.910000 665.000000 268.090000 ;
        RECT 710.000000 267.910000 715.000000 268.090000 ;
        RECT 710.000000 259.910000 715.000000 260.090000 ;
        RECT 710.000000 263.910000 715.000000 264.090000 ;
        RECT 610.000000 271.910000 615.000000 272.090000 ;
        RECT 610.000000 275.910000 615.000000 276.090000 ;
        RECT 610.000000 279.910000 615.000000 280.090000 ;
        RECT 610.000000 283.910000 615.000000 284.090000 ;
        RECT 610.000000 287.910000 615.000000 288.090000 ;
        RECT 610.000000 291.910000 615.000000 292.090000 ;
        RECT 610.000000 295.910000 615.000000 296.090000 ;
        RECT 610.000000 299.910000 615.000000 300.090000 ;
        RECT 610.000000 303.910000 615.000000 304.090000 ;
        RECT 660.000000 271.910000 665.000000 272.090000 ;
        RECT 660.000000 275.910000 665.000000 276.090000 ;
        RECT 660.000000 283.910000 665.000000 284.090000 ;
        RECT 660.000000 279.910000 665.000000 280.090000 ;
        RECT 660.000000 287.910000 665.000000 288.090000 ;
        RECT 660.000000 291.910000 665.000000 292.090000 ;
        RECT 660.000000 295.910000 665.000000 296.090000 ;
        RECT 660.000000 299.910000 665.000000 300.090000 ;
        RECT 660.000000 303.910000 665.000000 304.090000 ;
        RECT 610.000000 307.910000 615.000000 308.090000 ;
        RECT 610.000000 311.910000 615.000000 312.090000 ;
        RECT 610.000000 315.910000 615.000000 316.090000 ;
        RECT 610.000000 319.910000 615.000000 320.090000 ;
        RECT 610.000000 323.910000 615.000000 324.090000 ;
        RECT 610.000000 339.910000 615.000000 340.090000 ;
        RECT 610.000000 335.910000 615.000000 336.090000 ;
        RECT 610.000000 331.910000 615.000000 332.090000 ;
        RECT 610.000000 327.910000 615.000000 328.090000 ;
        RECT 660.000000 311.910000 665.000000 312.090000 ;
        RECT 660.000000 307.910000 665.000000 308.090000 ;
        RECT 660.000000 315.910000 665.000000 316.090000 ;
        RECT 660.000000 319.910000 665.000000 320.090000 ;
        RECT 660.000000 323.910000 665.000000 324.090000 ;
        RECT 660.000000 331.910000 665.000000 332.090000 ;
        RECT 660.000000 327.910000 665.000000 328.090000 ;
        RECT 660.000000 335.910000 665.000000 336.090000 ;
        RECT 660.000000 339.910000 665.000000 340.090000 ;
        RECT 710.000000 271.910000 715.000000 272.090000 ;
        RECT 710.000000 275.910000 715.000000 276.090000 ;
        RECT 710.000000 279.910000 715.000000 280.090000 ;
        RECT 710.000000 283.910000 715.000000 284.090000 ;
        RECT 710.000000 295.910000 715.000000 296.090000 ;
        RECT 710.000000 291.910000 715.000000 292.090000 ;
        RECT 710.000000 287.910000 715.000000 288.090000 ;
        RECT 710.000000 303.910000 715.000000 304.090000 ;
        RECT 710.000000 299.910000 715.000000 300.090000 ;
        RECT 710.000000 323.910000 715.000000 324.090000 ;
        RECT 710.000000 319.910000 715.000000 320.090000 ;
        RECT 710.000000 315.910000 715.000000 316.090000 ;
        RECT 710.000000 311.910000 715.000000 312.090000 ;
        RECT 710.000000 307.910000 715.000000 308.090000 ;
        RECT 710.000000 331.910000 715.000000 332.090000 ;
        RECT 710.000000 327.910000 715.000000 328.090000 ;
        RECT 710.000000 339.910000 715.000000 340.090000 ;
        RECT 710.000000 335.910000 715.000000 336.090000 ;
        RECT 760.000000 267.910000 765.000000 268.090000 ;
        RECT 760.000000 263.910000 765.000000 264.090000 ;
        RECT 760.000000 259.910000 765.000000 260.090000 ;
        RECT 810.000000 259.910000 815.000000 260.090000 ;
        RECT 810.000000 263.910000 815.000000 264.090000 ;
        RECT 810.000000 267.910000 815.000000 268.090000 ;
        RECT 860.000000 267.910000 865.000000 268.090000 ;
        RECT 860.000000 259.910000 865.000000 260.090000 ;
        RECT 860.000000 263.910000 865.000000 264.090000 ;
        RECT 760.000000 283.910000 765.000000 284.090000 ;
        RECT 760.000000 279.910000 765.000000 280.090000 ;
        RECT 760.000000 275.910000 765.000000 276.090000 ;
        RECT 760.000000 271.910000 765.000000 272.090000 ;
        RECT 760.000000 287.910000 765.000000 288.090000 ;
        RECT 760.000000 291.910000 765.000000 292.090000 ;
        RECT 760.000000 295.910000 765.000000 296.090000 ;
        RECT 760.000000 299.910000 765.000000 300.090000 ;
        RECT 760.000000 303.910000 765.000000 304.090000 ;
        RECT 810.000000 271.910000 815.000000 272.090000 ;
        RECT 810.000000 275.910000 815.000000 276.090000 ;
        RECT 810.000000 283.910000 815.000000 284.090000 ;
        RECT 810.000000 279.910000 815.000000 280.090000 ;
        RECT 810.000000 287.910000 815.000000 288.090000 ;
        RECT 810.000000 291.910000 815.000000 292.090000 ;
        RECT 810.000000 295.910000 815.000000 296.090000 ;
        RECT 810.000000 303.910000 815.000000 304.090000 ;
        RECT 810.000000 299.910000 815.000000 300.090000 ;
        RECT 760.000000 307.910000 765.000000 308.090000 ;
        RECT 760.000000 311.910000 765.000000 312.090000 ;
        RECT 760.000000 315.910000 765.000000 316.090000 ;
        RECT 760.000000 319.910000 765.000000 320.090000 ;
        RECT 760.000000 323.910000 765.000000 324.090000 ;
        RECT 760.000000 339.910000 765.000000 340.090000 ;
        RECT 760.000000 335.910000 765.000000 336.090000 ;
        RECT 760.000000 331.910000 765.000000 332.090000 ;
        RECT 760.000000 327.910000 765.000000 328.090000 ;
        RECT 810.000000 307.910000 815.000000 308.090000 ;
        RECT 810.000000 311.910000 815.000000 312.090000 ;
        RECT 810.000000 315.910000 815.000000 316.090000 ;
        RECT 810.000000 323.910000 815.000000 324.090000 ;
        RECT 810.000000 319.910000 815.000000 320.090000 ;
        RECT 810.000000 327.910000 815.000000 328.090000 ;
        RECT 810.000000 331.910000 815.000000 332.090000 ;
        RECT 810.000000 335.910000 815.000000 336.090000 ;
        RECT 810.000000 339.910000 815.000000 340.090000 ;
        RECT 860.000000 271.910000 865.000000 272.090000 ;
        RECT 860.000000 275.910000 865.000000 276.090000 ;
        RECT 860.000000 279.910000 865.000000 280.090000 ;
        RECT 860.000000 283.910000 865.000000 284.090000 ;
        RECT 860.000000 295.910000 865.000000 296.090000 ;
        RECT 860.000000 291.910000 865.000000 292.090000 ;
        RECT 860.000000 287.910000 865.000000 288.090000 ;
        RECT 860.000000 303.910000 865.000000 304.090000 ;
        RECT 860.000000 299.910000 865.000000 300.090000 ;
        RECT 860.000000 307.910000 865.000000 308.090000 ;
        RECT 860.000000 311.910000 865.000000 312.090000 ;
        RECT 860.000000 315.910000 865.000000 316.090000 ;
        RECT 860.000000 319.910000 865.000000 320.090000 ;
        RECT 860.000000 323.910000 865.000000 324.090000 ;
        RECT 860.000000 339.910000 865.000000 340.090000 ;
        RECT 860.000000 335.910000 865.000000 336.090000 ;
        RECT 860.000000 331.910000 865.000000 332.090000 ;
        RECT 860.000000 327.910000 865.000000 328.090000 ;
        RECT 1158.000000 47.910000 1168.000000 48.090000 ;
        RECT 1158.000000 51.910000 1168.000000 52.090000 ;
        RECT 1158.000000 63.910000 1168.000000 64.090000 ;
        RECT 1158.000000 55.910000 1168.000000 56.090000 ;
        RECT 1158.000000 59.910000 1168.000000 60.090000 ;
        RECT 1158.000000 67.910000 1168.000000 68.090000 ;
        RECT 1158.000000 71.910000 1168.000000 72.090000 ;
        RECT 1158.000000 79.910000 1168.000000 80.090000 ;
        RECT 1158.000000 75.910000 1168.000000 76.090000 ;
        RECT 1158.000000 83.910000 1168.000000 84.090000 ;
        RECT 1158.000000 87.910000 1168.000000 88.090000 ;
        RECT 1158.000000 91.910000 1168.000000 92.090000 ;
        RECT 1158.000000 99.910000 1168.000000 100.090000 ;
        RECT 1158.000000 95.910000 1168.000000 96.090000 ;
        RECT 1158.000000 103.910000 1168.000000 104.090000 ;
        RECT 1158.000000 107.910000 1168.000000 108.090000 ;
        RECT 1158.000000 119.910000 1168.000000 120.090000 ;
        RECT 1158.000000 115.910000 1168.000000 116.090000 ;
        RECT 1158.000000 111.910000 1168.000000 112.090000 ;
        RECT 1158.000000 123.910000 1168.000000 124.090000 ;
        RECT 1158.000000 127.910000 1168.000000 128.090000 ;
        RECT 1158.000000 135.910000 1168.000000 136.090000 ;
        RECT 1158.000000 131.910000 1168.000000 132.090000 ;
        RECT 1158.000000 139.910000 1168.000000 140.090000 ;
        RECT 1158.000000 143.910000 1168.000000 144.090000 ;
        RECT 1158.000000 147.910000 1168.000000 148.090000 ;
        RECT 1158.000000 155.910000 1168.000000 156.090000 ;
        RECT 1158.000000 151.910000 1168.000000 152.090000 ;
        RECT 1158.000000 159.910000 1168.000000 160.090000 ;
        RECT 1158.000000 163.910000 1168.000000 164.090000 ;
        RECT 1158.000000 175.910000 1168.000000 176.090000 ;
        RECT 1158.000000 171.910000 1168.000000 172.090000 ;
        RECT 1158.000000 167.910000 1168.000000 168.090000 ;
        RECT 1158.000000 179.910000 1168.000000 180.090000 ;
        RECT 1158.000000 183.910000 1168.000000 184.090000 ;
        RECT 1158.000000 191.910000 1168.000000 192.090000 ;
        RECT 1158.000000 187.910000 1168.000000 188.090000 ;
        RECT 960.000000 267.910000 965.000000 268.090000 ;
        RECT 960.000000 263.910000 965.000000 264.090000 ;
        RECT 960.000000 259.910000 965.000000 260.090000 ;
        RECT 910.000000 267.910000 915.000000 268.090000 ;
        RECT 910.000000 263.910000 915.000000 264.090000 ;
        RECT 910.000000 259.910000 915.000000 260.090000 ;
        RECT 1010.000000 259.910000 1015.000000 260.090000 ;
        RECT 1010.000000 263.910000 1015.000000 264.090000 ;
        RECT 1010.000000 267.910000 1015.000000 268.090000 ;
        RECT 960.000000 283.910000 965.000000 284.090000 ;
        RECT 960.000000 279.910000 965.000000 280.090000 ;
        RECT 960.000000 275.910000 965.000000 276.090000 ;
        RECT 960.000000 271.910000 965.000000 272.090000 ;
        RECT 960.000000 287.910000 965.000000 288.090000 ;
        RECT 960.000000 291.910000 965.000000 292.090000 ;
        RECT 960.000000 295.910000 965.000000 296.090000 ;
        RECT 960.000000 299.910000 965.000000 300.090000 ;
        RECT 960.000000 303.910000 965.000000 304.090000 ;
        RECT 960.000000 311.910000 965.000000 312.090000 ;
        RECT 960.000000 307.910000 965.000000 308.090000 ;
        RECT 960.000000 323.910000 965.000000 324.090000 ;
        RECT 960.000000 319.910000 965.000000 320.090000 ;
        RECT 960.000000 315.910000 965.000000 316.090000 ;
        RECT 960.000000 339.910000 965.000000 340.090000 ;
        RECT 960.000000 335.910000 965.000000 336.090000 ;
        RECT 960.000000 331.910000 965.000000 332.090000 ;
        RECT 960.000000 327.910000 965.000000 328.090000 ;
        RECT 910.000000 283.910000 915.000000 284.090000 ;
        RECT 910.000000 279.910000 915.000000 280.090000 ;
        RECT 910.000000 275.910000 915.000000 276.090000 ;
        RECT 910.000000 271.910000 915.000000 272.090000 ;
        RECT 910.000000 287.910000 915.000000 288.090000 ;
        RECT 910.000000 291.910000 915.000000 292.090000 ;
        RECT 910.000000 295.910000 915.000000 296.090000 ;
        RECT 910.000000 299.910000 915.000000 300.090000 ;
        RECT 910.000000 303.910000 915.000000 304.090000 ;
        RECT 910.000000 307.910000 915.000000 308.090000 ;
        RECT 910.000000 311.910000 915.000000 312.090000 ;
        RECT 910.000000 315.910000 915.000000 316.090000 ;
        RECT 910.000000 319.910000 915.000000 320.090000 ;
        RECT 910.000000 323.910000 915.000000 324.090000 ;
        RECT 910.000000 339.910000 915.000000 340.090000 ;
        RECT 910.000000 335.910000 915.000000 336.090000 ;
        RECT 910.000000 331.910000 915.000000 332.090000 ;
        RECT 910.000000 327.910000 915.000000 328.090000 ;
        RECT 1010.000000 271.910000 1015.000000 272.090000 ;
        RECT 1010.000000 275.910000 1015.000000 276.090000 ;
        RECT 1010.000000 283.910000 1015.000000 284.090000 ;
        RECT 1010.000000 279.910000 1015.000000 280.090000 ;
        RECT 1010.000000 287.910000 1015.000000 288.090000 ;
        RECT 1010.000000 291.910000 1015.000000 292.090000 ;
        RECT 1010.000000 295.910000 1015.000000 296.090000 ;
        RECT 1010.000000 303.910000 1015.000000 304.090000 ;
        RECT 1010.000000 299.910000 1015.000000 300.090000 ;
        RECT 1010.000000 311.910000 1015.000000 312.090000 ;
        RECT 1010.000000 307.910000 1015.000000 308.090000 ;
        RECT 1010.000000 315.910000 1015.000000 316.090000 ;
        RECT 1010.000000 319.910000 1015.000000 320.090000 ;
        RECT 1010.000000 323.910000 1015.000000 324.090000 ;
        RECT 1010.000000 331.910000 1015.000000 332.090000 ;
        RECT 1010.000000 327.910000 1015.000000 328.090000 ;
        RECT 1010.000000 335.910000 1015.000000 336.090000 ;
        RECT 1010.000000 339.910000 1015.000000 340.090000 ;
        RECT 1110.000000 267.910000 1115.000000 268.090000 ;
        RECT 1110.000000 263.910000 1115.000000 264.090000 ;
        RECT 1110.000000 259.910000 1115.000000 260.090000 ;
        RECT 1060.000000 267.910000 1065.000000 268.090000 ;
        RECT 1060.000000 263.910000 1065.000000 264.090000 ;
        RECT 1060.000000 259.910000 1065.000000 260.090000 ;
        RECT 1158.000000 203.910000 1168.000000 204.090000 ;
        RECT 1158.000000 195.910000 1168.000000 196.090000 ;
        RECT 1158.000000 199.910000 1168.000000 200.090000 ;
        RECT 1158.000000 211.910000 1168.000000 212.090000 ;
        RECT 1158.000000 207.910000 1168.000000 208.090000 ;
        RECT 1158.000000 215.910000 1168.000000 216.090000 ;
        RECT 1158.000000 219.910000 1168.000000 220.090000 ;
        RECT 1158.000000 227.910000 1168.000000 228.090000 ;
        RECT 1158.000000 223.910000 1168.000000 224.090000 ;
        RECT 1158.000000 231.910000 1168.000000 232.090000 ;
        RECT 1158.000000 235.910000 1168.000000 236.090000 ;
        RECT 1158.000000 239.910000 1168.000000 240.090000 ;
        RECT 1158.000000 247.910000 1168.000000 248.090000 ;
        RECT 1158.000000 243.910000 1168.000000 244.090000 ;
        RECT 1158.000000 251.910000 1168.000000 252.090000 ;
        RECT 1158.000000 255.910000 1168.000000 256.090000 ;
        RECT 1158.000000 267.910000 1168.000000 268.090000 ;
        RECT 1158.000000 259.910000 1168.000000 260.090000 ;
        RECT 1158.000000 263.910000 1168.000000 264.090000 ;
        RECT 1110.000000 283.910000 1115.000000 284.090000 ;
        RECT 1110.000000 279.910000 1115.000000 280.090000 ;
        RECT 1110.000000 275.910000 1115.000000 276.090000 ;
        RECT 1110.000000 271.910000 1115.000000 272.090000 ;
        RECT 1110.000000 287.910000 1115.000000 288.090000 ;
        RECT 1110.000000 291.910000 1115.000000 292.090000 ;
        RECT 1110.000000 295.910000 1115.000000 296.090000 ;
        RECT 1110.000000 299.910000 1115.000000 300.090000 ;
        RECT 1110.000000 303.910000 1115.000000 304.090000 ;
        RECT 1110.000000 311.910000 1115.000000 312.090000 ;
        RECT 1110.000000 307.910000 1115.000000 308.090000 ;
        RECT 1110.000000 323.910000 1115.000000 324.090000 ;
        RECT 1110.000000 319.910000 1115.000000 320.090000 ;
        RECT 1110.000000 315.910000 1115.000000 316.090000 ;
        RECT 1110.000000 339.910000 1115.000000 340.090000 ;
        RECT 1110.000000 335.910000 1115.000000 336.090000 ;
        RECT 1110.000000 331.910000 1115.000000 332.090000 ;
        RECT 1110.000000 327.910000 1115.000000 328.090000 ;
        RECT 1060.000000 283.910000 1065.000000 284.090000 ;
        RECT 1060.000000 279.910000 1065.000000 280.090000 ;
        RECT 1060.000000 275.910000 1065.000000 276.090000 ;
        RECT 1060.000000 271.910000 1065.000000 272.090000 ;
        RECT 1060.000000 287.910000 1065.000000 288.090000 ;
        RECT 1060.000000 291.910000 1065.000000 292.090000 ;
        RECT 1060.000000 295.910000 1065.000000 296.090000 ;
        RECT 1060.000000 299.910000 1065.000000 300.090000 ;
        RECT 1060.000000 303.910000 1065.000000 304.090000 ;
        RECT 1060.000000 307.910000 1065.000000 308.090000 ;
        RECT 1060.000000 311.910000 1065.000000 312.090000 ;
        RECT 1060.000000 315.910000 1065.000000 316.090000 ;
        RECT 1060.000000 319.910000 1065.000000 320.090000 ;
        RECT 1060.000000 323.910000 1065.000000 324.090000 ;
        RECT 1060.000000 339.910000 1065.000000 340.090000 ;
        RECT 1060.000000 335.910000 1065.000000 336.090000 ;
        RECT 1060.000000 331.910000 1065.000000 332.090000 ;
        RECT 1060.000000 327.910000 1065.000000 328.090000 ;
        RECT 1158.000000 283.910000 1168.000000 284.090000 ;
        RECT 1158.000000 279.910000 1168.000000 280.090000 ;
        RECT 1158.000000 275.910000 1168.000000 276.090000 ;
        RECT 1158.000000 271.910000 1168.000000 272.090000 ;
        RECT 1158.000000 287.910000 1168.000000 288.090000 ;
        RECT 1158.000000 291.910000 1168.000000 292.090000 ;
        RECT 1158.000000 295.910000 1168.000000 296.090000 ;
        RECT 1158.000000 299.910000 1168.000000 300.090000 ;
        RECT 1158.000000 303.910000 1168.000000 304.090000 ;
        RECT 1158.000000 307.910000 1168.000000 308.090000 ;
        RECT 1158.000000 311.910000 1168.000000 312.090000 ;
        RECT 1158.000000 315.910000 1168.000000 316.090000 ;
        RECT 1158.000000 319.910000 1168.000000 320.090000 ;
        RECT 1158.000000 323.910000 1168.000000 324.090000 ;
        RECT 1158.000000 339.910000 1168.000000 340.090000 ;
        RECT 1158.000000 335.910000 1168.000000 336.090000 ;
        RECT 1158.000000 331.910000 1168.000000 332.090000 ;
        RECT 1158.000000 327.910000 1168.000000 328.090000 ;
        RECT 60.000000 379.910000 65.000000 380.090000 ;
        RECT 18.000000 379.910000 28.000000 380.090000 ;
        RECT 18.000000 343.910000 28.000000 344.090000 ;
        RECT 18.000000 347.910000 28.000000 348.090000 ;
        RECT 18.000000 351.910000 28.000000 352.090000 ;
        RECT 18.000000 359.910000 28.000000 360.090000 ;
        RECT 18.000000 355.910000 28.000000 356.090000 ;
        RECT 18.000000 375.910000 28.000000 376.090000 ;
        RECT 18.000000 371.910000 28.000000 372.090000 ;
        RECT 18.000000 367.910000 28.000000 368.090000 ;
        RECT 18.000000 363.910000 28.000000 364.090000 ;
        RECT 60.000000 347.910000 65.000000 348.090000 ;
        RECT 60.000000 343.910000 65.000000 344.090000 ;
        RECT 60.000000 352.445000 64.080000 352.745000 ;
        RECT 60.000000 375.910000 65.000000 376.090000 ;
        RECT 60.000000 371.910000 65.000000 372.090000 ;
        RECT 60.000000 367.910000 65.000000 368.090000 ;
        RECT 60.000000 363.910000 65.000000 364.090000 ;
        RECT 18.000000 395.910000 28.000000 396.090000 ;
        RECT 18.000000 391.910000 28.000000 392.090000 ;
        RECT 18.000000 387.910000 28.000000 388.090000 ;
        RECT 18.000000 383.910000 28.000000 384.090000 ;
        RECT 18.000000 399.910000 28.000000 400.090000 ;
        RECT 18.000000 403.910000 28.000000 404.090000 ;
        RECT 18.000000 407.910000 28.000000 408.090000 ;
        RECT 18.000000 411.910000 28.000000 412.090000 ;
        RECT 18.000000 415.910000 28.000000 416.090000 ;
        RECT 60.000000 395.910000 65.000000 396.090000 ;
        RECT 60.000000 391.910000 65.000000 392.090000 ;
        RECT 60.000000 387.910000 65.000000 388.090000 ;
        RECT 60.000000 383.910000 65.000000 384.090000 ;
        RECT 60.000000 399.910000 65.000000 400.090000 ;
        RECT 60.000000 403.910000 65.000000 404.090000 ;
        RECT 60.000000 407.910000 65.000000 408.090000 ;
        RECT 60.000000 411.910000 65.000000 412.090000 ;
        RECT 60.000000 415.910000 65.000000 416.090000 ;
        RECT 110.000000 379.910000 115.000000 380.090000 ;
        RECT 110.000000 351.910000 115.000000 352.090000 ;
        RECT 110.000000 347.910000 115.000000 348.090000 ;
        RECT 110.000000 343.910000 115.000000 344.090000 ;
        RECT 110.000000 359.910000 115.000000 360.090000 ;
        RECT 110.000000 355.910000 115.000000 356.090000 ;
        RECT 110.000000 375.910000 115.000000 376.090000 ;
        RECT 110.000000 371.910000 115.000000 372.090000 ;
        RECT 110.000000 367.910000 115.000000 368.090000 ;
        RECT 110.000000 363.910000 115.000000 364.090000 ;
        RECT 110.000000 383.910000 115.000000 384.090000 ;
        RECT 110.000000 387.910000 115.000000 388.090000 ;
        RECT 110.000000 391.910000 115.000000 392.090000 ;
        RECT 110.000000 395.910000 115.000000 396.090000 ;
        RECT 110.000000 399.910000 115.000000 400.090000 ;
        RECT 110.000000 403.910000 115.000000 404.090000 ;
        RECT 110.000000 407.910000 115.000000 408.090000 ;
        RECT 110.000000 411.910000 115.000000 412.090000 ;
        RECT 110.000000 415.910000 115.000000 416.090000 ;
        RECT 18.000000 431.910000 28.000000 432.090000 ;
        RECT 18.000000 427.910000 28.000000 428.090000 ;
        RECT 18.000000 423.910000 28.000000 424.090000 ;
        RECT 18.000000 419.910000 28.000000 420.090000 ;
        RECT 18.000000 435.910000 28.000000 436.090000 ;
        RECT 18.000000 439.910000 28.000000 440.090000 ;
        RECT 18.000000 443.910000 28.000000 444.090000 ;
        RECT 18.000000 447.910000 28.000000 448.090000 ;
        RECT 18.000000 451.910000 28.000000 452.090000 ;
        RECT 60.000000 431.910000 65.000000 432.090000 ;
        RECT 60.000000 427.910000 65.000000 428.090000 ;
        RECT 60.000000 423.910000 65.000000 424.090000 ;
        RECT 60.000000 419.910000 65.000000 420.090000 ;
        RECT 60.000000 435.910000 65.000000 436.090000 ;
        RECT 60.000000 439.910000 65.000000 440.090000 ;
        RECT 60.000000 443.910000 65.000000 444.090000 ;
        RECT 60.000000 447.910000 65.000000 448.090000 ;
        RECT 60.000000 451.910000 65.000000 452.090000 ;
        RECT 18.000000 455.910000 28.000000 456.090000 ;
        RECT 18.000000 459.910000 28.000000 460.090000 ;
        RECT 18.000000 463.910000 28.000000 464.090000 ;
        RECT 18.000000 467.910000 28.000000 468.090000 ;
        RECT 18.000000 471.910000 28.000000 472.090000 ;
        RECT 18.000000 487.910000 28.000000 488.090000 ;
        RECT 18.000000 483.910000 28.000000 484.090000 ;
        RECT 18.000000 479.910000 28.000000 480.090000 ;
        RECT 18.000000 475.910000 28.000000 476.090000 ;
        RECT 60.000000 455.910000 65.000000 456.090000 ;
        RECT 60.000000 459.910000 65.000000 460.090000 ;
        RECT 60.000000 463.910000 65.000000 464.090000 ;
        RECT 60.000000 467.910000 65.000000 468.090000 ;
        RECT 60.000000 471.910000 65.000000 472.090000 ;
        RECT 60.000000 487.910000 65.000000 488.090000 ;
        RECT 60.000000 483.910000 65.000000 484.090000 ;
        RECT 60.000000 479.910000 65.000000 480.090000 ;
        RECT 60.000000 475.910000 65.000000 476.090000 ;
        RECT 110.000000 419.910000 115.000000 420.090000 ;
        RECT 110.000000 423.910000 115.000000 424.090000 ;
        RECT 110.000000 427.910000 115.000000 428.090000 ;
        RECT 110.000000 431.910000 115.000000 432.090000 ;
        RECT 110.000000 435.910000 115.000000 436.090000 ;
        RECT 110.000000 439.910000 115.000000 440.090000 ;
        RECT 110.000000 443.910000 115.000000 444.090000 ;
        RECT 110.000000 447.910000 115.000000 448.090000 ;
        RECT 110.000000 451.910000 115.000000 452.090000 ;
        RECT 110.000000 459.910000 115.000000 460.090000 ;
        RECT 110.000000 455.910000 115.000000 456.090000 ;
        RECT 110.000000 471.910000 115.000000 472.090000 ;
        RECT 110.000000 467.910000 115.000000 468.090000 ;
        RECT 110.000000 463.910000 115.000000 464.090000 ;
        RECT 110.000000 487.910000 115.000000 488.090000 ;
        RECT 110.000000 483.910000 115.000000 484.090000 ;
        RECT 110.000000 479.910000 115.000000 480.090000 ;
        RECT 110.000000 475.910000 115.000000 476.090000 ;
        RECT 210.000000 379.910000 215.000000 380.090000 ;
        RECT 160.000000 379.910000 165.000000 380.090000 ;
        RECT 160.000000 343.910000 165.000000 344.090000 ;
        RECT 160.000000 347.910000 165.000000 348.090000 ;
        RECT 160.000000 351.910000 165.000000 352.090000 ;
        RECT 160.000000 359.910000 165.000000 360.090000 ;
        RECT 160.000000 355.910000 165.000000 356.090000 ;
        RECT 160.000000 363.910000 165.000000 364.090000 ;
        RECT 160.000000 367.910000 165.000000 368.090000 ;
        RECT 160.000000 371.910000 165.000000 372.090000 ;
        RECT 160.000000 375.910000 165.000000 376.090000 ;
        RECT 210.000000 343.910000 215.000000 344.090000 ;
        RECT 210.000000 347.910000 215.000000 348.090000 ;
        RECT 210.000000 351.910000 215.000000 352.090000 ;
        RECT 210.000000 355.910000 215.000000 356.090000 ;
        RECT 210.000000 359.910000 215.000000 360.090000 ;
        RECT 210.000000 375.910000 215.000000 376.090000 ;
        RECT 210.000000 371.910000 215.000000 372.090000 ;
        RECT 210.000000 367.910000 215.000000 368.090000 ;
        RECT 210.000000 363.910000 215.000000 364.090000 ;
        RECT 160.000000 383.910000 165.000000 384.090000 ;
        RECT 160.000000 387.910000 165.000000 388.090000 ;
        RECT 160.000000 391.910000 165.000000 392.090000 ;
        RECT 160.000000 395.910000 165.000000 396.090000 ;
        RECT 160.000000 403.910000 165.000000 404.090000 ;
        RECT 160.000000 399.910000 165.000000 400.090000 ;
        RECT 160.000000 407.910000 165.000000 408.090000 ;
        RECT 210.000000 383.910000 215.000000 384.090000 ;
        RECT 210.000000 387.910000 215.000000 388.090000 ;
        RECT 210.000000 391.910000 215.000000 392.090000 ;
        RECT 210.000000 395.910000 215.000000 396.090000 ;
        RECT 210.000000 399.910000 215.000000 400.090000 ;
        RECT 210.000000 403.910000 215.000000 404.090000 ;
        RECT 210.000000 407.910000 215.000000 408.090000 ;
        RECT 210.000000 411.910000 215.000000 412.090000 ;
        RECT 210.000000 415.910000 215.000000 416.090000 ;
        RECT 260.000000 379.910000 265.000000 380.090000 ;
        RECT 260.000000 351.910000 265.000000 352.090000 ;
        RECT 260.000000 347.910000 265.000000 348.090000 ;
        RECT 260.000000 343.910000 265.000000 344.090000 ;
        RECT 260.000000 359.910000 265.000000 360.090000 ;
        RECT 260.000000 355.910000 265.000000 356.090000 ;
        RECT 260.000000 367.910000 265.000000 368.090000 ;
        RECT 260.000000 363.910000 265.000000 364.090000 ;
        RECT 260.000000 375.910000 265.000000 376.090000 ;
        RECT 260.000000 371.910000 265.000000 372.090000 ;
        RECT 260.000000 383.910000 265.000000 384.090000 ;
        RECT 260.000000 387.910000 265.000000 388.090000 ;
        RECT 260.000000 391.910000 265.000000 392.090000 ;
        RECT 260.000000 395.910000 265.000000 396.090000 ;
        RECT 260.000000 399.910000 265.000000 400.090000 ;
        RECT 260.000000 403.910000 265.000000 404.090000 ;
        RECT 260.000000 407.910000 265.000000 408.090000 ;
        RECT 210.000000 431.910000 215.000000 432.090000 ;
        RECT 210.000000 427.910000 215.000000 428.090000 ;
        RECT 210.000000 423.910000 215.000000 424.090000 ;
        RECT 210.000000 419.910000 215.000000 420.090000 ;
        RECT 210.000000 435.910000 215.000000 436.090000 ;
        RECT 210.000000 439.910000 215.000000 440.090000 ;
        RECT 210.000000 443.910000 215.000000 444.090000 ;
        RECT 210.000000 447.910000 215.000000 448.090000 ;
        RECT 210.000000 451.910000 215.000000 452.090000 ;
        RECT 160.000000 463.910000 165.000000 464.090000 ;
        RECT 160.000000 467.910000 165.000000 468.090000 ;
        RECT 160.000000 471.910000 165.000000 472.090000 ;
        RECT 160.000000 479.910000 165.000000 480.090000 ;
        RECT 160.000000 475.910000 165.000000 476.090000 ;
        RECT 160.000000 487.910000 165.000000 488.090000 ;
        RECT 160.000000 483.910000 165.000000 484.090000 ;
        RECT 210.000000 455.910000 215.000000 456.090000 ;
        RECT 210.000000 459.910000 215.000000 460.090000 ;
        RECT 210.000000 467.910000 215.000000 468.090000 ;
        RECT 210.000000 463.910000 215.000000 464.090000 ;
        RECT 210.000000 471.910000 215.000000 472.090000 ;
        RECT 210.000000 487.910000 215.000000 488.090000 ;
        RECT 210.000000 483.910000 215.000000 484.090000 ;
        RECT 210.000000 479.910000 215.000000 480.090000 ;
        RECT 210.000000 475.910000 215.000000 476.090000 ;
        RECT 260.000000 471.910000 265.000000 472.090000 ;
        RECT 260.000000 467.910000 265.000000 468.090000 ;
        RECT 260.000000 463.910000 265.000000 464.090000 ;
        RECT 260.000000 479.910000 265.000000 480.090000 ;
        RECT 260.000000 475.910000 265.000000 476.090000 ;
        RECT 260.000000 483.910000 265.000000 484.090000 ;
        RECT 260.000000 487.910000 265.000000 488.090000 ;
        RECT 18.000000 491.910000 28.000000 492.090000 ;
        RECT 18.000000 495.910000 28.000000 496.090000 ;
        RECT 18.000000 499.910000 28.000000 500.090000 ;
        RECT 18.000000 503.910000 28.000000 504.090000 ;
        RECT 18.000000 507.910000 28.000000 508.090000 ;
        RECT 18.000000 515.910000 28.000000 516.090000 ;
        RECT 18.000000 511.910000 28.000000 512.090000 ;
        RECT 60.000000 491.910000 65.000000 492.090000 ;
        RECT 60.000000 495.910000 65.000000 496.090000 ;
        RECT 60.000000 499.910000 65.000000 500.090000 ;
        RECT 60.000000 503.910000 65.000000 504.090000 ;
        RECT 60.000000 507.910000 65.000000 508.090000 ;
        RECT 60.000000 515.910000 65.000000 516.090000 ;
        RECT 60.000000 511.910000 65.000000 512.090000 ;
        RECT 110.000000 499.910000 115.000000 500.090000 ;
        RECT 110.000000 495.910000 115.000000 496.090000 ;
        RECT 110.000000 491.910000 115.000000 492.090000 ;
        RECT 110.000000 507.910000 115.000000 508.090000 ;
        RECT 110.000000 503.910000 115.000000 504.090000 ;
        RECT 110.000000 515.910000 115.000000 516.090000 ;
        RECT 110.000000 511.910000 115.000000 512.090000 ;
        RECT 160.000000 491.910000 165.000000 492.090000 ;
        RECT 160.000000 495.910000 165.000000 496.090000 ;
        RECT 160.000000 499.910000 165.000000 500.090000 ;
        RECT 160.000000 507.910000 165.000000 508.090000 ;
        RECT 160.000000 503.910000 165.000000 504.090000 ;
        RECT 160.000000 511.910000 165.000000 512.090000 ;
        RECT 160.000000 515.910000 165.000000 516.090000 ;
        RECT 210.000000 491.910000 215.000000 492.090000 ;
        RECT 210.000000 495.910000 215.000000 496.090000 ;
        RECT 210.000000 499.910000 215.000000 500.090000 ;
        RECT 210.000000 503.910000 215.000000 504.090000 ;
        RECT 210.000000 507.910000 215.000000 508.090000 ;
        RECT 210.000000 515.910000 215.000000 516.090000 ;
        RECT 210.000000 511.910000 215.000000 512.090000 ;
        RECT 260.000000 491.910000 265.000000 492.090000 ;
        RECT 260.000000 495.910000 265.000000 496.090000 ;
        RECT 260.000000 499.910000 265.000000 500.090000 ;
        RECT 260.000000 503.910000 265.000000 504.090000 ;
        RECT 260.000000 507.910000 265.000000 508.090000 ;
        RECT 260.000000 511.910000 265.000000 512.090000 ;
        RECT 260.000000 515.910000 265.000000 516.090000 ;
        RECT 310.000000 379.910000 315.000000 380.090000 ;
        RECT 360.000000 379.910000 365.000000 380.090000 ;
        RECT 310.000000 343.910000 315.000000 344.090000 ;
        RECT 310.000000 351.910000 315.000000 352.090000 ;
        RECT 310.000000 347.910000 315.000000 348.090000 ;
        RECT 310.000000 355.910000 315.000000 356.090000 ;
        RECT 310.000000 359.910000 315.000000 360.090000 ;
        RECT 310.000000 363.910000 315.000000 364.090000 ;
        RECT 310.000000 367.910000 315.000000 368.090000 ;
        RECT 310.000000 371.910000 315.000000 372.090000 ;
        RECT 310.000000 375.910000 315.000000 376.090000 ;
        RECT 360.000000 343.910000 365.000000 344.090000 ;
        RECT 360.000000 347.910000 365.000000 348.090000 ;
        RECT 360.000000 351.910000 365.000000 352.090000 ;
        RECT 360.000000 355.910000 365.000000 356.090000 ;
        RECT 360.000000 359.910000 365.000000 360.090000 ;
        RECT 360.000000 363.910000 365.000000 364.090000 ;
        RECT 360.000000 367.910000 365.000000 368.090000 ;
        RECT 360.000000 371.910000 365.000000 372.090000 ;
        RECT 360.000000 375.910000 365.000000 376.090000 ;
        RECT 310.000000 383.910000 315.000000 384.090000 ;
        RECT 310.000000 387.910000 315.000000 388.090000 ;
        RECT 310.000000 391.910000 315.000000 392.090000 ;
        RECT 310.000000 395.910000 315.000000 396.090000 ;
        RECT 310.000000 399.910000 315.000000 400.090000 ;
        RECT 310.000000 403.910000 315.000000 404.090000 ;
        RECT 310.000000 411.910000 315.000000 412.090000 ;
        RECT 310.000000 407.910000 315.000000 408.090000 ;
        RECT 310.000000 415.910000 315.000000 416.090000 ;
        RECT 360.000000 383.910000 365.000000 384.090000 ;
        RECT 360.000000 387.910000 365.000000 388.090000 ;
        RECT 360.000000 391.910000 365.000000 392.090000 ;
        RECT 360.000000 395.910000 365.000000 396.090000 ;
        RECT 360.000000 399.910000 365.000000 400.090000 ;
        RECT 360.000000 403.910000 365.000000 404.090000 ;
        RECT 360.000000 407.910000 365.000000 408.090000 ;
        RECT 360.000000 411.910000 365.000000 412.090000 ;
        RECT 360.000000 415.910000 365.000000 416.090000 ;
        RECT 410.000000 379.910000 415.000000 380.090000 ;
        RECT 410.000000 343.910000 415.000000 344.090000 ;
        RECT 410.000000 347.910000 415.000000 348.090000 ;
        RECT 410.000000 351.910000 415.000000 352.090000 ;
        RECT 410.000000 355.910000 415.000000 356.090000 ;
        RECT 410.000000 359.910000 415.000000 360.090000 ;
        RECT 410.000000 363.910000 415.000000 364.090000 ;
        RECT 410.000000 367.910000 415.000000 368.090000 ;
        RECT 410.000000 371.910000 415.000000 372.090000 ;
        RECT 410.000000 375.910000 415.000000 376.090000 ;
        RECT 410.000000 383.910000 415.000000 384.090000 ;
        RECT 410.000000 387.910000 415.000000 388.090000 ;
        RECT 410.000000 391.910000 415.000000 392.090000 ;
        RECT 410.000000 395.910000 415.000000 396.090000 ;
        RECT 410.000000 399.910000 415.000000 400.090000 ;
        RECT 410.000000 403.910000 415.000000 404.090000 ;
        RECT 410.000000 411.910000 415.000000 412.090000 ;
        RECT 410.000000 407.910000 415.000000 408.090000 ;
        RECT 410.000000 415.910000 415.000000 416.090000 ;
        RECT 361.000000 479.910000 371.000000 480.090000 ;
        RECT 361.000000 483.910000 371.000000 484.090000 ;
        RECT 361.000000 487.910000 371.000000 488.090000 ;
        RECT 310.000000 419.910000 315.000000 420.090000 ;
        RECT 310.000000 423.910000 315.000000 424.090000 ;
        RECT 310.000000 427.910000 315.000000 428.090000 ;
        RECT 310.000000 431.910000 315.000000 432.090000 ;
        RECT 310.000000 439.910000 315.000000 440.090000 ;
        RECT 310.000000 435.910000 315.000000 436.090000 ;
        RECT 310.000000 443.910000 315.000000 444.090000 ;
        RECT 310.000000 447.910000 315.000000 448.090000 ;
        RECT 310.000000 451.910000 315.000000 452.090000 ;
        RECT 360.000000 419.910000 365.000000 420.090000 ;
        RECT 360.000000 423.910000 365.000000 424.090000 ;
        RECT 360.000000 427.910000 365.000000 428.090000 ;
        RECT 360.000000 431.910000 365.000000 432.090000 ;
        RECT 360.000000 435.910000 365.000000 436.090000 ;
        RECT 360.000000 439.910000 365.000000 440.090000 ;
        RECT 360.000000 443.910000 365.000000 444.090000 ;
        RECT 360.000000 447.910000 365.000000 448.090000 ;
        RECT 360.000000 451.910000 365.000000 452.090000 ;
        RECT 310.000000 455.910000 315.000000 456.090000 ;
        RECT 310.000000 459.910000 315.000000 460.090000 ;
        RECT 310.000000 467.910000 315.000000 468.090000 ;
        RECT 310.000000 463.910000 315.000000 464.090000 ;
        RECT 310.000000 471.910000 315.000000 472.090000 ;
        RECT 310.000000 475.910000 315.000000 476.090000 ;
        RECT 310.000000 479.910000 315.000000 480.090000 ;
        RECT 310.000000 487.910000 315.000000 488.090000 ;
        RECT 310.000000 483.910000 315.000000 484.090000 ;
        RECT 360.000000 455.910000 365.000000 456.090000 ;
        RECT 360.000000 459.910000 365.000000 460.090000 ;
        RECT 360.000000 471.910000 368.500000 472.090000 ;
        RECT 360.000000 463.910000 365.000000 464.090000 ;
        RECT 360.000000 467.910000 365.000000 468.090000 ;
        RECT 363.500000 475.910000 368.500000 476.090000 ;
        RECT 410.000000 419.910000 415.000000 420.090000 ;
        RECT 410.000000 423.910000 415.000000 424.090000 ;
        RECT 410.000000 427.910000 415.000000 428.090000 ;
        RECT 410.000000 431.910000 415.000000 432.090000 ;
        RECT 410.000000 439.910000 415.000000 440.090000 ;
        RECT 410.000000 435.910000 415.000000 436.090000 ;
        RECT 410.000000 443.910000 415.000000 444.090000 ;
        RECT 410.000000 451.910000 415.000000 452.090000 ;
        RECT 410.000000 447.910000 415.000000 448.090000 ;
        RECT 410.000000 455.910000 415.000000 456.090000 ;
        RECT 410.000000 459.910000 415.000000 460.090000 ;
        RECT 410.000000 467.910000 415.000000 468.090000 ;
        RECT 410.000000 463.910000 415.000000 464.090000 ;
        RECT 410.000000 471.910000 415.000000 472.090000 ;
        RECT 410.000000 475.910000 415.000000 476.090000 ;
        RECT 410.000000 479.910000 415.000000 480.090000 ;
        RECT 410.000000 483.910000 415.000000 484.090000 ;
        RECT 410.000000 487.910000 415.000000 488.090000 ;
        RECT 460.000000 379.910000 465.000000 380.090000 ;
        RECT 510.000000 379.910000 515.000000 380.090000 ;
        RECT 460.000000 347.910000 465.000000 348.090000 ;
        RECT 460.000000 343.910000 465.000000 344.090000 ;
        RECT 460.000000 351.230000 465.000000 352.230000 ;
        RECT 460.000000 375.910000 465.000000 376.090000 ;
        RECT 460.000000 371.910000 465.000000 372.090000 ;
        RECT 510.000000 343.910000 515.000000 344.090000 ;
        RECT 510.000000 351.910000 515.000000 352.090000 ;
        RECT 510.000000 347.910000 515.000000 348.090000 ;
        RECT 510.000000 359.910000 515.000000 360.090000 ;
        RECT 510.000000 355.910000 515.000000 356.090000 ;
        RECT 510.000000 363.910000 515.000000 364.090000 ;
        RECT 510.000000 367.910000 515.000000 368.090000 ;
        RECT 510.000000 375.910000 515.000000 376.090000 ;
        RECT 510.000000 371.910000 515.000000 372.090000 ;
        RECT 460.000000 383.910000 465.000000 384.090000 ;
        RECT 460.000000 387.910000 465.000000 388.090000 ;
        RECT 460.000000 391.910000 465.000000 392.090000 ;
        RECT 460.000000 395.910000 465.000000 396.090000 ;
        RECT 460.000000 401.230000 465.000000 402.230000 ;
        RECT 510.000000 383.910000 515.000000 384.090000 ;
        RECT 510.000000 387.910000 515.000000 388.090000 ;
        RECT 510.000000 391.910000 515.000000 392.090000 ;
        RECT 510.000000 395.910000 515.000000 396.090000 ;
        RECT 510.000000 399.910000 515.000000 400.090000 ;
        RECT 510.000000 403.910000 515.000000 404.090000 ;
        RECT 510.000000 407.910000 515.000000 408.090000 ;
        RECT 510.000000 411.910000 515.000000 412.090000 ;
        RECT 510.000000 415.910000 515.000000 416.090000 ;
        RECT 560.000000 379.910000 565.000000 380.090000 ;
        RECT 560.000000 343.910000 565.000000 344.090000 ;
        RECT 560.000000 347.910000 565.000000 348.090000 ;
        RECT 560.000000 351.910000 565.000000 352.090000 ;
        RECT 560.000000 355.910000 565.000000 356.090000 ;
        RECT 560.000000 359.910000 565.000000 360.090000 ;
        RECT 560.000000 363.910000 565.000000 364.090000 ;
        RECT 560.000000 367.910000 565.000000 368.090000 ;
        RECT 560.000000 371.910000 565.000000 372.090000 ;
        RECT 560.000000 375.910000 565.000000 376.090000 ;
        RECT 560.000000 383.910000 565.000000 384.090000 ;
        RECT 560.000000 387.910000 565.000000 388.090000 ;
        RECT 560.000000 391.910000 565.000000 392.090000 ;
        RECT 560.000000 395.910000 565.000000 396.090000 ;
        RECT 560.000000 403.910000 565.000000 404.090000 ;
        RECT 560.000000 399.910000 565.000000 400.090000 ;
        RECT 560.000000 411.910000 565.000000 412.090000 ;
        RECT 560.000000 407.910000 565.000000 408.090000 ;
        RECT 560.000000 415.910000 565.000000 416.090000 ;
        RECT 460.000000 423.910000 465.000000 424.090000 ;
        RECT 460.000000 419.910000 465.000000 420.090000 ;
        RECT 460.000000 427.910000 465.000000 428.090000 ;
        RECT 460.000000 431.910000 465.000000 432.090000 ;
        RECT 460.000000 435.910000 465.000000 436.090000 ;
        RECT 460.000000 439.910000 465.000000 440.090000 ;
        RECT 460.000000 443.910000 465.000000 444.090000 ;
        RECT 460.000000 447.910000 465.000000 448.090000 ;
        RECT 460.000000 451.910000 465.000000 452.090000 ;
        RECT 510.000000 419.910000 515.000000 420.090000 ;
        RECT 510.000000 423.910000 515.000000 424.090000 ;
        RECT 510.000000 431.910000 515.000000 432.090000 ;
        RECT 510.000000 427.910000 515.000000 428.090000 ;
        RECT 510.000000 435.910000 515.000000 436.090000 ;
        RECT 510.000000 439.910000 515.000000 440.090000 ;
        RECT 510.000000 443.910000 515.000000 444.090000 ;
        RECT 510.000000 447.910000 515.000000 448.090000 ;
        RECT 510.000000 451.910000 515.000000 452.090000 ;
        RECT 460.000000 455.910000 465.000000 456.090000 ;
        RECT 460.000000 459.910000 465.000000 460.090000 ;
        RECT 460.000000 463.910000 465.000000 464.090000 ;
        RECT 460.000000 467.910000 465.000000 468.090000 ;
        RECT 460.000000 471.910000 465.000000 472.090000 ;
        RECT 460.000000 475.910000 465.000000 476.090000 ;
        RECT 460.000000 479.910000 465.000000 480.090000 ;
        RECT 460.000000 483.910000 465.000000 484.090000 ;
        RECT 460.000000 487.910000 465.000000 488.090000 ;
        RECT 510.000000 459.910000 515.000000 460.090000 ;
        RECT 510.000000 455.910000 515.000000 456.090000 ;
        RECT 510.000000 463.910000 515.000000 464.090000 ;
        RECT 510.000000 467.910000 515.000000 468.090000 ;
        RECT 510.000000 471.910000 515.000000 472.090000 ;
        RECT 510.000000 479.910000 515.000000 480.090000 ;
        RECT 510.000000 475.910000 515.000000 476.090000 ;
        RECT 510.000000 487.910000 515.000000 488.090000 ;
        RECT 510.000000 483.910000 515.000000 484.090000 ;
        RECT 560.000000 419.910000 565.000000 420.090000 ;
        RECT 560.000000 423.910000 565.000000 424.090000 ;
        RECT 560.000000 427.910000 565.000000 428.090000 ;
        RECT 560.000000 431.910000 565.000000 432.090000 ;
        RECT 560.000000 443.910000 565.000000 444.090000 ;
        RECT 560.000000 439.910000 565.000000 440.090000 ;
        RECT 560.000000 435.910000 565.000000 436.090000 ;
        RECT 560.000000 451.910000 565.000000 452.090000 ;
        RECT 560.000000 447.910000 565.000000 448.090000 ;
        RECT 560.000000 455.910000 565.000000 456.090000 ;
        RECT 560.000000 459.910000 565.000000 460.090000 ;
        RECT 560.000000 463.910000 565.000000 464.090000 ;
        RECT 560.000000 467.910000 565.000000 468.090000 ;
        RECT 560.000000 471.910000 565.000000 472.090000 ;
        RECT 560.000000 475.910000 565.000000 476.090000 ;
        RECT 560.000000 479.910000 565.000000 480.090000 ;
        RECT 560.000000 483.910000 565.000000 484.090000 ;
        RECT 560.000000 487.910000 565.000000 488.090000 ;
        RECT 360.000000 499.910000 371.000000 500.090000 ;
        RECT 360.000000 491.910000 371.000000 492.090000 ;
        RECT 360.000000 495.910000 371.000000 496.090000 ;
        RECT 360.000000 507.910000 371.000000 508.090000 ;
        RECT 360.000000 503.910000 371.000000 504.090000 ;
        RECT 360.000000 511.910000 371.000000 512.090000 ;
        RECT 360.000000 515.910000 371.000000 516.090000 ;
        RECT 360.000000 519.910000 371.000000 520.090000 ;
        RECT 360.000000 523.910000 371.000000 524.090000 ;
        RECT 360.000000 527.910000 371.000000 528.090000 ;
        RECT 360.000000 535.910000 371.000000 536.090000 ;
        RECT 360.000000 531.910000 371.000000 532.090000 ;
        RECT 360.000000 543.910000 371.000000 544.090000 ;
        RECT 360.000000 539.910000 371.000000 540.090000 ;
        RECT 360.000000 547.910000 371.000000 548.090000 ;
        RECT 360.000000 551.910000 371.000000 552.090000 ;
        RECT 360.000000 555.910000 371.000000 556.090000 ;
        RECT 360.000000 563.910000 371.000000 564.090000 ;
        RECT 360.000000 559.910000 371.000000 560.090000 ;
        RECT 310.000000 491.910000 315.000000 492.090000 ;
        RECT 310.000000 495.910000 315.000000 496.090000 ;
        RECT 310.000000 499.910000 315.000000 500.090000 ;
        RECT 310.000000 507.910000 315.000000 508.090000 ;
        RECT 310.000000 503.910000 315.000000 504.090000 ;
        RECT 310.000000 511.910000 315.000000 512.090000 ;
        RECT 310.000000 515.910000 315.000000 516.090000 ;
        RECT 410.000000 491.910000 415.000000 492.090000 ;
        RECT 410.000000 495.910000 415.000000 496.090000 ;
        RECT 410.000000 499.910000 415.000000 500.090000 ;
        RECT 410.000000 503.910000 415.000000 504.090000 ;
        RECT 360.000000 571.910000 371.000000 572.090000 ;
        RECT 360.000000 567.910000 371.000000 568.090000 ;
        RECT 360.000000 579.910000 371.000000 580.090000 ;
        RECT 360.000000 575.910000 371.000000 576.090000 ;
        RECT 360.000000 583.910000 371.000000 584.090000 ;
        RECT 360.000000 587.910000 371.000000 588.090000 ;
        RECT 360.000000 591.910000 371.000000 592.090000 ;
        RECT 360.000000 599.910000 371.000000 600.090000 ;
        RECT 360.000000 595.910000 371.000000 596.090000 ;
        RECT 360.000000 607.910000 371.000000 608.090000 ;
        RECT 360.000000 603.910000 371.000000 604.090000 ;
        RECT 360.000000 619.910000 371.000000 620.090000 ;
        RECT 360.000000 615.910000 371.000000 616.090000 ;
        RECT 360.000000 611.910000 371.000000 612.090000 ;
        RECT 360.000000 623.910000 371.000000 624.090000 ;
        RECT 360.000000 627.910000 371.000000 628.090000 ;
        RECT 360.000000 635.910000 371.000000 636.090000 ;
        RECT 360.000000 631.910000 371.000000 632.090000 ;
        RECT 460.000000 503.910000 465.000000 504.090000 ;
        RECT 460.000000 499.910000 465.000000 500.090000 ;
        RECT 460.000000 491.910000 465.000000 492.090000 ;
        RECT 460.000000 495.910000 465.000000 496.090000 ;
        RECT 510.000000 495.910000 515.000000 496.090000 ;
        RECT 510.000000 491.910000 515.000000 492.090000 ;
        RECT 510.000000 499.910000 515.000000 500.090000 ;
        RECT 510.000000 503.910000 515.000000 504.090000 ;
        RECT 560.000000 499.910000 565.000000 500.090000 ;
        RECT 560.000000 495.910000 565.000000 496.090000 ;
        RECT 560.000000 491.910000 565.000000 492.090000 ;
        RECT 560.000000 503.910000 565.000000 504.090000 ;
        RECT 360.000000 639.910000 371.000000 640.090000 ;
        RECT 360.000000 643.910000 371.000000 644.090000 ;
        RECT 360.000000 647.910000 371.000000 648.090000 ;
        RECT 360.000000 655.910000 371.000000 656.090000 ;
        RECT 360.000000 651.910000 371.000000 652.090000 ;
        RECT 360.000000 667.910000 371.000000 668.090000 ;
        RECT 360.000000 663.910000 371.000000 664.090000 ;
        RECT 360.000000 659.910000 371.000000 660.090000 ;
        RECT 360.000000 675.910000 365.000000 676.090000 ;
        RECT 360.000000 671.910000 365.000000 672.090000 ;
        RECT 310.000000 679.910000 315.000000 680.090000 ;
        RECT 310.000000 683.910000 315.000000 684.090000 ;
        RECT 360.000000 679.910000 365.000000 680.090000 ;
        RECT 360.000000 683.910000 365.000000 684.090000 ;
        RECT 410.000000 659.910000 415.000000 660.090000 ;
        RECT 410.000000 663.910000 415.000000 664.090000 ;
        RECT 410.000000 667.910000 415.000000 668.090000 ;
        RECT 410.000000 671.910000 415.000000 672.090000 ;
        RECT 410.000000 675.910000 415.000000 676.090000 ;
        RECT 410.000000 683.910000 415.000000 684.090000 ;
        RECT 410.000000 679.910000 415.000000 680.090000 ;
        RECT 460.000000 659.910000 465.000000 660.090000 ;
        RECT 460.000000 663.910000 465.000000 664.090000 ;
        RECT 460.000000 667.910000 465.000000 668.090000 ;
        RECT 460.000000 671.910000 465.000000 672.090000 ;
        RECT 460.000000 675.910000 465.000000 676.090000 ;
        RECT 510.000000 663.910000 515.000000 664.090000 ;
        RECT 510.000000 659.910000 515.000000 660.090000 ;
        RECT 510.000000 667.910000 515.000000 668.090000 ;
        RECT 510.000000 671.910000 515.000000 672.090000 ;
        RECT 510.000000 675.910000 515.000000 676.090000 ;
        RECT 460.000000 683.910000 465.000000 684.090000 ;
        RECT 460.000000 679.910000 465.000000 680.090000 ;
        RECT 510.000000 683.910000 515.000000 684.090000 ;
        RECT 510.000000 679.910000 515.000000 680.090000 ;
        RECT 560.000000 659.910000 565.000000 660.090000 ;
        RECT 560.000000 663.910000 565.000000 664.090000 ;
        RECT 560.000000 667.910000 565.000000 668.090000 ;
        RECT 560.000000 671.910000 565.000000 672.090000 ;
        RECT 560.000000 675.910000 565.000000 676.090000 ;
        RECT 560.000000 683.910000 565.000000 684.090000 ;
        RECT 560.000000 679.910000 565.000000 680.090000 ;
        RECT 610.000000 379.910000 615.000000 380.090000 ;
        RECT 660.000000 379.910000 665.000000 380.090000 ;
        RECT 610.000000 343.910000 615.000000 344.090000 ;
        RECT 610.000000 347.910000 615.000000 348.090000 ;
        RECT 610.000000 351.910000 615.000000 352.090000 ;
        RECT 610.000000 355.910000 615.000000 356.090000 ;
        RECT 610.000000 359.910000 615.000000 360.090000 ;
        RECT 610.000000 363.910000 615.000000 364.090000 ;
        RECT 610.000000 367.910000 615.000000 368.090000 ;
        RECT 610.000000 371.910000 615.000000 372.090000 ;
        RECT 610.000000 375.910000 615.000000 376.090000 ;
        RECT 660.000000 343.910000 665.000000 344.090000 ;
        RECT 660.000000 351.910000 665.000000 352.090000 ;
        RECT 660.000000 347.910000 665.000000 348.090000 ;
        RECT 660.000000 355.910000 665.000000 356.090000 ;
        RECT 660.000000 359.910000 665.000000 360.090000 ;
        RECT 660.000000 363.910000 665.000000 364.090000 ;
        RECT 660.000000 367.910000 665.000000 368.090000 ;
        RECT 660.000000 371.910000 665.000000 372.090000 ;
        RECT 660.000000 375.910000 665.000000 376.090000 ;
        RECT 610.000000 395.910000 615.000000 396.090000 ;
        RECT 610.000000 391.910000 615.000000 392.090000 ;
        RECT 610.000000 387.910000 615.000000 388.090000 ;
        RECT 610.000000 383.910000 615.000000 384.090000 ;
        RECT 610.000000 399.910000 615.000000 400.090000 ;
        RECT 610.000000 403.910000 615.000000 404.090000 ;
        RECT 610.000000 407.910000 615.000000 408.090000 ;
        RECT 610.000000 411.910000 615.000000 412.090000 ;
        RECT 610.000000 415.910000 615.000000 416.090000 ;
        RECT 660.000000 383.910000 665.000000 384.090000 ;
        RECT 660.000000 387.910000 665.000000 388.090000 ;
        RECT 660.000000 391.910000 665.000000 392.090000 ;
        RECT 660.000000 395.910000 665.000000 396.090000 ;
        RECT 660.000000 403.910000 665.000000 404.090000 ;
        RECT 660.000000 399.910000 665.000000 400.090000 ;
        RECT 660.000000 407.910000 665.000000 408.090000 ;
        RECT 660.000000 411.910000 665.000000 412.090000 ;
        RECT 660.000000 415.910000 665.000000 416.090000 ;
        RECT 710.000000 379.910000 715.000000 380.090000 ;
        RECT 710.000000 343.910000 715.000000 344.090000 ;
        RECT 710.000000 347.910000 715.000000 348.090000 ;
        RECT 710.000000 351.910000 715.000000 352.090000 ;
        RECT 710.000000 355.910000 715.000000 356.090000 ;
        RECT 710.000000 359.910000 715.000000 360.090000 ;
        RECT 710.000000 367.910000 715.000000 368.090000 ;
        RECT 710.000000 363.910000 715.000000 364.090000 ;
        RECT 710.000000 375.910000 715.000000 376.090000 ;
        RECT 710.000000 371.910000 715.000000 372.090000 ;
        RECT 710.000000 383.910000 715.000000 384.090000 ;
        RECT 710.000000 387.910000 715.000000 388.090000 ;
        RECT 710.000000 391.910000 715.000000 392.090000 ;
        RECT 710.000000 395.910000 715.000000 396.090000 ;
        RECT 710.000000 403.910000 715.000000 404.090000 ;
        RECT 710.000000 399.910000 715.000000 400.090000 ;
        RECT 713.500000 415.910000 718.500000 416.090000 ;
        RECT 710.000000 411.910000 718.500000 412.090000 ;
        RECT 710.000000 407.910000 715.000000 408.090000 ;
        RECT 610.000000 431.910000 615.000000 432.090000 ;
        RECT 610.000000 427.910000 615.000000 428.090000 ;
        RECT 610.000000 423.910000 615.000000 424.090000 ;
        RECT 610.000000 419.910000 615.000000 420.090000 ;
        RECT 610.000000 435.910000 615.000000 436.090000 ;
        RECT 610.000000 439.910000 615.000000 440.090000 ;
        RECT 610.000000 443.910000 615.000000 444.090000 ;
        RECT 610.000000 447.910000 615.000000 448.090000 ;
        RECT 610.000000 451.910000 615.000000 452.090000 ;
        RECT 660.000000 419.910000 665.000000 420.090000 ;
        RECT 660.000000 423.910000 665.000000 424.090000 ;
        RECT 660.000000 427.910000 665.000000 428.090000 ;
        RECT 660.000000 431.910000 665.000000 432.090000 ;
        RECT 660.000000 439.910000 665.000000 440.090000 ;
        RECT 660.000000 435.910000 665.000000 436.090000 ;
        RECT 660.000000 443.910000 665.000000 444.090000 ;
        RECT 660.000000 447.910000 665.000000 448.090000 ;
        RECT 660.000000 451.910000 665.000000 452.090000 ;
        RECT 610.000000 455.910000 615.000000 456.090000 ;
        RECT 610.000000 459.910000 615.000000 460.090000 ;
        RECT 610.000000 463.910000 615.000000 464.090000 ;
        RECT 610.000000 467.910000 615.000000 468.090000 ;
        RECT 610.000000 471.910000 615.000000 472.090000 ;
        RECT 610.000000 475.910000 615.000000 476.090000 ;
        RECT 610.000000 479.910000 615.000000 480.090000 ;
        RECT 610.000000 483.910000 615.000000 484.090000 ;
        RECT 610.000000 487.910000 615.000000 488.090000 ;
        RECT 660.000000 459.910000 665.000000 460.090000 ;
        RECT 660.000000 455.910000 665.000000 456.090000 ;
        RECT 660.000000 463.910000 665.000000 464.090000 ;
        RECT 660.000000 467.910000 665.000000 468.090000 ;
        RECT 660.000000 471.910000 665.000000 472.090000 ;
        RECT 660.000000 479.910000 665.000000 480.090000 ;
        RECT 660.000000 475.910000 665.000000 476.090000 ;
        RECT 660.000000 487.910000 665.000000 488.090000 ;
        RECT 660.000000 483.910000 665.000000 484.090000 ;
        RECT 711.000000 423.910000 721.000000 424.090000 ;
        RECT 711.000000 419.910000 721.000000 420.090000 ;
        RECT 710.000000 431.910000 721.000000 432.090000 ;
        RECT 711.000000 427.910000 721.000000 428.090000 ;
        RECT 710.000000 435.910000 721.000000 436.090000 ;
        RECT 710.000000 439.910000 721.000000 440.090000 ;
        RECT 710.000000 443.910000 721.000000 444.090000 ;
        RECT 710.000000 451.910000 721.000000 452.090000 ;
        RECT 710.000000 447.910000 721.000000 448.090000 ;
        RECT 710.000000 455.910000 721.000000 456.090000 ;
        RECT 710.000000 459.910000 721.000000 460.090000 ;
        RECT 710.000000 471.910000 721.000000 472.090000 ;
        RECT 710.000000 463.910000 721.000000 464.090000 ;
        RECT 710.000000 467.910000 721.000000 468.090000 ;
        RECT 710.000000 475.910000 721.000000 476.090000 ;
        RECT 710.000000 479.910000 721.000000 480.090000 ;
        RECT 710.000000 483.910000 721.000000 484.090000 ;
        RECT 710.000000 487.910000 721.000000 488.090000 ;
        RECT 810.000000 379.910000 815.000000 380.090000 ;
        RECT 760.000000 379.910000 765.000000 380.090000 ;
        RECT 760.000000 343.910000 765.000000 344.090000 ;
        RECT 760.000000 347.910000 765.000000 348.090000 ;
        RECT 760.000000 351.910000 765.000000 352.090000 ;
        RECT 760.000000 355.910000 765.000000 356.090000 ;
        RECT 760.000000 359.910000 765.000000 360.090000 ;
        RECT 760.000000 363.910000 765.000000 364.090000 ;
        RECT 760.000000 367.910000 765.000000 368.090000 ;
        RECT 760.000000 375.910000 765.000000 376.090000 ;
        RECT 760.000000 371.910000 765.000000 372.090000 ;
        RECT 810.000000 343.910000 815.000000 344.090000 ;
        RECT 810.000000 347.910000 815.000000 348.090000 ;
        RECT 810.000000 351.910000 815.000000 352.090000 ;
        RECT 810.000000 359.910000 815.000000 360.090000 ;
        RECT 810.000000 355.910000 815.000000 356.090000 ;
        RECT 810.000000 363.910000 815.000000 364.090000 ;
        RECT 810.000000 367.910000 815.000000 368.090000 ;
        RECT 810.000000 371.910000 815.000000 372.090000 ;
        RECT 810.000000 375.910000 815.000000 376.090000 ;
        RECT 760.000000 395.910000 765.000000 396.090000 ;
        RECT 760.000000 391.910000 765.000000 392.090000 ;
        RECT 760.000000 387.910000 765.000000 388.090000 ;
        RECT 760.000000 383.910000 765.000000 384.090000 ;
        RECT 760.000000 399.910000 765.000000 400.090000 ;
        RECT 760.000000 403.910000 765.000000 404.090000 ;
        RECT 760.000000 407.910000 765.000000 408.090000 ;
        RECT 760.000000 411.910000 765.000000 412.090000 ;
        RECT 760.000000 415.910000 765.000000 416.090000 ;
        RECT 810.000000 387.910000 815.000000 388.090000 ;
        RECT 810.000000 383.910000 815.000000 384.090000 ;
        RECT 810.000000 391.910000 815.000000 392.090000 ;
        RECT 810.000000 395.910000 815.000000 396.090000 ;
        RECT 810.000000 403.910000 815.000000 404.090000 ;
        RECT 810.000000 399.910000 815.000000 400.090000 ;
        RECT 810.000000 407.910000 815.000000 408.090000 ;
        RECT 810.000000 411.910000 815.000000 412.090000 ;
        RECT 810.000000 415.910000 815.000000 416.090000 ;
        RECT 860.000000 379.910000 865.000000 380.090000 ;
        RECT 860.000000 359.910000 865.000000 360.090000 ;
        RECT 860.000000 355.910000 865.000000 356.090000 ;
        RECT 860.000000 351.910000 865.000000 352.090000 ;
        RECT 860.000000 347.910000 865.000000 348.090000 ;
        RECT 860.000000 343.910000 865.000000 344.090000 ;
        RECT 860.000000 363.910000 865.000000 364.090000 ;
        RECT 860.000000 367.910000 865.000000 368.090000 ;
        RECT 860.000000 371.910000 865.000000 372.090000 ;
        RECT 860.000000 375.910000 865.000000 376.090000 ;
        RECT 860.000000 383.910000 865.000000 384.090000 ;
        RECT 860.000000 387.910000 865.000000 388.090000 ;
        RECT 860.000000 391.910000 865.000000 392.090000 ;
        RECT 860.000000 395.910000 865.000000 396.090000 ;
        RECT 860.000000 403.910000 865.000000 404.090000 ;
        RECT 860.000000 399.910000 865.000000 400.090000 ;
        RECT 860.000000 415.910000 865.000000 416.090000 ;
        RECT 860.000000 411.910000 865.000000 412.090000 ;
        RECT 860.000000 407.910000 865.000000 408.090000 ;
        RECT 760.000000 419.910000 765.000000 420.090000 ;
        RECT 760.000000 423.910000 765.000000 424.090000 ;
        RECT 760.000000 427.910000 765.000000 428.090000 ;
        RECT 760.000000 431.910000 765.000000 432.090000 ;
        RECT 760.000000 435.910000 765.000000 436.090000 ;
        RECT 760.000000 439.910000 765.000000 440.090000 ;
        RECT 760.000000 443.910000 765.000000 444.090000 ;
        RECT 810.000000 419.910000 815.000000 420.090000 ;
        RECT 810.000000 423.910000 815.000000 424.090000 ;
        RECT 810.000000 431.910000 815.000000 432.090000 ;
        RECT 810.000000 427.910000 815.000000 428.090000 ;
        RECT 810.000000 435.910000 815.000000 436.090000 ;
        RECT 810.000000 439.910000 815.000000 440.090000 ;
        RECT 810.000000 443.910000 815.000000 444.090000 ;
        RECT 860.000000 419.910000 865.000000 420.090000 ;
        RECT 860.000000 423.910000 865.000000 424.090000 ;
        RECT 860.000000 427.910000 865.000000 428.090000 ;
        RECT 860.000000 431.910000 865.000000 432.090000 ;
        RECT 860.000000 443.910000 865.000000 444.090000 ;
        RECT 860.000000 439.910000 865.000000 440.090000 ;
        RECT 860.000000 435.910000 865.000000 436.090000 ;
        RECT 610.000000 491.910000 615.000000 492.090000 ;
        RECT 610.000000 499.910000 615.000000 500.090000 ;
        RECT 610.000000 495.910000 615.000000 496.090000 ;
        RECT 610.000000 503.910000 615.000000 504.090000 ;
        RECT 660.000000 495.910000 665.000000 496.090000 ;
        RECT 660.000000 491.910000 665.000000 492.090000 ;
        RECT 660.000000 499.910000 665.000000 500.090000 ;
        RECT 660.000000 503.910000 665.000000 504.090000 ;
        RECT 710.000000 503.910000 715.000000 504.090000 ;
        RECT 710.000000 499.910000 715.000000 500.090000 ;
        RECT 710.000000 495.910000 715.000000 496.090000 ;
        RECT 710.000000 491.910000 715.000000 492.090000 ;
        RECT 960.000000 379.910000 965.000000 380.090000 ;
        RECT 960.000000 343.910000 965.000000 344.090000 ;
        RECT 960.000000 347.910000 965.000000 348.090000 ;
        RECT 960.000000 351.910000 965.000000 352.090000 ;
        RECT 960.000000 355.910000 965.000000 356.090000 ;
        RECT 960.000000 359.910000 965.000000 360.090000 ;
        RECT 960.000000 375.910000 965.000000 376.090000 ;
        RECT 960.000000 371.910000 965.000000 372.090000 ;
        RECT 960.000000 367.910000 965.000000 368.090000 ;
        RECT 960.000000 363.910000 965.000000 364.090000 ;
        RECT 960.000000 383.910000 965.000000 384.090000 ;
        RECT 960.000000 387.910000 965.000000 388.090000 ;
        RECT 960.000000 391.910000 965.000000 392.090000 ;
        RECT 960.000000 395.910000 965.000000 396.090000 ;
        RECT 960.000000 399.910000 965.000000 400.090000 ;
        RECT 960.000000 403.910000 965.000000 404.090000 ;
        RECT 960.000000 407.910000 965.000000 408.090000 ;
        RECT 960.000000 411.910000 965.000000 412.090000 ;
        RECT 960.000000 415.910000 965.000000 416.090000 ;
        RECT 910.000000 379.910000 915.000000 380.090000 ;
        RECT 910.000000 343.910000 915.000000 344.090000 ;
        RECT 910.000000 347.910000 915.000000 348.090000 ;
        RECT 910.000000 351.910000 915.000000 352.090000 ;
        RECT 910.000000 355.910000 915.000000 356.090000 ;
        RECT 910.000000 359.910000 915.000000 360.090000 ;
        RECT 910.000000 363.910000 915.000000 364.090000 ;
        RECT 910.000000 367.910000 915.000000 368.090000 ;
        RECT 910.000000 371.910000 915.000000 372.090000 ;
        RECT 910.000000 375.910000 915.000000 376.090000 ;
        RECT 910.000000 395.910000 915.000000 396.090000 ;
        RECT 910.000000 391.910000 915.000000 392.090000 ;
        RECT 910.000000 387.910000 915.000000 388.090000 ;
        RECT 910.000000 383.910000 915.000000 384.090000 ;
        RECT 910.000000 399.910000 915.000000 400.090000 ;
        RECT 910.000000 403.910000 915.000000 404.090000 ;
        RECT 910.000000 407.910000 915.000000 408.090000 ;
        RECT 910.000000 411.910000 915.000000 412.090000 ;
        RECT 910.000000 415.910000 915.000000 416.090000 ;
        RECT 1010.000000 379.910000 1015.000000 380.090000 ;
        RECT 1010.000000 343.910000 1015.000000 344.090000 ;
        RECT 1010.000000 347.910000 1015.000000 348.090000 ;
        RECT 1010.000000 351.910000 1015.000000 352.090000 ;
        RECT 1010.000000 359.910000 1015.000000 360.090000 ;
        RECT 1010.000000 355.910000 1015.000000 356.090000 ;
        RECT 1010.000000 363.910000 1015.000000 364.090000 ;
        RECT 1010.000000 367.910000 1015.000000 368.090000 ;
        RECT 1010.000000 371.910000 1015.000000 372.090000 ;
        RECT 1010.000000 375.910000 1015.000000 376.090000 ;
        RECT 1010.000000 387.910000 1015.000000 388.090000 ;
        RECT 1010.000000 383.910000 1015.000000 384.090000 ;
        RECT 1010.000000 391.910000 1015.000000 392.090000 ;
        RECT 1010.000000 395.910000 1015.000000 396.090000 ;
        RECT 1010.000000 399.910000 1015.000000 400.090000 ;
        RECT 1010.000000 403.910000 1015.000000 404.090000 ;
        RECT 1010.000000 407.910000 1015.000000 408.090000 ;
        RECT 1010.000000 411.910000 1015.000000 412.090000 ;
        RECT 1010.000000 415.910000 1015.000000 416.090000 ;
        RECT 960.000000 431.910000 965.000000 432.090000 ;
        RECT 960.000000 427.910000 965.000000 428.090000 ;
        RECT 960.000000 423.910000 965.000000 424.090000 ;
        RECT 960.000000 419.910000 965.000000 420.090000 ;
        RECT 960.000000 443.910000 965.000000 444.090000 ;
        RECT 960.000000 439.910000 965.000000 440.090000 ;
        RECT 960.000000 435.910000 965.000000 436.090000 ;
        RECT 910.000000 431.910000 915.000000 432.090000 ;
        RECT 910.000000 427.910000 915.000000 428.090000 ;
        RECT 910.000000 423.910000 915.000000 424.090000 ;
        RECT 910.000000 419.910000 915.000000 420.090000 ;
        RECT 910.000000 435.910000 915.000000 436.090000 ;
        RECT 910.000000 439.910000 915.000000 440.090000 ;
        RECT 910.000000 443.910000 915.000000 444.090000 ;
        RECT 1010.000000 419.910000 1015.000000 420.090000 ;
        RECT 1010.000000 423.910000 1015.000000 424.090000 ;
        RECT 1010.000000 427.910000 1015.000000 428.090000 ;
        RECT 1010.000000 431.910000 1015.000000 432.090000 ;
        RECT 1010.000000 435.910000 1015.000000 436.090000 ;
        RECT 1010.000000 439.910000 1015.000000 440.090000 ;
        RECT 1010.000000 443.910000 1015.000000 444.090000 ;
        RECT 1110.000000 379.910000 1115.000000 380.090000 ;
        RECT 1110.000000 343.910000 1115.000000 344.090000 ;
        RECT 1110.000000 347.910000 1115.000000 348.090000 ;
        RECT 1110.000000 351.910000 1115.000000 352.090000 ;
        RECT 1110.000000 355.910000 1115.000000 356.090000 ;
        RECT 1110.000000 359.910000 1115.000000 360.090000 ;
        RECT 1110.000000 375.910000 1115.000000 376.090000 ;
        RECT 1110.000000 371.910000 1115.000000 372.090000 ;
        RECT 1110.000000 367.910000 1115.000000 368.090000 ;
        RECT 1110.000000 363.910000 1115.000000 364.090000 ;
        RECT 1110.000000 383.910000 1115.000000 384.090000 ;
        RECT 1110.000000 387.910000 1115.000000 388.090000 ;
        RECT 1110.000000 391.910000 1115.000000 392.090000 ;
        RECT 1110.000000 395.910000 1115.000000 396.090000 ;
        RECT 1110.000000 399.910000 1115.000000 400.090000 ;
        RECT 1110.000000 403.910000 1115.000000 404.090000 ;
        RECT 1110.000000 407.910000 1115.000000 408.090000 ;
        RECT 1110.000000 411.910000 1115.000000 412.090000 ;
        RECT 1110.000000 415.910000 1115.000000 416.090000 ;
        RECT 1060.000000 379.910000 1065.000000 380.090000 ;
        RECT 1060.000000 343.910000 1065.000000 344.090000 ;
        RECT 1060.000000 347.910000 1065.000000 348.090000 ;
        RECT 1060.000000 351.910000 1065.000000 352.090000 ;
        RECT 1060.000000 355.910000 1065.000000 356.090000 ;
        RECT 1060.000000 359.910000 1065.000000 360.090000 ;
        RECT 1060.000000 375.910000 1065.000000 376.090000 ;
        RECT 1060.000000 371.910000 1065.000000 372.090000 ;
        RECT 1060.000000 367.910000 1065.000000 368.090000 ;
        RECT 1060.000000 363.910000 1065.000000 364.090000 ;
        RECT 1060.000000 395.910000 1065.000000 396.090000 ;
        RECT 1060.000000 391.910000 1065.000000 392.090000 ;
        RECT 1060.000000 387.910000 1065.000000 388.090000 ;
        RECT 1060.000000 383.910000 1065.000000 384.090000 ;
        RECT 1060.000000 399.910000 1065.000000 400.090000 ;
        RECT 1060.000000 403.910000 1065.000000 404.090000 ;
        RECT 1060.000000 407.910000 1065.000000 408.090000 ;
        RECT 1060.000000 411.910000 1065.000000 412.090000 ;
        RECT 1060.000000 415.910000 1065.000000 416.090000 ;
        RECT 1158.000000 379.910000 1168.000000 380.090000 ;
        RECT 1158.000000 343.910000 1168.000000 344.090000 ;
        RECT 1158.000000 347.910000 1168.000000 348.090000 ;
        RECT 1158.000000 351.910000 1168.000000 352.090000 ;
        RECT 1158.000000 355.910000 1168.000000 356.090000 ;
        RECT 1158.000000 359.910000 1168.000000 360.090000 ;
        RECT 1158.000000 375.910000 1168.000000 376.090000 ;
        RECT 1158.000000 371.910000 1168.000000 372.090000 ;
        RECT 1158.000000 367.910000 1168.000000 368.090000 ;
        RECT 1158.000000 363.910000 1168.000000 364.090000 ;
        RECT 1158.000000 395.910000 1168.000000 396.090000 ;
        RECT 1158.000000 391.910000 1168.000000 392.090000 ;
        RECT 1158.000000 387.910000 1168.000000 388.090000 ;
        RECT 1158.000000 383.910000 1168.000000 384.090000 ;
        RECT 1158.000000 399.910000 1168.000000 400.090000 ;
        RECT 1158.000000 403.910000 1168.000000 404.090000 ;
        RECT 1158.000000 407.910000 1168.000000 408.090000 ;
        RECT 1158.000000 411.910000 1168.000000 412.090000 ;
        RECT 1158.000000 415.910000 1168.000000 416.090000 ;
        RECT 1110.000000 431.910000 1115.000000 432.090000 ;
        RECT 1110.000000 427.910000 1115.000000 428.090000 ;
        RECT 1110.000000 423.910000 1115.000000 424.090000 ;
        RECT 1110.000000 419.910000 1115.000000 420.090000 ;
        RECT 1110.000000 443.910000 1115.000000 444.090000 ;
        RECT 1110.000000 439.910000 1115.000000 440.090000 ;
        RECT 1110.000000 435.910000 1115.000000 436.090000 ;
        RECT 1060.000000 419.910000 1065.000000 420.090000 ;
        RECT 1060.000000 423.910000 1065.000000 424.090000 ;
        RECT 1060.000000 427.910000 1065.000000 428.090000 ;
        RECT 1060.000000 431.910000 1065.000000 432.090000 ;
        RECT 1060.000000 435.910000 1065.000000 436.090000 ;
        RECT 1060.000000 439.910000 1065.000000 440.090000 ;
        RECT 1060.000000 443.910000 1065.000000 444.090000 ;
        RECT 1158.000000 427.910000 1168.000000 428.090000 ;
        RECT 1158.000000 423.910000 1168.000000 424.090000 ;
        RECT 1158.000000 419.910000 1168.000000 420.090000 ;
        RECT 1160.000000 431.910000 1165.000000 432.090000 ;
        RECT 1160.000000 435.910000 1165.000000 436.090000 ;
        RECT 1160.000000 439.910000 1165.000000 440.090000 ;
        RECT 1160.000000 443.910000 1165.000000 444.090000 ;
        RECT 1160.000000 447.910000 1165.000000 448.090000 ;
        RECT 1160.000000 451.910000 1165.000000 452.090000 ;
        RECT 1160.000000 459.910000 1165.000000 460.090000 ;
        RECT 1160.000000 455.910000 1165.000000 456.090000 ;
        RECT 1160.000000 463.910000 1165.000000 464.090000 ;
        RECT 1160.000000 467.910000 1165.000000 468.090000 ;
        RECT 1160.000000 471.910000 1165.000000 472.090000 ;
        RECT 1160.000000 479.910000 1165.000000 480.090000 ;
        RECT 1160.000000 475.910000 1165.000000 476.090000 ;
        RECT 1160.000000 487.910000 1165.000000 488.090000 ;
        RECT 1160.000000 483.910000 1165.000000 484.090000 ;
        RECT 1160.000000 491.910000 1165.000000 492.090000 ;
        RECT 1160.000000 495.910000 1165.000000 496.090000 ;
        RECT 1160.000000 499.910000 1165.000000 500.090000 ;
        RECT 1160.000000 507.910000 1165.000000 508.090000 ;
        RECT 1160.000000 503.910000 1165.000000 504.090000 ;
        RECT 1160.000000 511.910000 1165.000000 512.090000 ;
        RECT 1160.000000 515.910000 1165.000000 516.090000 ;
        RECT 1160.000000 519.910000 1165.000000 520.090000 ;
        RECT 1160.000000 523.910000 1165.000000 524.090000 ;
        RECT 1160.000000 527.910000 1165.000000 528.090000 ;
        RECT 1160.000000 535.910000 1165.000000 536.090000 ;
        RECT 1160.000000 531.910000 1165.000000 532.090000 ;
        RECT 1160.000000 539.910000 1165.000000 540.090000 ;
        RECT 1160.000000 543.910000 1165.000000 544.090000 ;
        RECT 1160.000000 547.910000 1165.000000 548.090000 ;
        RECT 1160.000000 551.910000 1165.000000 552.090000 ;
        RECT 1160.000000 555.910000 1165.000000 556.090000 ;
        RECT 1160.000000 563.910000 1165.000000 564.090000 ;
        RECT 1160.000000 559.910000 1165.000000 560.090000 ;
        RECT 1160.000000 567.910000 1165.000000 568.090000 ;
        RECT 1160.000000 571.910000 1165.000000 572.090000 ;
        RECT 1160.000000 579.910000 1165.000000 580.090000 ;
        RECT 1160.000000 575.910000 1165.000000 576.090000 ;
        RECT 1160.000000 583.910000 1165.000000 584.090000 ;
        RECT 1160.000000 587.910000 1165.000000 588.090000 ;
        RECT 1160.000000 591.910000 1165.000000 592.090000 ;
        RECT 1160.000000 595.910000 1165.000000 596.090000 ;
        RECT 1160.000000 599.910000 1165.000000 600.090000 ;
        RECT 1160.000000 607.910000 1165.000000 608.090000 ;
        RECT 1160.000000 603.910000 1165.000000 604.090000 ;
        RECT 1160.000000 611.910000 1165.000000 612.090000 ;
        RECT 1160.000000 615.910000 1165.000000 616.090000 ;
        RECT 1160.000000 619.910000 1165.000000 620.090000 ;
        RECT 1160.000000 623.910000 1165.000000 624.090000 ;
        RECT 1160.000000 627.910000 1165.000000 628.090000 ;
        RECT 1160.000000 635.910000 1165.000000 636.090000 ;
        RECT 1160.000000 631.910000 1165.000000 632.090000 ;
        RECT 610.000000 659.910000 615.000000 660.090000 ;
        RECT 610.000000 663.910000 615.000000 664.090000 ;
        RECT 610.000000 667.910000 615.000000 668.090000 ;
        RECT 610.000000 671.910000 615.000000 672.090000 ;
        RECT 610.000000 675.910000 615.000000 676.090000 ;
        RECT 660.000000 663.910000 665.000000 664.090000 ;
        RECT 660.000000 659.910000 665.000000 660.090000 ;
        RECT 660.000000 667.910000 665.000000 668.090000 ;
        RECT 660.000000 671.910000 665.000000 672.090000 ;
        RECT 660.000000 675.910000 665.000000 676.090000 ;
        RECT 610.000000 683.910000 615.000000 684.090000 ;
        RECT 610.000000 679.910000 615.000000 680.090000 ;
        RECT 660.000000 683.910000 665.000000 684.090000 ;
        RECT 660.000000 679.910000 665.000000 680.090000 ;
        RECT 1160.000000 639.910000 1165.000000 640.090000 ;
        RECT 1160.000000 643.910000 1165.000000 644.090000 ;
        RECT 1160.000000 647.910000 1165.000000 648.090000 ;
        RECT 1160.000000 655.910000 1165.000000 656.090000 ;
        RECT 1160.000000 651.910000 1165.000000 652.090000 ;
        RECT 1160.000000 663.910000 1165.000000 664.090000 ;
        RECT 1160.000000 659.910000 1165.000000 660.090000 ;
        RECT 1160.000000 667.910000 1165.000000 668.090000 ;
        RECT 1160.000000 671.910000 1165.000000 672.090000 ;
        RECT 1160.000000 675.910000 1165.000000 676.090000 ;
        RECT 1160.000000 683.910000 1165.000000 684.090000 ;
        RECT 1160.000000 679.910000 1165.000000 680.090000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  OBS
    LAYER OVERLAP ;
      RECT 0.000000 656.000000 670.000000 686.000000 ;
      RECT 0.000000 506.000000 389.000000 656.000000 ;
      RECT 1139.000000 446.000000 1186.000000 686.000000 ;
      RECT 0.000000 446.000000 739.000000 506.000000 ;
      RECT 0.000000 0.000000 1186.000000 446.000000 ;
    LAYER M1 ;
      RECT 0.000000 656.000000 670.000000 686.000000 ;
      RECT 0.000000 506.000000 389.000000 656.000000 ;
      RECT 1139.000000 446.000000 1186.000000 686.000000 ;
      RECT 0.000000 446.000000 739.000000 506.000000 ;
      RECT 0.000000 0.000000 1186.000000 446.000000 ;
    LAYER M2 ;
      RECT 1139.000000 685.590000 1186.000000 686.000000 ;
      RECT 647.765000 685.590000 670.000000 686.000000 ;
      RECT 561.965000 685.590000 624.430000 686.000000 ;
      RECT 556.285000 685.590000 558.865000 686.000000 ;
      RECT 476.165000 685.590000 538.630000 686.000000 ;
      RECT 455.930000 685.590000 463.425000 686.000000 ;
      RECT 390.365000 685.590000 452.830000 686.000000 ;
      RECT 304.565000 685.590000 367.030000 686.000000 ;
      RECT 647.765000 683.980000 658.500000 685.590000 ;
      RECT 642.085000 683.980000 644.665000 686.000000 ;
      RECT 638.125000 683.980000 638.985000 686.000000 ;
      RECT 627.530000 683.980000 635.025000 686.000000 ;
      RECT 616.500000 683.980000 624.430000 685.590000 ;
      RECT 556.285000 683.980000 558.500000 685.590000 ;
      RECT 552.325000 683.980000 553.185000 686.000000 ;
      RECT 541.730000 683.980000 549.225000 686.000000 ;
      RECT 516.500000 683.980000 538.630000 685.590000 ;
      RECT 476.165000 683.980000 508.500000 685.590000 ;
      RECT 470.485000 683.980000 473.065000 686.000000 ;
      RECT 466.525000 683.980000 467.385000 686.000000 ;
      RECT 455.930000 683.980000 458.500000 685.590000 ;
      RECT 416.500000 683.980000 452.830000 685.590000 ;
      RECT 390.365000 683.980000 408.500000 685.590000 ;
      RECT 384.685000 683.980000 387.265000 686.000000 ;
      RECT 380.725000 683.980000 381.585000 686.000000 ;
      RECT 370.130000 683.980000 377.625000 686.000000 ;
      RECT 366.500000 683.980000 367.030000 685.590000 ;
      RECT 304.565000 683.980000 308.500000 685.590000 ;
      RECT 298.885000 683.980000 301.465000 686.000000 ;
      RECT 294.925000 683.980000 295.785000 686.000000 ;
      RECT 284.330000 683.980000 291.825000 686.000000 ;
      RECT 218.765000 683.980000 281.230000 686.000000 ;
      RECT 213.085000 683.980000 215.665000 686.000000 ;
      RECT 209.125000 683.980000 209.985000 686.000000 ;
      RECT 198.530000 683.980000 206.025000 686.000000 ;
      RECT 132.965000 683.980000 195.430000 686.000000 ;
      RECT 127.285000 683.980000 129.865000 686.000000 ;
      RECT 123.325000 683.980000 124.185000 686.000000 ;
      RECT 112.730000 683.980000 120.225000 686.000000 ;
      RECT 47.165000 683.980000 109.630000 686.000000 ;
      RECT 41.485000 683.980000 44.065000 686.000000 ;
      RECT 37.525000 683.980000 38.385000 686.000000 ;
      RECT 26.930000 683.980000 34.425000 686.000000 ;
      RECT 0.000000 683.980000 23.830000 686.000000 ;
      RECT 1139.000000 683.590000 1158.500000 685.590000 ;
      RECT 616.500000 683.590000 658.500000 683.980000 ;
      RECT 566.500000 683.590000 608.500000 685.590000 ;
      RECT 516.500000 683.590000 558.500000 683.980000 ;
      RECT 466.500000 683.590000 508.500000 683.980000 ;
      RECT 416.500000 683.590000 458.500000 683.980000 ;
      RECT 366.500000 683.590000 408.500000 683.980000 ;
      RECT 316.500000 683.590000 358.500000 685.590000 ;
      RECT 0.000000 683.590000 308.500000 683.980000 ;
      RECT 1166.500000 682.410000 1186.000000 685.590000 ;
      RECT 1157.500000 682.410000 1158.500000 683.590000 ;
      RECT 666.500000 682.410000 670.000000 685.590000 ;
      RECT 657.500000 682.410000 658.500000 683.590000 ;
      RECT 616.500000 682.410000 649.500000 683.590000 ;
      RECT 607.500000 682.410000 608.500000 683.590000 ;
      RECT 566.500000 682.410000 599.500000 683.590000 ;
      RECT 557.500000 682.410000 558.500000 683.590000 ;
      RECT 516.500000 682.410000 549.500000 683.590000 ;
      RECT 507.500000 682.410000 508.500000 683.590000 ;
      RECT 466.500000 682.410000 499.500000 683.590000 ;
      RECT 457.500000 682.410000 458.500000 683.590000 ;
      RECT 416.500000 682.410000 449.500000 683.590000 ;
      RECT 407.500000 682.410000 408.500000 683.590000 ;
      RECT 366.500000 682.410000 373.500000 683.590000 ;
      RECT 357.500000 682.410000 358.500000 683.590000 ;
      RECT 316.500000 682.410000 349.500000 683.590000 ;
      RECT 307.500000 682.410000 308.500000 683.590000 ;
      RECT 1157.500000 681.590000 1186.000000 682.410000 ;
      RECT 657.500000 681.590000 670.000000 682.410000 ;
      RECT 607.500000 681.590000 649.500000 682.410000 ;
      RECT 557.500000 681.590000 599.500000 682.410000 ;
      RECT 507.500000 681.590000 549.500000 682.410000 ;
      RECT 457.500000 681.590000 499.500000 682.410000 ;
      RECT 407.500000 681.590000 449.500000 682.410000 ;
      RECT 357.500000 681.590000 373.500000 682.410000 ;
      RECT 307.500000 681.590000 349.500000 682.410000 ;
      RECT 1157.500000 680.410000 1158.500000 681.590000 ;
      RECT 1139.000000 680.410000 1149.500000 683.590000 ;
      RECT 657.500000 680.410000 658.500000 681.590000 ;
      RECT 616.500000 680.410000 649.500000 681.590000 ;
      RECT 607.500000 680.410000 608.500000 681.590000 ;
      RECT 566.500000 680.410000 599.500000 681.590000 ;
      RECT 557.500000 680.410000 558.500000 681.590000 ;
      RECT 516.500000 680.410000 549.500000 681.590000 ;
      RECT 507.500000 680.410000 508.500000 681.590000 ;
      RECT 466.500000 680.410000 499.500000 681.590000 ;
      RECT 457.500000 680.410000 458.500000 681.590000 ;
      RECT 416.500000 680.410000 449.500000 681.590000 ;
      RECT 407.500000 680.410000 408.500000 681.590000 ;
      RECT 386.500000 680.410000 399.500000 683.590000 ;
      RECT 366.500000 680.410000 373.500000 681.590000 ;
      RECT 357.500000 680.410000 358.500000 681.590000 ;
      RECT 316.500000 680.410000 349.500000 681.590000 ;
      RECT 307.500000 680.410000 308.500000 681.590000 ;
      RECT 0.000000 680.410000 299.500000 683.590000 ;
      RECT 1139.000000 679.590000 1158.500000 680.410000 ;
      RECT 616.500000 679.590000 658.500000 680.410000 ;
      RECT 566.500000 679.590000 608.500000 680.410000 ;
      RECT 516.500000 679.590000 558.500000 680.410000 ;
      RECT 466.500000 679.590000 508.500000 680.410000 ;
      RECT 416.500000 679.590000 458.500000 680.410000 ;
      RECT 366.500000 679.590000 408.500000 680.410000 ;
      RECT 316.500000 679.590000 358.500000 680.410000 ;
      RECT 0.000000 679.590000 308.500000 680.410000 ;
      RECT 1166.500000 678.410000 1186.000000 681.590000 ;
      RECT 1157.500000 678.410000 1158.500000 679.590000 ;
      RECT 666.500000 678.410000 670.000000 681.590000 ;
      RECT 657.500000 678.410000 658.500000 679.590000 ;
      RECT 616.500000 678.410000 649.500000 679.590000 ;
      RECT 607.500000 678.410000 608.500000 679.590000 ;
      RECT 566.500000 678.410000 599.500000 679.590000 ;
      RECT 557.500000 678.410000 558.500000 679.590000 ;
      RECT 516.500000 678.410000 549.500000 679.590000 ;
      RECT 507.500000 678.410000 508.500000 679.590000 ;
      RECT 466.500000 678.410000 499.500000 679.590000 ;
      RECT 457.500000 678.410000 458.500000 679.590000 ;
      RECT 416.500000 678.410000 449.500000 679.590000 ;
      RECT 407.500000 678.410000 408.500000 679.590000 ;
      RECT 366.500000 678.410000 373.500000 679.590000 ;
      RECT 357.500000 678.410000 358.500000 679.590000 ;
      RECT 316.500000 678.410000 349.500000 679.590000 ;
      RECT 307.500000 678.410000 308.500000 679.590000 ;
      RECT 1157.500000 677.590000 1186.000000 678.410000 ;
      RECT 657.500000 677.590000 670.000000 678.410000 ;
      RECT 607.500000 677.590000 649.500000 678.410000 ;
      RECT 557.500000 677.590000 599.500000 678.410000 ;
      RECT 507.500000 677.590000 549.500000 678.410000 ;
      RECT 457.500000 677.590000 499.500000 678.410000 ;
      RECT 407.500000 677.590000 449.500000 678.410000 ;
      RECT 357.500000 677.590000 373.500000 678.410000 ;
      RECT 1157.500000 676.410000 1158.500000 677.590000 ;
      RECT 1139.000000 676.410000 1149.500000 679.590000 ;
      RECT 657.500000 676.410000 658.500000 677.590000 ;
      RECT 616.500000 676.410000 649.500000 677.590000 ;
      RECT 607.500000 676.410000 608.500000 677.590000 ;
      RECT 566.500000 676.410000 599.500000 677.590000 ;
      RECT 557.500000 676.410000 558.500000 677.590000 ;
      RECT 516.500000 676.410000 549.500000 677.590000 ;
      RECT 507.500000 676.410000 508.500000 677.590000 ;
      RECT 466.500000 676.410000 499.500000 677.590000 ;
      RECT 457.500000 676.410000 458.500000 677.590000 ;
      RECT 416.500000 676.410000 449.500000 677.590000 ;
      RECT 407.500000 676.410000 408.500000 677.590000 ;
      RECT 386.500000 676.410000 399.500000 679.590000 ;
      RECT 366.500000 676.410000 373.500000 677.590000 ;
      RECT 357.500000 676.410000 358.500000 677.590000 ;
      RECT 307.500000 676.410000 349.500000 678.410000 ;
      RECT 0.000000 676.410000 299.500000 679.590000 ;
      RECT 1139.000000 675.590000 1158.500000 676.410000 ;
      RECT 616.500000 675.590000 658.500000 676.410000 ;
      RECT 566.500000 675.590000 608.500000 676.410000 ;
      RECT 516.500000 675.590000 558.500000 676.410000 ;
      RECT 466.500000 675.590000 508.500000 676.410000 ;
      RECT 416.500000 675.590000 458.500000 676.410000 ;
      RECT 366.500000 675.590000 408.500000 676.410000 ;
      RECT 0.000000 675.590000 358.500000 676.410000 ;
      RECT 1166.500000 674.410000 1186.000000 677.590000 ;
      RECT 1157.500000 674.410000 1158.500000 675.590000 ;
      RECT 666.500000 674.410000 670.000000 677.590000 ;
      RECT 657.500000 674.410000 658.500000 675.590000 ;
      RECT 616.500000 674.410000 649.500000 675.590000 ;
      RECT 607.500000 674.410000 608.500000 675.590000 ;
      RECT 566.500000 674.410000 599.500000 675.590000 ;
      RECT 557.500000 674.410000 558.500000 675.590000 ;
      RECT 516.500000 674.410000 549.500000 675.590000 ;
      RECT 507.500000 674.410000 508.500000 675.590000 ;
      RECT 466.500000 674.410000 499.500000 675.590000 ;
      RECT 457.500000 674.410000 458.500000 675.590000 ;
      RECT 416.500000 674.410000 449.500000 675.590000 ;
      RECT 407.500000 674.410000 408.500000 675.590000 ;
      RECT 366.500000 674.410000 373.500000 675.590000 ;
      RECT 357.500000 674.410000 358.500000 675.590000 ;
      RECT 1157.500000 673.590000 1186.000000 674.410000 ;
      RECT 657.500000 673.590000 670.000000 674.410000 ;
      RECT 607.500000 673.590000 649.500000 674.410000 ;
      RECT 557.500000 673.590000 599.500000 674.410000 ;
      RECT 507.500000 673.590000 549.500000 674.410000 ;
      RECT 457.500000 673.590000 499.500000 674.410000 ;
      RECT 407.500000 673.590000 449.500000 674.410000 ;
      RECT 357.500000 673.590000 373.500000 674.410000 ;
      RECT 1157.500000 672.410000 1158.500000 673.590000 ;
      RECT 1139.000000 672.410000 1149.500000 675.590000 ;
      RECT 657.500000 672.410000 658.500000 673.590000 ;
      RECT 616.500000 672.410000 649.500000 673.590000 ;
      RECT 607.500000 672.410000 608.500000 673.590000 ;
      RECT 566.500000 672.410000 599.500000 673.590000 ;
      RECT 557.500000 672.410000 558.500000 673.590000 ;
      RECT 516.500000 672.410000 549.500000 673.590000 ;
      RECT 507.500000 672.410000 508.500000 673.590000 ;
      RECT 466.500000 672.410000 499.500000 673.590000 ;
      RECT 457.500000 672.410000 458.500000 673.590000 ;
      RECT 416.500000 672.410000 449.500000 673.590000 ;
      RECT 407.500000 672.410000 408.500000 673.590000 ;
      RECT 386.500000 672.410000 399.500000 675.590000 ;
      RECT 366.500000 672.410000 373.500000 673.590000 ;
      RECT 357.500000 672.410000 358.500000 673.590000 ;
      RECT 0.000000 672.410000 349.500000 675.590000 ;
      RECT 1139.000000 671.590000 1158.500000 672.410000 ;
      RECT 616.500000 671.590000 658.500000 672.410000 ;
      RECT 566.500000 671.590000 608.500000 672.410000 ;
      RECT 516.500000 671.590000 558.500000 672.410000 ;
      RECT 466.500000 671.590000 508.500000 672.410000 ;
      RECT 416.500000 671.590000 458.500000 672.410000 ;
      RECT 366.500000 671.590000 408.500000 672.410000 ;
      RECT 0.000000 671.590000 358.500000 672.410000 ;
      RECT 1166.500000 670.410000 1186.000000 673.590000 ;
      RECT 1157.500000 670.410000 1158.500000 671.590000 ;
      RECT 666.500000 670.410000 670.000000 673.590000 ;
      RECT 657.500000 670.410000 658.500000 671.590000 ;
      RECT 616.500000 670.410000 649.500000 671.590000 ;
      RECT 607.500000 670.410000 608.500000 671.590000 ;
      RECT 566.500000 670.410000 599.500000 671.590000 ;
      RECT 557.500000 670.410000 558.500000 671.590000 ;
      RECT 516.500000 670.410000 549.500000 671.590000 ;
      RECT 507.500000 670.410000 508.500000 671.590000 ;
      RECT 466.500000 670.410000 499.500000 671.590000 ;
      RECT 457.500000 670.410000 458.500000 671.590000 ;
      RECT 416.500000 670.410000 449.500000 671.590000 ;
      RECT 407.500000 670.410000 408.500000 671.590000 ;
      RECT 366.500000 670.410000 373.500000 671.590000 ;
      RECT 357.500000 670.410000 358.500000 671.590000 ;
      RECT 1157.500000 669.590000 1186.000000 670.410000 ;
      RECT 657.500000 669.590000 670.000000 670.410000 ;
      RECT 607.500000 669.590000 649.500000 670.410000 ;
      RECT 557.500000 669.590000 599.500000 670.410000 ;
      RECT 507.500000 669.590000 549.500000 670.410000 ;
      RECT 457.500000 669.590000 499.500000 670.410000 ;
      RECT 407.500000 669.590000 449.500000 670.410000 ;
      RECT 357.500000 669.590000 373.500000 670.410000 ;
      RECT 1157.500000 668.410000 1158.500000 669.590000 ;
      RECT 1139.000000 668.410000 1149.500000 671.590000 ;
      RECT 657.500000 668.410000 658.500000 669.590000 ;
      RECT 616.500000 668.410000 649.500000 669.590000 ;
      RECT 607.500000 668.410000 608.500000 669.590000 ;
      RECT 566.500000 668.410000 599.500000 669.590000 ;
      RECT 557.500000 668.410000 558.500000 669.590000 ;
      RECT 516.500000 668.410000 549.500000 669.590000 ;
      RECT 507.500000 668.410000 508.500000 669.590000 ;
      RECT 466.500000 668.410000 499.500000 669.590000 ;
      RECT 457.500000 668.410000 458.500000 669.590000 ;
      RECT 416.500000 668.410000 449.500000 669.590000 ;
      RECT 407.500000 668.410000 408.500000 669.590000 ;
      RECT 386.500000 668.410000 399.500000 671.590000 ;
      RECT 372.500000 668.410000 373.500000 669.590000 ;
      RECT 357.500000 668.410000 358.500000 669.590000 ;
      RECT 0.000000 668.410000 349.500000 671.590000 ;
      RECT 1139.000000 667.590000 1158.500000 668.410000 ;
      RECT 616.500000 667.590000 658.500000 668.410000 ;
      RECT 566.500000 667.590000 608.500000 668.410000 ;
      RECT 516.500000 667.590000 558.500000 668.410000 ;
      RECT 466.500000 667.590000 508.500000 668.410000 ;
      RECT 416.500000 667.590000 458.500000 668.410000 ;
      RECT 372.500000 667.590000 408.500000 668.410000 ;
      RECT 0.000000 667.590000 358.500000 668.410000 ;
      RECT 1166.500000 666.410000 1186.000000 669.590000 ;
      RECT 1157.500000 666.410000 1158.500000 667.590000 ;
      RECT 666.500000 666.410000 670.000000 669.590000 ;
      RECT 657.500000 666.410000 658.500000 667.590000 ;
      RECT 616.500000 666.410000 649.500000 667.590000 ;
      RECT 607.500000 666.410000 608.500000 667.590000 ;
      RECT 566.500000 666.410000 599.500000 667.590000 ;
      RECT 557.500000 666.410000 558.500000 667.590000 ;
      RECT 516.500000 666.410000 549.500000 667.590000 ;
      RECT 507.500000 666.410000 508.500000 667.590000 ;
      RECT 466.500000 666.410000 499.500000 667.590000 ;
      RECT 457.500000 666.410000 458.500000 667.590000 ;
      RECT 416.500000 666.410000 449.500000 667.590000 ;
      RECT 407.500000 666.410000 408.500000 667.590000 ;
      RECT 372.500000 666.410000 373.500000 667.590000 ;
      RECT 357.500000 666.410000 358.500000 667.590000 ;
      RECT 1157.500000 665.590000 1186.000000 666.410000 ;
      RECT 657.500000 665.590000 670.000000 666.410000 ;
      RECT 607.500000 665.590000 649.500000 666.410000 ;
      RECT 557.500000 665.590000 599.500000 666.410000 ;
      RECT 507.500000 665.590000 549.500000 666.410000 ;
      RECT 457.500000 665.590000 499.500000 666.410000 ;
      RECT 407.500000 665.590000 449.500000 666.410000 ;
      RECT 357.500000 665.590000 373.500000 666.410000 ;
      RECT 1157.500000 664.410000 1158.500000 665.590000 ;
      RECT 1139.000000 664.410000 1149.500000 667.590000 ;
      RECT 657.500000 664.410000 658.500000 665.590000 ;
      RECT 616.500000 664.410000 649.500000 665.590000 ;
      RECT 607.500000 664.410000 608.500000 665.590000 ;
      RECT 566.500000 664.410000 599.500000 665.590000 ;
      RECT 557.500000 664.410000 558.500000 665.590000 ;
      RECT 516.500000 664.410000 549.500000 665.590000 ;
      RECT 507.500000 664.410000 508.500000 665.590000 ;
      RECT 466.500000 664.410000 499.500000 665.590000 ;
      RECT 457.500000 664.410000 458.500000 665.590000 ;
      RECT 416.500000 664.410000 449.500000 665.590000 ;
      RECT 407.500000 664.410000 408.500000 665.590000 ;
      RECT 386.500000 664.410000 399.500000 667.590000 ;
      RECT 372.500000 664.410000 373.500000 665.590000 ;
      RECT 357.500000 664.410000 358.500000 665.590000 ;
      RECT 0.000000 664.410000 349.500000 667.590000 ;
      RECT 1139.000000 663.590000 1158.500000 664.410000 ;
      RECT 616.500000 663.590000 658.500000 664.410000 ;
      RECT 566.500000 663.590000 608.500000 664.410000 ;
      RECT 516.500000 663.590000 558.500000 664.410000 ;
      RECT 466.500000 663.590000 508.500000 664.410000 ;
      RECT 416.500000 663.590000 458.500000 664.410000 ;
      RECT 372.500000 663.590000 408.500000 664.410000 ;
      RECT 0.000000 663.590000 358.500000 664.410000 ;
      RECT 0.000000 663.170000 349.500000 663.590000 ;
      RECT 1166.500000 663.165000 1186.000000 665.590000 ;
      RECT 1166.500000 662.410000 1183.980000 663.165000 ;
      RECT 1157.500000 662.410000 1158.500000 663.590000 ;
      RECT 666.500000 662.410000 670.000000 665.590000 ;
      RECT 657.500000 662.410000 658.500000 663.590000 ;
      RECT 616.500000 662.410000 649.500000 663.590000 ;
      RECT 607.500000 662.410000 608.500000 663.590000 ;
      RECT 566.500000 662.410000 599.500000 663.590000 ;
      RECT 557.500000 662.410000 558.500000 663.590000 ;
      RECT 516.500000 662.410000 549.500000 663.590000 ;
      RECT 507.500000 662.410000 508.500000 663.590000 ;
      RECT 466.500000 662.410000 499.500000 663.590000 ;
      RECT 457.500000 662.410000 458.500000 663.590000 ;
      RECT 416.500000 662.410000 449.500000 663.590000 ;
      RECT 407.500000 662.410000 408.500000 663.590000 ;
      RECT 372.500000 662.410000 373.500000 663.590000 ;
      RECT 357.500000 662.410000 358.500000 663.590000 ;
      RECT 1157.500000 661.590000 1183.980000 662.410000 ;
      RECT 657.500000 661.590000 670.000000 662.410000 ;
      RECT 607.500000 661.590000 649.500000 662.410000 ;
      RECT 557.500000 661.590000 599.500000 662.410000 ;
      RECT 507.500000 661.590000 549.500000 662.410000 ;
      RECT 457.500000 661.590000 499.500000 662.410000 ;
      RECT 407.500000 661.590000 449.500000 662.410000 ;
      RECT 357.500000 661.590000 373.500000 662.410000 ;
      RECT 1157.500000 660.410000 1158.500000 661.590000 ;
      RECT 1139.000000 660.410000 1149.500000 663.590000 ;
      RECT 657.500000 660.410000 658.500000 661.590000 ;
      RECT 616.500000 660.410000 649.500000 661.590000 ;
      RECT 607.500000 660.410000 608.500000 661.590000 ;
      RECT 566.500000 660.410000 599.500000 661.590000 ;
      RECT 557.500000 660.410000 558.500000 661.590000 ;
      RECT 516.500000 660.410000 549.500000 661.590000 ;
      RECT 507.500000 660.410000 508.500000 661.590000 ;
      RECT 466.500000 660.410000 499.500000 661.590000 ;
      RECT 457.500000 660.410000 458.500000 661.590000 ;
      RECT 416.500000 660.410000 449.500000 661.590000 ;
      RECT 407.500000 660.410000 408.500000 661.590000 ;
      RECT 386.500000 660.410000 399.500000 663.590000 ;
      RECT 372.500000 660.410000 373.500000 661.590000 ;
      RECT 357.500000 660.410000 358.500000 661.590000 ;
      RECT 2.020000 660.410000 349.500000 663.170000 ;
      RECT 2.020000 660.070000 358.500000 660.410000 ;
      RECT 1166.500000 660.065000 1183.980000 661.590000 ;
      RECT 1139.000000 659.590000 1158.500000 660.410000 ;
      RECT 616.500000 659.590000 658.500000 660.410000 ;
      RECT 566.500000 659.590000 608.500000 660.410000 ;
      RECT 516.500000 659.590000 558.500000 660.410000 ;
      RECT 466.500000 659.590000 508.500000 660.410000 ;
      RECT 416.500000 659.590000 458.500000 660.410000 ;
      RECT 372.500000 659.590000 408.500000 660.410000 ;
      RECT 0.000000 659.590000 358.500000 660.070000 ;
      RECT 1166.500000 658.410000 1186.000000 660.065000 ;
      RECT 1157.500000 658.410000 1158.500000 659.590000 ;
      RECT 666.500000 658.410000 670.000000 661.590000 ;
      RECT 657.500000 658.410000 658.500000 659.590000 ;
      RECT 616.500000 658.410000 649.500000 659.590000 ;
      RECT 607.500000 658.410000 608.500000 659.590000 ;
      RECT 566.500000 658.410000 599.500000 659.590000 ;
      RECT 557.500000 658.410000 558.500000 659.590000 ;
      RECT 516.500000 658.410000 549.500000 659.590000 ;
      RECT 507.500000 658.410000 508.500000 659.590000 ;
      RECT 466.500000 658.410000 499.500000 659.590000 ;
      RECT 457.500000 658.410000 458.500000 659.590000 ;
      RECT 416.500000 658.410000 449.500000 659.590000 ;
      RECT 407.500000 658.410000 408.500000 659.590000 ;
      RECT 372.500000 658.410000 373.500000 659.590000 ;
      RECT 357.500000 658.410000 358.500000 659.590000 ;
      RECT 1157.500000 657.590000 1186.000000 658.410000 ;
      RECT 357.500000 657.590000 373.500000 658.410000 ;
      RECT 1166.500000 657.485000 1186.000000 657.590000 ;
      RECT 1157.500000 656.410000 1158.500000 657.590000 ;
      RECT 1139.000000 656.410000 1149.500000 659.590000 ;
      RECT 657.500000 656.410000 670.000000 658.410000 ;
      RECT 607.500000 656.410000 649.500000 658.410000 ;
      RECT 557.500000 656.410000 599.500000 658.410000 ;
      RECT 507.500000 656.410000 549.500000 658.410000 ;
      RECT 457.500000 656.410000 499.500000 658.410000 ;
      RECT 407.500000 656.410000 449.500000 658.410000 ;
      RECT 386.500000 656.410000 399.500000 659.590000 ;
      RECT 372.500000 656.410000 373.500000 657.590000 ;
      RECT 357.500000 656.410000 358.500000 657.590000 ;
      RECT 0.000000 656.410000 349.500000 659.590000 ;
      RECT 372.500000 656.000000 670.000000 656.410000 ;
      RECT 1139.000000 655.590000 1158.500000 656.410000 ;
      RECT 372.500000 655.590000 389.000000 656.000000 ;
      RECT 0.000000 655.590000 358.500000 656.410000 ;
      RECT 1166.500000 654.410000 1183.980000 657.485000 ;
      RECT 1157.500000 654.410000 1158.500000 655.590000 ;
      RECT 372.500000 654.410000 373.500000 655.590000 ;
      RECT 357.500000 654.410000 358.500000 655.590000 ;
      RECT 1157.500000 654.385000 1183.980000 654.410000 ;
      RECT 1157.500000 653.590000 1186.000000 654.385000 ;
      RECT 357.500000 653.590000 373.500000 654.410000 ;
      RECT 1166.500000 653.525000 1186.000000 653.590000 ;
      RECT 0.000000 652.575000 349.500000 655.590000 ;
      RECT 1157.500000 652.410000 1158.500000 653.590000 ;
      RECT 1139.000000 652.410000 1149.500000 655.590000 ;
      RECT 386.500000 652.410000 389.000000 655.590000 ;
      RECT 372.500000 652.410000 373.500000 653.590000 ;
      RECT 357.500000 652.410000 358.500000 653.590000 ;
      RECT 2.020000 652.410000 349.500000 652.575000 ;
      RECT 1139.000000 651.590000 1158.500000 652.410000 ;
      RECT 372.500000 651.590000 389.000000 652.410000 ;
      RECT 2.020000 651.590000 358.500000 652.410000 ;
      RECT 1166.500000 650.425000 1183.980000 653.525000 ;
      RECT 1166.500000 650.410000 1186.000000 650.425000 ;
      RECT 1157.500000 650.410000 1158.500000 651.590000 ;
      RECT 372.500000 650.410000 373.500000 651.590000 ;
      RECT 357.500000 650.410000 358.500000 651.590000 ;
      RECT 1157.500000 649.590000 1186.000000 650.410000 ;
      RECT 357.500000 649.590000 373.500000 650.410000 ;
      RECT 2.020000 649.475000 349.500000 651.590000 ;
      RECT 0.000000 648.615000 349.500000 649.475000 ;
      RECT 1157.500000 648.410000 1158.500000 649.590000 ;
      RECT 1139.000000 648.410000 1149.500000 651.590000 ;
      RECT 386.500000 648.410000 389.000000 651.590000 ;
      RECT 372.500000 648.410000 373.500000 649.590000 ;
      RECT 357.500000 648.410000 358.500000 649.590000 ;
      RECT 2.020000 648.410000 349.500000 648.615000 ;
      RECT 1139.000000 647.590000 1158.500000 648.410000 ;
      RECT 372.500000 647.590000 389.000000 648.410000 ;
      RECT 2.020000 647.590000 358.500000 648.410000 ;
      RECT 1166.500000 646.410000 1186.000000 649.590000 ;
      RECT 1157.500000 646.410000 1158.500000 647.590000 ;
      RECT 372.500000 646.410000 373.500000 647.590000 ;
      RECT 357.500000 646.410000 358.500000 647.590000 ;
      RECT 1157.500000 645.590000 1186.000000 646.410000 ;
      RECT 357.500000 645.590000 373.500000 646.410000 ;
      RECT 2.020000 645.515000 349.500000 647.590000 ;
      RECT 1157.500000 644.410000 1158.500000 645.590000 ;
      RECT 1139.000000 644.410000 1149.500000 647.590000 ;
      RECT 386.500000 644.410000 389.000000 647.590000 ;
      RECT 372.500000 644.410000 373.500000 645.590000 ;
      RECT 357.500000 644.410000 358.500000 645.590000 ;
      RECT 0.000000 644.410000 349.500000 645.515000 ;
      RECT 1139.000000 643.590000 1158.500000 644.410000 ;
      RECT 372.500000 643.590000 389.000000 644.410000 ;
      RECT 0.000000 643.590000 358.500000 644.410000 ;
      RECT 0.000000 642.935000 349.500000 643.590000 ;
      RECT 1166.500000 642.930000 1186.000000 645.590000 ;
      RECT 1166.500000 642.410000 1183.980000 642.930000 ;
      RECT 1157.500000 642.410000 1158.500000 643.590000 ;
      RECT 372.500000 642.410000 373.500000 643.590000 ;
      RECT 357.500000 642.410000 358.500000 643.590000 ;
      RECT 1157.500000 641.590000 1183.980000 642.410000 ;
      RECT 357.500000 641.590000 373.500000 642.410000 ;
      RECT 1157.500000 640.410000 1158.500000 641.590000 ;
      RECT 1139.000000 640.410000 1149.500000 643.590000 ;
      RECT 386.500000 640.410000 389.000000 643.590000 ;
      RECT 372.500000 640.410000 373.500000 641.590000 ;
      RECT 357.500000 640.410000 358.500000 641.590000 ;
      RECT 2.020000 640.410000 349.500000 642.935000 ;
      RECT 2.020000 639.835000 358.500000 640.410000 ;
      RECT 1166.500000 639.830000 1183.980000 641.590000 ;
      RECT 1139.000000 639.590000 1158.500000 640.410000 ;
      RECT 372.500000 639.590000 389.000000 640.410000 ;
      RECT 0.000000 639.590000 358.500000 639.835000 ;
      RECT 1166.500000 638.410000 1186.000000 639.830000 ;
      RECT 1157.500000 638.410000 1158.500000 639.590000 ;
      RECT 372.500000 638.410000 373.500000 639.590000 ;
      RECT 357.500000 638.410000 358.500000 639.590000 ;
      RECT 1157.500000 637.590000 1186.000000 638.410000 ;
      RECT 357.500000 637.590000 373.500000 638.410000 ;
      RECT 1157.500000 636.410000 1158.500000 637.590000 ;
      RECT 1139.000000 636.410000 1149.500000 639.590000 ;
      RECT 386.500000 636.410000 389.000000 639.590000 ;
      RECT 372.500000 636.410000 373.500000 637.590000 ;
      RECT 357.500000 636.410000 358.500000 637.590000 ;
      RECT 0.000000 636.410000 349.500000 639.590000 ;
      RECT 1139.000000 635.590000 1158.500000 636.410000 ;
      RECT 372.500000 635.590000 389.000000 636.410000 ;
      RECT 0.000000 635.590000 358.500000 636.410000 ;
      RECT 1166.500000 634.410000 1186.000000 637.590000 ;
      RECT 1157.500000 634.410000 1158.500000 635.590000 ;
      RECT 372.500000 634.410000 373.500000 635.590000 ;
      RECT 357.500000 634.410000 358.500000 635.590000 ;
      RECT 1157.500000 633.590000 1186.000000 634.410000 ;
      RECT 357.500000 633.590000 373.500000 634.410000 ;
      RECT 1157.500000 632.410000 1158.500000 633.590000 ;
      RECT 1139.000000 632.410000 1149.500000 635.590000 ;
      RECT 386.500000 632.410000 389.000000 635.590000 ;
      RECT 372.500000 632.410000 373.500000 633.590000 ;
      RECT 357.500000 632.410000 358.500000 633.590000 ;
      RECT 0.000000 632.410000 349.500000 635.590000 ;
      RECT 1139.000000 631.590000 1158.500000 632.410000 ;
      RECT 372.500000 631.590000 389.000000 632.410000 ;
      RECT 0.000000 631.590000 358.500000 632.410000 ;
      RECT 1166.500000 630.410000 1186.000000 633.590000 ;
      RECT 1157.500000 630.410000 1158.500000 631.590000 ;
      RECT 372.500000 630.410000 373.500000 631.590000 ;
      RECT 357.500000 630.410000 358.500000 631.590000 ;
      RECT 1157.500000 629.590000 1186.000000 630.410000 ;
      RECT 357.500000 629.590000 373.500000 630.410000 ;
      RECT 1157.500000 628.410000 1158.500000 629.590000 ;
      RECT 1139.000000 628.410000 1149.500000 631.590000 ;
      RECT 386.500000 628.410000 389.000000 631.590000 ;
      RECT 372.500000 628.410000 373.500000 629.590000 ;
      RECT 357.500000 628.410000 358.500000 629.590000 ;
      RECT 0.000000 628.410000 349.500000 631.590000 ;
      RECT 1139.000000 627.590000 1158.500000 628.410000 ;
      RECT 372.500000 627.590000 389.000000 628.410000 ;
      RECT 0.000000 627.590000 358.500000 628.410000 ;
      RECT 1166.500000 626.410000 1186.000000 629.590000 ;
      RECT 1157.500000 626.410000 1158.500000 627.590000 ;
      RECT 372.500000 626.410000 373.500000 627.590000 ;
      RECT 357.500000 626.410000 358.500000 627.590000 ;
      RECT 1157.500000 625.590000 1186.000000 626.410000 ;
      RECT 357.500000 625.590000 373.500000 626.410000 ;
      RECT 1157.500000 624.410000 1158.500000 625.590000 ;
      RECT 1139.000000 624.410000 1149.500000 627.590000 ;
      RECT 386.500000 624.410000 389.000000 627.590000 ;
      RECT 372.500000 624.410000 373.500000 625.590000 ;
      RECT 357.500000 624.410000 358.500000 625.590000 ;
      RECT 0.000000 624.410000 349.500000 627.590000 ;
      RECT 1139.000000 623.590000 1158.500000 624.410000 ;
      RECT 372.500000 623.590000 389.000000 624.410000 ;
      RECT 0.000000 623.590000 358.500000 624.410000 ;
      RECT 1166.500000 622.410000 1186.000000 625.590000 ;
      RECT 1157.500000 622.410000 1158.500000 623.590000 ;
      RECT 372.500000 622.410000 373.500000 623.590000 ;
      RECT 357.500000 622.410000 358.500000 623.590000 ;
      RECT 1157.500000 621.590000 1186.000000 622.410000 ;
      RECT 357.500000 621.590000 373.500000 622.410000 ;
      RECT 1157.500000 620.410000 1158.500000 621.590000 ;
      RECT 1139.000000 620.410000 1149.500000 623.590000 ;
      RECT 386.500000 620.410000 389.000000 623.590000 ;
      RECT 372.500000 620.410000 373.500000 621.590000 ;
      RECT 357.500000 620.410000 358.500000 621.590000 ;
      RECT 0.000000 620.410000 349.500000 623.590000 ;
      RECT 1139.000000 619.590000 1158.500000 620.410000 ;
      RECT 372.500000 619.590000 389.000000 620.410000 ;
      RECT 0.000000 619.590000 358.500000 620.410000 ;
      RECT 1166.500000 618.410000 1186.000000 621.590000 ;
      RECT 1157.500000 618.410000 1158.500000 619.590000 ;
      RECT 372.500000 618.410000 373.500000 619.590000 ;
      RECT 357.500000 618.410000 358.500000 619.590000 ;
      RECT 1157.500000 617.590000 1186.000000 618.410000 ;
      RECT 357.500000 617.590000 373.500000 618.410000 ;
      RECT 1157.500000 616.410000 1158.500000 617.590000 ;
      RECT 1139.000000 616.410000 1149.500000 619.590000 ;
      RECT 386.500000 616.410000 389.000000 619.590000 ;
      RECT 372.500000 616.410000 373.500000 617.590000 ;
      RECT 357.500000 616.410000 358.500000 617.590000 ;
      RECT 0.000000 616.410000 349.500000 619.590000 ;
      RECT 372.500000 616.115000 389.000000 616.410000 ;
      RECT 1139.000000 615.695000 1158.500000 616.410000 ;
      RECT 1141.020000 615.590000 1158.500000 615.695000 ;
      RECT 372.500000 615.590000 386.980000 616.115000 ;
      RECT 0.000000 615.590000 358.500000 616.410000 ;
      RECT 1166.500000 614.410000 1186.000000 617.590000 ;
      RECT 1157.500000 614.410000 1158.500000 615.590000 ;
      RECT 372.500000 614.410000 373.500000 615.590000 ;
      RECT 357.500000 614.410000 358.500000 615.590000 ;
      RECT 1157.500000 613.590000 1186.000000 614.410000 ;
      RECT 357.500000 613.590000 373.500000 614.410000 ;
      RECT 1157.500000 612.410000 1158.500000 613.590000 ;
      RECT 1141.020000 612.410000 1149.500000 615.590000 ;
      RECT 386.500000 612.410000 386.980000 615.590000 ;
      RECT 372.500000 612.410000 373.500000 613.590000 ;
      RECT 357.500000 612.410000 358.500000 613.590000 ;
      RECT 0.000000 612.410000 349.500000 615.590000 ;
      RECT 1141.020000 611.590000 1158.500000 612.410000 ;
      RECT 372.500000 611.590000 386.980000 612.410000 ;
      RECT 0.000000 611.590000 358.500000 612.410000 ;
      RECT 1166.500000 610.410000 1186.000000 613.590000 ;
      RECT 1157.500000 610.410000 1158.500000 611.590000 ;
      RECT 372.500000 610.410000 373.500000 611.590000 ;
      RECT 357.500000 610.410000 358.500000 611.590000 ;
      RECT 1157.500000 609.590000 1186.000000 610.410000 ;
      RECT 357.500000 609.590000 373.500000 610.410000 ;
      RECT 1157.500000 608.410000 1158.500000 609.590000 ;
      RECT 1141.020000 608.410000 1149.500000 611.590000 ;
      RECT 386.500000 608.410000 386.980000 611.590000 ;
      RECT 372.500000 608.410000 373.500000 609.590000 ;
      RECT 357.500000 608.410000 358.500000 609.590000 ;
      RECT 0.000000 608.410000 349.500000 611.590000 ;
      RECT 1141.020000 607.590000 1158.500000 608.410000 ;
      RECT 372.500000 607.590000 386.980000 608.410000 ;
      RECT 0.000000 607.590000 358.500000 608.410000 ;
      RECT 1166.500000 606.410000 1186.000000 609.590000 ;
      RECT 1157.500000 606.410000 1158.500000 607.590000 ;
      RECT 372.500000 606.410000 373.500000 607.590000 ;
      RECT 357.500000 606.410000 358.500000 607.590000 ;
      RECT 1157.500000 605.590000 1186.000000 606.410000 ;
      RECT 357.500000 605.590000 373.500000 606.410000 ;
      RECT 1157.500000 604.410000 1158.500000 605.590000 ;
      RECT 1141.020000 604.410000 1149.500000 607.590000 ;
      RECT 386.500000 604.410000 386.980000 607.590000 ;
      RECT 372.500000 604.410000 373.500000 605.590000 ;
      RECT 357.500000 604.410000 358.500000 605.590000 ;
      RECT 0.000000 604.410000 349.500000 607.590000 ;
      RECT 1141.020000 603.590000 1158.500000 604.410000 ;
      RECT 372.500000 603.590000 386.980000 604.410000 ;
      RECT 0.000000 603.590000 358.500000 604.410000 ;
      RECT 1166.500000 602.410000 1186.000000 605.590000 ;
      RECT 1157.500000 602.410000 1158.500000 603.590000 ;
      RECT 372.500000 602.410000 373.500000 603.590000 ;
      RECT 357.500000 602.410000 358.500000 603.590000 ;
      RECT 1157.500000 601.590000 1186.000000 602.410000 ;
      RECT 357.500000 601.590000 373.500000 602.410000 ;
      RECT 1157.500000 600.410000 1158.500000 601.590000 ;
      RECT 1141.020000 600.410000 1149.500000 603.590000 ;
      RECT 386.500000 600.410000 386.980000 603.590000 ;
      RECT 372.500000 600.410000 373.500000 601.590000 ;
      RECT 357.500000 600.410000 358.500000 601.590000 ;
      RECT 0.000000 600.410000 349.500000 603.590000 ;
      RECT 1141.020000 599.590000 1158.500000 600.410000 ;
      RECT 372.500000 599.590000 386.980000 600.410000 ;
      RECT 0.000000 599.590000 358.500000 600.410000 ;
      RECT 1166.500000 598.410000 1186.000000 601.590000 ;
      RECT 1157.500000 598.410000 1158.500000 599.590000 ;
      RECT 372.500000 598.410000 373.500000 599.590000 ;
      RECT 357.500000 598.410000 358.500000 599.590000 ;
      RECT 1141.020000 597.880000 1149.500000 599.590000 ;
      RECT 1157.500000 597.590000 1186.000000 598.410000 ;
      RECT 357.500000 597.590000 373.500000 598.410000 ;
      RECT 1157.500000 596.410000 1158.500000 597.590000 ;
      RECT 1139.000000 596.410000 1149.500000 597.880000 ;
      RECT 386.500000 596.410000 386.980000 599.590000 ;
      RECT 372.500000 596.410000 373.500000 597.590000 ;
      RECT 357.500000 596.410000 358.500000 597.590000 ;
      RECT 0.000000 596.410000 349.500000 599.590000 ;
      RECT 1139.000000 595.590000 1158.500000 596.410000 ;
      RECT 372.500000 595.590000 386.980000 596.410000 ;
      RECT 0.000000 595.590000 358.500000 596.410000 ;
      RECT 1166.500000 594.410000 1186.000000 597.590000 ;
      RECT 1157.500000 594.410000 1158.500000 595.590000 ;
      RECT 372.500000 594.410000 373.500000 595.590000 ;
      RECT 357.500000 594.410000 358.500000 595.590000 ;
      RECT 1157.500000 593.590000 1186.000000 594.410000 ;
      RECT 357.500000 593.590000 373.500000 594.410000 ;
      RECT 1157.500000 592.410000 1158.500000 593.590000 ;
      RECT 1139.000000 592.410000 1149.500000 595.590000 ;
      RECT 386.500000 592.410000 386.980000 595.590000 ;
      RECT 372.500000 592.410000 373.500000 593.590000 ;
      RECT 357.500000 592.410000 358.500000 593.590000 ;
      RECT 0.000000 592.410000 349.500000 595.590000 ;
      RECT 1139.000000 591.590000 1158.500000 592.410000 ;
      RECT 372.500000 591.590000 386.980000 592.410000 ;
      RECT 0.000000 591.590000 358.500000 592.410000 ;
      RECT 1166.500000 590.410000 1186.000000 593.590000 ;
      RECT 1157.500000 590.410000 1158.500000 591.590000 ;
      RECT 372.500000 590.410000 373.500000 591.590000 ;
      RECT 357.500000 590.410000 358.500000 591.590000 ;
      RECT 1157.500000 589.590000 1186.000000 590.410000 ;
      RECT 357.500000 589.590000 373.500000 590.410000 ;
      RECT 1157.500000 588.410000 1158.500000 589.590000 ;
      RECT 1139.000000 588.410000 1149.500000 591.590000 ;
      RECT 386.500000 588.410000 386.980000 591.590000 ;
      RECT 372.500000 588.410000 373.500000 589.590000 ;
      RECT 357.500000 588.410000 358.500000 589.590000 ;
      RECT 0.000000 588.410000 349.500000 591.590000 ;
      RECT 1139.000000 587.590000 1158.500000 588.410000 ;
      RECT 372.500000 587.590000 386.980000 588.410000 ;
      RECT 0.000000 587.590000 358.500000 588.410000 ;
      RECT 1166.500000 586.410000 1186.000000 589.590000 ;
      RECT 1157.500000 586.410000 1158.500000 587.590000 ;
      RECT 372.500000 586.410000 373.500000 587.590000 ;
      RECT 357.500000 586.410000 358.500000 587.590000 ;
      RECT 1157.500000 585.590000 1186.000000 586.410000 ;
      RECT 357.500000 585.590000 373.500000 586.410000 ;
      RECT 1157.500000 584.410000 1158.500000 585.590000 ;
      RECT 1139.000000 584.410000 1149.500000 587.590000 ;
      RECT 386.500000 584.410000 386.980000 587.590000 ;
      RECT 372.500000 584.410000 373.500000 585.590000 ;
      RECT 357.500000 584.410000 358.500000 585.590000 ;
      RECT 0.000000 584.410000 349.500000 587.590000 ;
      RECT 1139.000000 583.590000 1158.500000 584.410000 ;
      RECT 372.500000 583.590000 386.980000 584.410000 ;
      RECT 0.000000 583.590000 358.500000 584.410000 ;
      RECT 1166.500000 582.410000 1186.000000 585.590000 ;
      RECT 1157.500000 582.410000 1158.500000 583.590000 ;
      RECT 372.500000 582.410000 373.500000 583.590000 ;
      RECT 357.500000 582.410000 358.500000 583.590000 ;
      RECT 1157.500000 581.590000 1186.000000 582.410000 ;
      RECT 357.500000 581.590000 373.500000 582.410000 ;
      RECT 1157.500000 580.410000 1158.500000 581.590000 ;
      RECT 1139.000000 580.410000 1149.500000 583.590000 ;
      RECT 386.500000 580.410000 386.980000 583.590000 ;
      RECT 372.500000 580.410000 373.500000 581.590000 ;
      RECT 357.500000 580.410000 358.500000 581.590000 ;
      RECT 0.000000 580.410000 349.500000 583.590000 ;
      RECT 1139.000000 579.590000 1158.500000 580.410000 ;
      RECT 372.500000 579.590000 386.980000 580.410000 ;
      RECT 0.000000 579.590000 358.500000 580.410000 ;
      RECT 1166.500000 578.410000 1186.000000 581.590000 ;
      RECT 1157.500000 578.410000 1158.500000 579.590000 ;
      RECT 372.500000 578.410000 373.500000 579.590000 ;
      RECT 357.500000 578.410000 358.500000 579.590000 ;
      RECT 1157.500000 577.590000 1186.000000 578.410000 ;
      RECT 386.500000 577.590000 386.980000 579.590000 ;
      RECT 357.500000 577.590000 373.500000 578.410000 ;
      RECT 1157.500000 576.410000 1158.500000 577.590000 ;
      RECT 1139.000000 576.410000 1149.500000 579.590000 ;
      RECT 386.500000 576.410000 389.000000 577.590000 ;
      RECT 372.500000 576.410000 373.500000 577.590000 ;
      RECT 357.500000 576.410000 358.500000 577.590000 ;
      RECT 0.000000 576.410000 349.500000 579.590000 ;
      RECT 1139.000000 575.590000 1158.500000 576.410000 ;
      RECT 372.500000 575.590000 389.000000 576.410000 ;
      RECT 0.000000 575.590000 358.500000 576.410000 ;
      RECT 0.000000 575.170000 349.500000 575.590000 ;
      RECT 1166.500000 575.165000 1186.000000 577.590000 ;
      RECT 1166.500000 574.410000 1183.980000 575.165000 ;
      RECT 1157.500000 574.410000 1158.500000 575.590000 ;
      RECT 372.500000 574.410000 373.500000 575.590000 ;
      RECT 357.500000 574.410000 358.500000 575.590000 ;
      RECT 1157.500000 573.590000 1183.980000 574.410000 ;
      RECT 357.500000 573.590000 373.500000 574.410000 ;
      RECT 1157.500000 572.410000 1158.500000 573.590000 ;
      RECT 1139.000000 572.410000 1149.500000 575.590000 ;
      RECT 386.500000 572.410000 389.000000 575.590000 ;
      RECT 372.500000 572.410000 373.500000 573.590000 ;
      RECT 357.500000 572.410000 358.500000 573.590000 ;
      RECT 2.020000 572.410000 349.500000 575.170000 ;
      RECT 2.020000 572.070000 358.500000 572.410000 ;
      RECT 1166.500000 572.065000 1183.980000 573.590000 ;
      RECT 1139.000000 571.590000 1158.500000 572.410000 ;
      RECT 372.500000 571.590000 389.000000 572.410000 ;
      RECT 0.000000 571.590000 358.500000 572.070000 ;
      RECT 1166.500000 570.410000 1186.000000 572.065000 ;
      RECT 1157.500000 570.410000 1158.500000 571.590000 ;
      RECT 372.500000 570.410000 373.500000 571.590000 ;
      RECT 357.500000 570.410000 358.500000 571.590000 ;
      RECT 1157.500000 569.590000 1186.000000 570.410000 ;
      RECT 357.500000 569.590000 373.500000 570.410000 ;
      RECT 1166.500000 569.485000 1186.000000 569.590000 ;
      RECT 1157.500000 568.410000 1158.500000 569.590000 ;
      RECT 1139.000000 568.410000 1149.500000 571.590000 ;
      RECT 386.500000 568.410000 389.000000 571.590000 ;
      RECT 372.500000 568.410000 373.500000 569.590000 ;
      RECT 357.500000 568.410000 358.500000 569.590000 ;
      RECT 0.000000 568.410000 349.500000 571.590000 ;
      RECT 1139.000000 567.590000 1158.500000 568.410000 ;
      RECT 372.500000 567.590000 389.000000 568.410000 ;
      RECT 0.000000 567.590000 358.500000 568.410000 ;
      RECT 1166.500000 566.410000 1183.980000 569.485000 ;
      RECT 1157.500000 566.410000 1158.500000 567.590000 ;
      RECT 372.500000 566.410000 373.500000 567.590000 ;
      RECT 357.500000 566.410000 358.500000 567.590000 ;
      RECT 1157.500000 566.385000 1183.980000 566.410000 ;
      RECT 1157.500000 565.590000 1186.000000 566.385000 ;
      RECT 357.500000 565.590000 373.500000 566.410000 ;
      RECT 1166.500000 565.525000 1186.000000 565.590000 ;
      RECT 0.000000 564.575000 349.500000 567.590000 ;
      RECT 1157.500000 564.410000 1158.500000 565.590000 ;
      RECT 1139.000000 564.410000 1149.500000 567.590000 ;
      RECT 386.500000 564.410000 389.000000 567.590000 ;
      RECT 372.500000 564.410000 373.500000 565.590000 ;
      RECT 357.500000 564.410000 358.500000 565.590000 ;
      RECT 2.020000 564.410000 349.500000 564.575000 ;
      RECT 1139.000000 563.590000 1158.500000 564.410000 ;
      RECT 372.500000 563.590000 389.000000 564.410000 ;
      RECT 2.020000 563.590000 358.500000 564.410000 ;
      RECT 1166.500000 562.425000 1183.980000 565.525000 ;
      RECT 1166.500000 562.410000 1186.000000 562.425000 ;
      RECT 1157.500000 562.410000 1158.500000 563.590000 ;
      RECT 372.500000 562.410000 373.500000 563.590000 ;
      RECT 357.500000 562.410000 358.500000 563.590000 ;
      RECT 1157.500000 561.590000 1186.000000 562.410000 ;
      RECT 357.500000 561.590000 373.500000 562.410000 ;
      RECT 2.020000 561.475000 349.500000 563.590000 ;
      RECT 0.000000 560.615000 349.500000 561.475000 ;
      RECT 1157.500000 560.410000 1158.500000 561.590000 ;
      RECT 1139.000000 560.410000 1149.500000 563.590000 ;
      RECT 386.500000 560.410000 389.000000 563.590000 ;
      RECT 372.500000 560.410000 373.500000 561.590000 ;
      RECT 357.500000 560.410000 358.500000 561.590000 ;
      RECT 2.020000 560.410000 349.500000 560.615000 ;
      RECT 1139.000000 559.590000 1158.500000 560.410000 ;
      RECT 372.500000 559.590000 389.000000 560.410000 ;
      RECT 2.020000 559.590000 358.500000 560.410000 ;
      RECT 1166.500000 558.410000 1186.000000 561.590000 ;
      RECT 1157.500000 558.410000 1158.500000 559.590000 ;
      RECT 372.500000 558.410000 373.500000 559.590000 ;
      RECT 357.500000 558.410000 358.500000 559.590000 ;
      RECT 1157.500000 557.590000 1186.000000 558.410000 ;
      RECT 357.500000 557.590000 373.500000 558.410000 ;
      RECT 2.020000 557.515000 349.500000 559.590000 ;
      RECT 1157.500000 556.410000 1158.500000 557.590000 ;
      RECT 1139.000000 556.410000 1149.500000 559.590000 ;
      RECT 386.500000 556.410000 389.000000 559.590000 ;
      RECT 372.500000 556.410000 373.500000 557.590000 ;
      RECT 357.500000 556.410000 358.500000 557.590000 ;
      RECT 0.000000 556.410000 349.500000 557.515000 ;
      RECT 1139.000000 555.590000 1158.500000 556.410000 ;
      RECT 372.500000 555.590000 389.000000 556.410000 ;
      RECT 0.000000 555.590000 358.500000 556.410000 ;
      RECT 0.000000 554.935000 349.500000 555.590000 ;
      RECT 1166.500000 554.930000 1186.000000 557.590000 ;
      RECT 1166.500000 554.410000 1183.980000 554.930000 ;
      RECT 1157.500000 554.410000 1158.500000 555.590000 ;
      RECT 372.500000 554.410000 373.500000 555.590000 ;
      RECT 357.500000 554.410000 358.500000 555.590000 ;
      RECT 1157.500000 553.590000 1183.980000 554.410000 ;
      RECT 357.500000 553.590000 373.500000 554.410000 ;
      RECT 1157.500000 552.410000 1158.500000 553.590000 ;
      RECT 1139.000000 552.410000 1149.500000 555.590000 ;
      RECT 386.500000 552.410000 389.000000 555.590000 ;
      RECT 372.500000 552.410000 373.500000 553.590000 ;
      RECT 357.500000 552.410000 358.500000 553.590000 ;
      RECT 2.020000 552.410000 349.500000 554.935000 ;
      RECT 2.020000 551.835000 358.500000 552.410000 ;
      RECT 1166.500000 551.830000 1183.980000 553.590000 ;
      RECT 1139.000000 551.590000 1158.500000 552.410000 ;
      RECT 372.500000 551.590000 389.000000 552.410000 ;
      RECT 0.000000 551.590000 358.500000 551.835000 ;
      RECT 1166.500000 550.410000 1186.000000 551.830000 ;
      RECT 1157.500000 550.410000 1158.500000 551.590000 ;
      RECT 372.500000 550.410000 373.500000 551.590000 ;
      RECT 357.500000 550.410000 358.500000 551.590000 ;
      RECT 1157.500000 549.590000 1186.000000 550.410000 ;
      RECT 357.500000 549.590000 373.500000 550.410000 ;
      RECT 1157.500000 548.410000 1158.500000 549.590000 ;
      RECT 1139.000000 548.410000 1149.500000 551.590000 ;
      RECT 386.500000 548.410000 389.000000 551.590000 ;
      RECT 372.500000 548.410000 373.500000 549.590000 ;
      RECT 357.500000 548.410000 358.500000 549.590000 ;
      RECT 0.000000 548.410000 349.500000 551.590000 ;
      RECT 1139.000000 547.590000 1158.500000 548.410000 ;
      RECT 372.500000 547.590000 389.000000 548.410000 ;
      RECT 0.000000 547.590000 358.500000 548.410000 ;
      RECT 1166.500000 546.410000 1186.000000 549.590000 ;
      RECT 1157.500000 546.410000 1158.500000 547.590000 ;
      RECT 372.500000 546.410000 373.500000 547.590000 ;
      RECT 357.500000 546.410000 358.500000 547.590000 ;
      RECT 1157.500000 545.590000 1186.000000 546.410000 ;
      RECT 357.500000 545.590000 373.500000 546.410000 ;
      RECT 1157.500000 544.410000 1158.500000 545.590000 ;
      RECT 1139.000000 544.410000 1149.500000 547.590000 ;
      RECT 386.500000 544.410000 389.000000 547.590000 ;
      RECT 372.500000 544.410000 373.500000 545.590000 ;
      RECT 357.500000 544.410000 358.500000 545.590000 ;
      RECT 0.000000 544.410000 349.500000 547.590000 ;
      RECT 1139.000000 543.590000 1158.500000 544.410000 ;
      RECT 372.500000 543.590000 389.000000 544.410000 ;
      RECT 0.000000 543.590000 358.500000 544.410000 ;
      RECT 1166.500000 542.410000 1186.000000 545.590000 ;
      RECT 1157.500000 542.410000 1158.500000 543.590000 ;
      RECT 372.500000 542.410000 373.500000 543.590000 ;
      RECT 357.500000 542.410000 358.500000 543.590000 ;
      RECT 1157.500000 541.590000 1186.000000 542.410000 ;
      RECT 357.500000 541.590000 373.500000 542.410000 ;
      RECT 1157.500000 540.410000 1158.500000 541.590000 ;
      RECT 1139.000000 540.410000 1149.500000 543.590000 ;
      RECT 386.500000 540.410000 389.000000 543.590000 ;
      RECT 372.500000 540.410000 373.500000 541.590000 ;
      RECT 357.500000 540.410000 358.500000 541.590000 ;
      RECT 0.000000 540.410000 349.500000 543.590000 ;
      RECT 1139.000000 539.590000 1158.500000 540.410000 ;
      RECT 372.500000 539.590000 389.000000 540.410000 ;
      RECT 0.000000 539.590000 358.500000 540.410000 ;
      RECT 1166.500000 538.410000 1186.000000 541.590000 ;
      RECT 1157.500000 538.410000 1158.500000 539.590000 ;
      RECT 372.500000 538.410000 373.500000 539.590000 ;
      RECT 357.500000 538.410000 358.500000 539.590000 ;
      RECT 1157.500000 537.590000 1186.000000 538.410000 ;
      RECT 357.500000 537.590000 373.500000 538.410000 ;
      RECT 1157.500000 536.410000 1158.500000 537.590000 ;
      RECT 1139.000000 536.410000 1149.500000 539.590000 ;
      RECT 386.500000 536.410000 389.000000 539.590000 ;
      RECT 372.500000 536.410000 373.500000 537.590000 ;
      RECT 357.500000 536.410000 358.500000 537.590000 ;
      RECT 0.000000 536.410000 349.500000 539.590000 ;
      RECT 1139.000000 535.590000 1158.500000 536.410000 ;
      RECT 372.500000 535.590000 389.000000 536.410000 ;
      RECT 0.000000 535.590000 358.500000 536.410000 ;
      RECT 1166.500000 534.410000 1186.000000 537.590000 ;
      RECT 1157.500000 534.410000 1158.500000 535.590000 ;
      RECT 372.500000 534.410000 373.500000 535.590000 ;
      RECT 357.500000 534.410000 358.500000 535.590000 ;
      RECT 1157.500000 533.590000 1186.000000 534.410000 ;
      RECT 357.500000 533.590000 373.500000 534.410000 ;
      RECT 1157.500000 532.410000 1158.500000 533.590000 ;
      RECT 1139.000000 532.410000 1149.500000 535.590000 ;
      RECT 386.500000 532.410000 389.000000 535.590000 ;
      RECT 372.500000 532.410000 373.500000 533.590000 ;
      RECT 357.500000 532.410000 358.500000 533.590000 ;
      RECT 0.000000 532.410000 349.500000 535.590000 ;
      RECT 1139.000000 531.590000 1158.500000 532.410000 ;
      RECT 372.500000 531.590000 389.000000 532.410000 ;
      RECT 0.000000 531.590000 358.500000 532.410000 ;
      RECT 1166.500000 530.410000 1186.000000 533.590000 ;
      RECT 1157.500000 530.410000 1158.500000 531.590000 ;
      RECT 372.500000 530.410000 373.500000 531.590000 ;
      RECT 357.500000 530.410000 358.500000 531.590000 ;
      RECT 1157.500000 529.590000 1186.000000 530.410000 ;
      RECT 357.500000 529.590000 373.500000 530.410000 ;
      RECT 1157.500000 528.410000 1158.500000 529.590000 ;
      RECT 1139.000000 528.410000 1149.500000 531.590000 ;
      RECT 386.500000 528.410000 389.000000 531.590000 ;
      RECT 372.500000 528.410000 373.500000 529.590000 ;
      RECT 357.500000 528.410000 358.500000 529.590000 ;
      RECT 0.000000 528.410000 349.500000 531.590000 ;
      RECT 1139.000000 527.590000 1158.500000 528.410000 ;
      RECT 372.500000 527.590000 389.000000 528.410000 ;
      RECT 0.000000 527.590000 358.500000 528.410000 ;
      RECT 1166.500000 526.410000 1186.000000 529.590000 ;
      RECT 1157.500000 526.410000 1158.500000 527.590000 ;
      RECT 372.500000 526.410000 373.500000 527.590000 ;
      RECT 357.500000 526.410000 358.500000 527.590000 ;
      RECT 1157.500000 525.590000 1186.000000 526.410000 ;
      RECT 357.500000 525.590000 373.500000 526.410000 ;
      RECT 1157.500000 524.410000 1158.500000 525.590000 ;
      RECT 1139.000000 524.410000 1149.500000 527.590000 ;
      RECT 386.500000 524.410000 389.000000 527.590000 ;
      RECT 372.500000 524.410000 373.500000 525.590000 ;
      RECT 357.500000 524.410000 358.500000 525.590000 ;
      RECT 0.000000 524.410000 349.500000 527.590000 ;
      RECT 1139.000000 523.590000 1158.500000 524.410000 ;
      RECT 372.500000 523.590000 389.000000 524.410000 ;
      RECT 0.000000 523.590000 358.500000 524.410000 ;
      RECT 1166.500000 522.410000 1186.000000 525.590000 ;
      RECT 1157.500000 522.410000 1158.500000 523.590000 ;
      RECT 372.500000 522.410000 373.500000 523.590000 ;
      RECT 357.500000 522.410000 358.500000 523.590000 ;
      RECT 1157.500000 521.590000 1186.000000 522.410000 ;
      RECT 357.500000 521.590000 373.500000 522.410000 ;
      RECT 1157.500000 520.410000 1158.500000 521.590000 ;
      RECT 1139.000000 520.410000 1149.500000 523.590000 ;
      RECT 386.500000 520.410000 389.000000 523.590000 ;
      RECT 372.500000 520.410000 373.500000 521.590000 ;
      RECT 357.500000 520.410000 358.500000 521.590000 ;
      RECT 0.000000 520.410000 349.500000 523.590000 ;
      RECT 1139.000000 519.590000 1158.500000 520.410000 ;
      RECT 372.500000 519.590000 389.000000 520.410000 ;
      RECT 0.000000 519.590000 358.500000 520.410000 ;
      RECT 1166.500000 518.410000 1186.000000 521.590000 ;
      RECT 1157.500000 518.410000 1158.500000 519.590000 ;
      RECT 372.500000 518.410000 373.500000 519.590000 ;
      RECT 357.500000 518.410000 358.500000 519.590000 ;
      RECT 1157.500000 517.590000 1186.000000 518.410000 ;
      RECT 357.500000 517.590000 373.500000 518.410000 ;
      RECT 307.500000 517.590000 349.500000 519.590000 ;
      RECT 0.000000 517.590000 299.500000 519.590000 ;
      RECT 1157.500000 516.410000 1158.500000 517.590000 ;
      RECT 1139.000000 516.410000 1149.500000 519.590000 ;
      RECT 386.500000 516.410000 389.000000 519.590000 ;
      RECT 372.500000 516.410000 373.500000 517.590000 ;
      RECT 357.500000 516.410000 358.500000 517.590000 ;
      RECT 316.500000 516.410000 349.500000 517.590000 ;
      RECT 307.500000 516.410000 308.500000 517.590000 ;
      RECT 266.500000 516.410000 299.500000 517.590000 ;
      RECT 1139.000000 515.590000 1158.500000 516.410000 ;
      RECT 372.500000 515.590000 389.000000 516.410000 ;
      RECT 316.500000 515.590000 358.500000 516.410000 ;
      RECT 266.500000 515.590000 308.500000 516.410000 ;
      RECT 216.500000 515.590000 258.500000 517.590000 ;
      RECT 166.500000 515.590000 208.500000 517.590000 ;
      RECT 116.500000 515.590000 158.500000 517.590000 ;
      RECT 66.500000 515.590000 108.500000 517.590000 ;
      RECT 29.500000 515.590000 58.500000 517.590000 ;
      RECT 0.000000 515.590000 16.500000 517.590000 ;
      RECT 1166.500000 514.410000 1186.000000 517.590000 ;
      RECT 1157.500000 514.410000 1158.500000 515.590000 ;
      RECT 372.500000 514.410000 373.500000 515.590000 ;
      RECT 357.500000 514.410000 358.500000 515.590000 ;
      RECT 316.500000 514.410000 349.500000 515.590000 ;
      RECT 307.500000 514.410000 308.500000 515.590000 ;
      RECT 266.500000 514.410000 299.500000 515.590000 ;
      RECT 257.500000 514.410000 258.500000 515.590000 ;
      RECT 216.500000 514.410000 249.500000 515.590000 ;
      RECT 207.500000 514.410000 208.500000 515.590000 ;
      RECT 166.500000 514.410000 199.500000 515.590000 ;
      RECT 157.500000 514.410000 158.500000 515.590000 ;
      RECT 116.500000 514.410000 149.500000 515.590000 ;
      RECT 107.500000 514.410000 108.500000 515.590000 ;
      RECT 66.500000 514.410000 99.500000 515.590000 ;
      RECT 57.500000 514.410000 58.500000 515.590000 ;
      RECT 29.500000 514.410000 49.500000 515.590000 ;
      RECT 15.500000 514.410000 16.500000 515.590000 ;
      RECT 1157.500000 513.590000 1186.000000 514.410000 ;
      RECT 357.500000 513.590000 373.500000 514.410000 ;
      RECT 307.500000 513.590000 349.500000 514.410000 ;
      RECT 257.500000 513.590000 299.500000 514.410000 ;
      RECT 207.500000 513.590000 249.500000 514.410000 ;
      RECT 157.500000 513.590000 199.500000 514.410000 ;
      RECT 107.500000 513.590000 149.500000 514.410000 ;
      RECT 57.500000 513.590000 99.500000 514.410000 ;
      RECT 15.500000 513.590000 49.500000 514.410000 ;
      RECT 1157.500000 512.410000 1158.500000 513.590000 ;
      RECT 1139.000000 512.410000 1149.500000 515.590000 ;
      RECT 386.500000 512.410000 389.000000 515.590000 ;
      RECT 372.500000 512.410000 373.500000 513.590000 ;
      RECT 357.500000 512.410000 358.500000 513.590000 ;
      RECT 316.500000 512.410000 349.500000 513.590000 ;
      RECT 307.500000 512.410000 308.500000 513.590000 ;
      RECT 266.500000 512.410000 299.500000 513.590000 ;
      RECT 257.500000 512.410000 258.500000 513.590000 ;
      RECT 216.500000 512.410000 249.500000 513.590000 ;
      RECT 207.500000 512.410000 208.500000 513.590000 ;
      RECT 166.500000 512.410000 199.500000 513.590000 ;
      RECT 157.500000 512.410000 158.500000 513.590000 ;
      RECT 116.500000 512.410000 149.500000 513.590000 ;
      RECT 107.500000 512.410000 108.500000 513.590000 ;
      RECT 66.500000 512.410000 99.500000 513.590000 ;
      RECT 57.500000 512.410000 58.500000 513.590000 ;
      RECT 29.500000 512.410000 49.500000 513.590000 ;
      RECT 15.500000 512.410000 16.500000 513.590000 ;
      RECT 0.000000 512.410000 2.500000 515.590000 ;
      RECT 1139.000000 511.590000 1158.500000 512.410000 ;
      RECT 372.500000 511.590000 389.000000 512.410000 ;
      RECT 316.500000 511.590000 358.500000 512.410000 ;
      RECT 266.500000 511.590000 308.500000 512.410000 ;
      RECT 216.500000 511.590000 258.500000 512.410000 ;
      RECT 166.500000 511.590000 208.500000 512.410000 ;
      RECT 116.500000 511.590000 158.500000 512.410000 ;
      RECT 66.500000 511.590000 108.500000 512.410000 ;
      RECT 29.500000 511.590000 58.500000 512.410000 ;
      RECT 0.000000 511.590000 16.500000 512.410000 ;
      RECT 1166.500000 510.410000 1186.000000 513.590000 ;
      RECT 1157.500000 510.410000 1158.500000 511.590000 ;
      RECT 372.500000 510.410000 373.500000 511.590000 ;
      RECT 357.500000 510.410000 358.500000 511.590000 ;
      RECT 316.500000 510.410000 349.500000 511.590000 ;
      RECT 307.500000 510.410000 308.500000 511.590000 ;
      RECT 266.500000 510.410000 299.500000 511.590000 ;
      RECT 257.500000 510.410000 258.500000 511.590000 ;
      RECT 216.500000 510.410000 249.500000 511.590000 ;
      RECT 207.500000 510.410000 208.500000 511.590000 ;
      RECT 166.500000 510.410000 199.500000 511.590000 ;
      RECT 157.500000 510.410000 158.500000 511.590000 ;
      RECT 116.500000 510.410000 149.500000 511.590000 ;
      RECT 107.500000 510.410000 108.500000 511.590000 ;
      RECT 66.500000 510.410000 99.500000 511.590000 ;
      RECT 57.500000 510.410000 58.500000 511.590000 ;
      RECT 29.500000 510.410000 49.500000 511.590000 ;
      RECT 15.500000 510.410000 16.500000 511.590000 ;
      RECT 1157.500000 509.590000 1186.000000 510.410000 ;
      RECT 357.500000 509.590000 373.500000 510.410000 ;
      RECT 307.500000 509.590000 349.500000 510.410000 ;
      RECT 257.500000 509.590000 299.500000 510.410000 ;
      RECT 207.500000 509.590000 249.500000 510.410000 ;
      RECT 157.500000 509.590000 199.500000 510.410000 ;
      RECT 107.500000 509.590000 149.500000 510.410000 ;
      RECT 57.500000 509.590000 99.500000 510.410000 ;
      RECT 15.500000 509.590000 49.500000 510.410000 ;
      RECT 1157.500000 508.410000 1158.500000 509.590000 ;
      RECT 1139.000000 508.410000 1149.500000 511.590000 ;
      RECT 386.500000 508.410000 389.000000 511.590000 ;
      RECT 372.500000 508.410000 373.500000 509.590000 ;
      RECT 357.500000 508.410000 358.500000 509.590000 ;
      RECT 316.500000 508.410000 349.500000 509.590000 ;
      RECT 307.500000 508.410000 308.500000 509.590000 ;
      RECT 266.500000 508.410000 299.500000 509.590000 ;
      RECT 257.500000 508.410000 258.500000 509.590000 ;
      RECT 216.500000 508.410000 249.500000 509.590000 ;
      RECT 207.500000 508.410000 208.500000 509.590000 ;
      RECT 166.500000 508.410000 199.500000 509.590000 ;
      RECT 157.500000 508.410000 158.500000 509.590000 ;
      RECT 116.500000 508.410000 149.500000 509.590000 ;
      RECT 107.500000 508.410000 108.500000 509.590000 ;
      RECT 66.500000 508.410000 99.500000 509.590000 ;
      RECT 57.500000 508.410000 58.500000 509.590000 ;
      RECT 29.500000 508.410000 49.500000 509.590000 ;
      RECT 15.500000 508.410000 16.500000 509.590000 ;
      RECT 0.000000 508.410000 2.500000 511.590000 ;
      RECT 1139.000000 507.590000 1158.500000 508.410000 ;
      RECT 372.500000 507.590000 389.000000 508.410000 ;
      RECT 316.500000 507.590000 358.500000 508.410000 ;
      RECT 266.500000 507.590000 308.500000 508.410000 ;
      RECT 216.500000 507.590000 258.500000 508.410000 ;
      RECT 166.500000 507.590000 208.500000 508.410000 ;
      RECT 116.500000 507.590000 158.500000 508.410000 ;
      RECT 66.500000 507.590000 108.500000 508.410000 ;
      RECT 29.500000 507.590000 58.500000 508.410000 ;
      RECT 0.000000 507.590000 16.500000 508.410000 ;
      RECT 1166.500000 506.410000 1186.000000 509.590000 ;
      RECT 1157.500000 506.410000 1158.500000 507.590000 ;
      RECT 372.500000 506.410000 373.500000 507.590000 ;
      RECT 357.500000 506.410000 358.500000 507.590000 ;
      RECT 316.500000 506.410000 349.500000 507.590000 ;
      RECT 307.500000 506.410000 308.500000 507.590000 ;
      RECT 266.500000 506.410000 299.500000 507.590000 ;
      RECT 257.500000 506.410000 258.500000 507.590000 ;
      RECT 216.500000 506.410000 249.500000 507.590000 ;
      RECT 207.500000 506.410000 208.500000 507.590000 ;
      RECT 166.500000 506.410000 199.500000 507.590000 ;
      RECT 157.500000 506.410000 158.500000 507.590000 ;
      RECT 116.500000 506.410000 149.500000 507.590000 ;
      RECT 107.500000 506.410000 108.500000 507.590000 ;
      RECT 66.500000 506.410000 99.500000 507.590000 ;
      RECT 57.500000 506.410000 58.500000 507.590000 ;
      RECT 29.500000 506.410000 49.500000 507.590000 ;
      RECT 15.500000 506.410000 16.500000 507.590000 ;
      RECT 386.500000 506.000000 389.000000 507.590000 ;
      RECT 1157.500000 505.590000 1186.000000 506.410000 ;
      RECT 386.500000 505.590000 739.000000 506.000000 ;
      RECT 357.500000 505.590000 373.500000 506.410000 ;
      RECT 307.500000 505.590000 349.500000 506.410000 ;
      RECT 257.500000 505.590000 299.500000 506.410000 ;
      RECT 207.500000 505.590000 249.500000 506.410000 ;
      RECT 157.500000 505.590000 199.500000 506.410000 ;
      RECT 107.500000 505.590000 149.500000 506.410000 ;
      RECT 57.500000 505.590000 99.500000 506.410000 ;
      RECT 15.500000 505.590000 49.500000 506.410000 ;
      RECT 1157.500000 504.410000 1158.500000 505.590000 ;
      RECT 1139.000000 504.410000 1149.500000 507.590000 ;
      RECT 386.500000 504.410000 408.500000 505.590000 ;
      RECT 372.500000 504.410000 373.500000 505.590000 ;
      RECT 357.500000 504.410000 358.500000 505.590000 ;
      RECT 316.500000 504.410000 349.500000 505.590000 ;
      RECT 307.500000 504.410000 308.500000 505.590000 ;
      RECT 266.500000 504.410000 299.500000 505.590000 ;
      RECT 257.500000 504.410000 258.500000 505.590000 ;
      RECT 216.500000 504.410000 249.500000 505.590000 ;
      RECT 207.500000 504.410000 208.500000 505.590000 ;
      RECT 166.500000 504.410000 199.500000 505.590000 ;
      RECT 157.500000 504.410000 158.500000 505.590000 ;
      RECT 116.500000 504.410000 149.500000 505.590000 ;
      RECT 107.500000 504.410000 108.500000 505.590000 ;
      RECT 66.500000 504.410000 99.500000 505.590000 ;
      RECT 57.500000 504.410000 58.500000 505.590000 ;
      RECT 29.500000 504.410000 49.500000 505.590000 ;
      RECT 15.500000 504.410000 16.500000 505.590000 ;
      RECT 0.000000 504.410000 2.500000 507.590000 ;
      RECT 1139.000000 503.590000 1158.500000 504.410000 ;
      RECT 716.500000 503.590000 739.000000 505.590000 ;
      RECT 666.500000 503.590000 708.500000 505.590000 ;
      RECT 616.500000 503.590000 658.500000 505.590000 ;
      RECT 566.500000 503.590000 608.500000 505.590000 ;
      RECT 516.500000 503.590000 558.500000 505.590000 ;
      RECT 466.500000 503.590000 508.500000 505.590000 ;
      RECT 416.500000 503.590000 458.500000 505.590000 ;
      RECT 372.500000 503.590000 408.500000 504.410000 ;
      RECT 316.500000 503.590000 358.500000 504.410000 ;
      RECT 266.500000 503.590000 308.500000 504.410000 ;
      RECT 216.500000 503.590000 258.500000 504.410000 ;
      RECT 166.500000 503.590000 208.500000 504.410000 ;
      RECT 116.500000 503.590000 158.500000 504.410000 ;
      RECT 66.500000 503.590000 108.500000 504.410000 ;
      RECT 29.500000 503.590000 58.500000 504.410000 ;
      RECT 0.000000 503.590000 16.500000 504.410000 ;
      RECT 1166.500000 502.410000 1186.000000 505.590000 ;
      RECT 1157.500000 502.410000 1158.500000 503.590000 ;
      RECT 716.500000 502.410000 723.500000 503.590000 ;
      RECT 707.500000 502.410000 708.500000 503.590000 ;
      RECT 666.500000 502.410000 699.500000 503.590000 ;
      RECT 657.500000 502.410000 658.500000 503.590000 ;
      RECT 616.500000 502.410000 649.500000 503.590000 ;
      RECT 607.500000 502.410000 608.500000 503.590000 ;
      RECT 566.500000 502.410000 599.500000 503.590000 ;
      RECT 557.500000 502.410000 558.500000 503.590000 ;
      RECT 516.500000 502.410000 549.500000 503.590000 ;
      RECT 507.500000 502.410000 508.500000 503.590000 ;
      RECT 466.500000 502.410000 499.500000 503.590000 ;
      RECT 457.500000 502.410000 458.500000 503.590000 ;
      RECT 416.500000 502.410000 449.500000 503.590000 ;
      RECT 407.500000 502.410000 408.500000 503.590000 ;
      RECT 372.500000 502.410000 373.500000 503.590000 ;
      RECT 357.500000 502.410000 358.500000 503.590000 ;
      RECT 316.500000 502.410000 349.500000 503.590000 ;
      RECT 307.500000 502.410000 308.500000 503.590000 ;
      RECT 266.500000 502.410000 299.500000 503.590000 ;
      RECT 257.500000 502.410000 258.500000 503.590000 ;
      RECT 216.500000 502.410000 249.500000 503.590000 ;
      RECT 207.500000 502.410000 208.500000 503.590000 ;
      RECT 166.500000 502.410000 199.500000 503.590000 ;
      RECT 157.500000 502.410000 158.500000 503.590000 ;
      RECT 116.500000 502.410000 149.500000 503.590000 ;
      RECT 107.500000 502.410000 108.500000 503.590000 ;
      RECT 66.500000 502.410000 99.500000 503.590000 ;
      RECT 57.500000 502.410000 58.500000 503.590000 ;
      RECT 29.500000 502.410000 49.500000 503.590000 ;
      RECT 15.500000 502.410000 16.500000 503.590000 ;
      RECT 1157.500000 501.590000 1186.000000 502.410000 ;
      RECT 707.500000 501.590000 723.500000 502.410000 ;
      RECT 657.500000 501.590000 699.500000 502.410000 ;
      RECT 607.500000 501.590000 649.500000 502.410000 ;
      RECT 557.500000 501.590000 599.500000 502.410000 ;
      RECT 507.500000 501.590000 549.500000 502.410000 ;
      RECT 457.500000 501.590000 499.500000 502.410000 ;
      RECT 407.500000 501.590000 449.500000 502.410000 ;
      RECT 357.500000 501.590000 373.500000 502.410000 ;
      RECT 307.500000 501.590000 349.500000 502.410000 ;
      RECT 257.500000 501.590000 299.500000 502.410000 ;
      RECT 207.500000 501.590000 249.500000 502.410000 ;
      RECT 157.500000 501.590000 199.500000 502.410000 ;
      RECT 107.500000 501.590000 149.500000 502.410000 ;
      RECT 57.500000 501.590000 99.500000 502.410000 ;
      RECT 15.500000 501.590000 49.500000 502.410000 ;
      RECT 1157.500000 500.410000 1158.500000 501.590000 ;
      RECT 1139.000000 500.410000 1149.500000 503.590000 ;
      RECT 736.500000 500.410000 739.000000 503.590000 ;
      RECT 716.500000 500.410000 723.500000 501.590000 ;
      RECT 707.500000 500.410000 708.500000 501.590000 ;
      RECT 666.500000 500.410000 699.500000 501.590000 ;
      RECT 657.500000 500.410000 658.500000 501.590000 ;
      RECT 616.500000 500.410000 649.500000 501.590000 ;
      RECT 607.500000 500.410000 608.500000 501.590000 ;
      RECT 566.500000 500.410000 599.500000 501.590000 ;
      RECT 557.500000 500.410000 558.500000 501.590000 ;
      RECT 516.500000 500.410000 549.500000 501.590000 ;
      RECT 507.500000 500.410000 508.500000 501.590000 ;
      RECT 466.500000 500.410000 499.500000 501.590000 ;
      RECT 457.500000 500.410000 458.500000 501.590000 ;
      RECT 416.500000 500.410000 449.500000 501.590000 ;
      RECT 407.500000 500.410000 408.500000 501.590000 ;
      RECT 386.500000 500.410000 399.500000 503.590000 ;
      RECT 372.500000 500.410000 373.500000 501.590000 ;
      RECT 357.500000 500.410000 358.500000 501.590000 ;
      RECT 316.500000 500.410000 349.500000 501.590000 ;
      RECT 307.500000 500.410000 308.500000 501.590000 ;
      RECT 266.500000 500.410000 299.500000 501.590000 ;
      RECT 257.500000 500.410000 258.500000 501.590000 ;
      RECT 216.500000 500.410000 249.500000 501.590000 ;
      RECT 207.500000 500.410000 208.500000 501.590000 ;
      RECT 166.500000 500.410000 199.500000 501.590000 ;
      RECT 157.500000 500.410000 158.500000 501.590000 ;
      RECT 116.500000 500.410000 149.500000 501.590000 ;
      RECT 107.500000 500.410000 108.500000 501.590000 ;
      RECT 66.500000 500.410000 99.500000 501.590000 ;
      RECT 57.500000 500.410000 58.500000 501.590000 ;
      RECT 29.500000 500.410000 49.500000 501.590000 ;
      RECT 15.500000 500.410000 16.500000 501.590000 ;
      RECT 0.000000 500.410000 2.500000 503.590000 ;
      RECT 1139.000000 499.590000 1158.500000 500.410000 ;
      RECT 716.500000 499.590000 739.000000 500.410000 ;
      RECT 666.500000 499.590000 708.500000 500.410000 ;
      RECT 616.500000 499.590000 658.500000 500.410000 ;
      RECT 566.500000 499.590000 608.500000 500.410000 ;
      RECT 516.500000 499.590000 558.500000 500.410000 ;
      RECT 466.500000 499.590000 508.500000 500.410000 ;
      RECT 416.500000 499.590000 458.500000 500.410000 ;
      RECT 372.500000 499.590000 408.500000 500.410000 ;
      RECT 316.500000 499.590000 358.500000 500.410000 ;
      RECT 266.500000 499.590000 308.500000 500.410000 ;
      RECT 216.500000 499.590000 258.500000 500.410000 ;
      RECT 166.500000 499.590000 208.500000 500.410000 ;
      RECT 116.500000 499.590000 158.500000 500.410000 ;
      RECT 66.500000 499.590000 108.500000 500.410000 ;
      RECT 29.500000 499.590000 58.500000 500.410000 ;
      RECT 0.000000 499.590000 16.500000 500.410000 ;
      RECT 1166.500000 498.410000 1186.000000 501.590000 ;
      RECT 1157.500000 498.410000 1158.500000 499.590000 ;
      RECT 716.500000 498.410000 723.500000 499.590000 ;
      RECT 707.500000 498.410000 708.500000 499.590000 ;
      RECT 666.500000 498.410000 699.500000 499.590000 ;
      RECT 657.500000 498.410000 658.500000 499.590000 ;
      RECT 616.500000 498.410000 649.500000 499.590000 ;
      RECT 607.500000 498.410000 608.500000 499.590000 ;
      RECT 566.500000 498.410000 599.500000 499.590000 ;
      RECT 557.500000 498.410000 558.500000 499.590000 ;
      RECT 516.500000 498.410000 549.500000 499.590000 ;
      RECT 507.500000 498.410000 508.500000 499.590000 ;
      RECT 466.500000 498.410000 499.500000 499.590000 ;
      RECT 457.500000 498.410000 458.500000 499.590000 ;
      RECT 416.500000 498.410000 449.500000 499.590000 ;
      RECT 407.500000 498.410000 408.500000 499.590000 ;
      RECT 372.500000 498.410000 373.500000 499.590000 ;
      RECT 357.500000 498.410000 358.500000 499.590000 ;
      RECT 316.500000 498.410000 349.500000 499.590000 ;
      RECT 307.500000 498.410000 308.500000 499.590000 ;
      RECT 266.500000 498.410000 299.500000 499.590000 ;
      RECT 257.500000 498.410000 258.500000 499.590000 ;
      RECT 216.500000 498.410000 249.500000 499.590000 ;
      RECT 207.500000 498.410000 208.500000 499.590000 ;
      RECT 166.500000 498.410000 199.500000 499.590000 ;
      RECT 157.500000 498.410000 158.500000 499.590000 ;
      RECT 116.500000 498.410000 149.500000 499.590000 ;
      RECT 107.500000 498.410000 108.500000 499.590000 ;
      RECT 66.500000 498.410000 99.500000 499.590000 ;
      RECT 57.500000 498.410000 58.500000 499.590000 ;
      RECT 29.500000 498.410000 49.500000 499.590000 ;
      RECT 15.500000 498.410000 16.500000 499.590000 ;
      RECT 1157.500000 497.590000 1186.000000 498.410000 ;
      RECT 707.500000 497.590000 723.500000 498.410000 ;
      RECT 657.500000 497.590000 699.500000 498.410000 ;
      RECT 607.500000 497.590000 649.500000 498.410000 ;
      RECT 557.500000 497.590000 599.500000 498.410000 ;
      RECT 507.500000 497.590000 549.500000 498.410000 ;
      RECT 457.500000 497.590000 499.500000 498.410000 ;
      RECT 407.500000 497.590000 449.500000 498.410000 ;
      RECT 357.500000 497.590000 373.500000 498.410000 ;
      RECT 307.500000 497.590000 349.500000 498.410000 ;
      RECT 257.500000 497.590000 299.500000 498.410000 ;
      RECT 207.500000 497.590000 249.500000 498.410000 ;
      RECT 157.500000 497.590000 199.500000 498.410000 ;
      RECT 107.500000 497.590000 149.500000 498.410000 ;
      RECT 57.500000 497.590000 99.500000 498.410000 ;
      RECT 15.500000 497.590000 49.500000 498.410000 ;
      RECT 1157.500000 496.410000 1158.500000 497.590000 ;
      RECT 1139.000000 496.410000 1149.500000 499.590000 ;
      RECT 736.500000 496.410000 739.000000 499.590000 ;
      RECT 716.500000 496.410000 723.500000 497.590000 ;
      RECT 707.500000 496.410000 708.500000 497.590000 ;
      RECT 666.500000 496.410000 699.500000 497.590000 ;
      RECT 657.500000 496.410000 658.500000 497.590000 ;
      RECT 616.500000 496.410000 649.500000 497.590000 ;
      RECT 607.500000 496.410000 608.500000 497.590000 ;
      RECT 566.500000 496.410000 599.500000 497.590000 ;
      RECT 557.500000 496.410000 558.500000 497.590000 ;
      RECT 516.500000 496.410000 549.500000 497.590000 ;
      RECT 507.500000 496.410000 508.500000 497.590000 ;
      RECT 466.500000 496.410000 499.500000 497.590000 ;
      RECT 457.500000 496.410000 458.500000 497.590000 ;
      RECT 416.500000 496.410000 449.500000 497.590000 ;
      RECT 407.500000 496.410000 408.500000 497.590000 ;
      RECT 386.500000 496.410000 399.500000 499.590000 ;
      RECT 372.500000 496.410000 373.500000 497.590000 ;
      RECT 357.500000 496.410000 358.500000 497.590000 ;
      RECT 316.500000 496.410000 349.500000 497.590000 ;
      RECT 307.500000 496.410000 308.500000 497.590000 ;
      RECT 266.500000 496.410000 299.500000 497.590000 ;
      RECT 257.500000 496.410000 258.500000 497.590000 ;
      RECT 216.500000 496.410000 249.500000 497.590000 ;
      RECT 207.500000 496.410000 208.500000 497.590000 ;
      RECT 166.500000 496.410000 199.500000 497.590000 ;
      RECT 157.500000 496.410000 158.500000 497.590000 ;
      RECT 116.500000 496.410000 149.500000 497.590000 ;
      RECT 107.500000 496.410000 108.500000 497.590000 ;
      RECT 66.500000 496.410000 99.500000 497.590000 ;
      RECT 57.500000 496.410000 58.500000 497.590000 ;
      RECT 29.500000 496.410000 49.500000 497.590000 ;
      RECT 15.500000 496.410000 16.500000 497.590000 ;
      RECT 0.000000 496.410000 2.500000 499.590000 ;
      RECT 1139.000000 495.590000 1158.500000 496.410000 ;
      RECT 716.500000 495.590000 739.000000 496.410000 ;
      RECT 666.500000 495.590000 708.500000 496.410000 ;
      RECT 616.500000 495.590000 658.500000 496.410000 ;
      RECT 566.500000 495.590000 608.500000 496.410000 ;
      RECT 516.500000 495.590000 558.500000 496.410000 ;
      RECT 466.500000 495.590000 508.500000 496.410000 ;
      RECT 416.500000 495.590000 458.500000 496.410000 ;
      RECT 372.500000 495.590000 408.500000 496.410000 ;
      RECT 316.500000 495.590000 358.500000 496.410000 ;
      RECT 266.500000 495.590000 308.500000 496.410000 ;
      RECT 216.500000 495.590000 258.500000 496.410000 ;
      RECT 166.500000 495.590000 208.500000 496.410000 ;
      RECT 116.500000 495.590000 158.500000 496.410000 ;
      RECT 66.500000 495.590000 108.500000 496.410000 ;
      RECT 29.500000 495.590000 58.500000 496.410000 ;
      RECT 0.000000 495.590000 16.500000 496.410000 ;
      RECT 1166.500000 494.410000 1186.000000 497.590000 ;
      RECT 1157.500000 494.410000 1158.500000 495.590000 ;
      RECT 716.500000 494.410000 723.500000 495.590000 ;
      RECT 707.500000 494.410000 708.500000 495.590000 ;
      RECT 666.500000 494.410000 699.500000 495.590000 ;
      RECT 657.500000 494.410000 658.500000 495.590000 ;
      RECT 616.500000 494.410000 649.500000 495.590000 ;
      RECT 607.500000 494.410000 608.500000 495.590000 ;
      RECT 566.500000 494.410000 599.500000 495.590000 ;
      RECT 557.500000 494.410000 558.500000 495.590000 ;
      RECT 516.500000 494.410000 549.500000 495.590000 ;
      RECT 507.500000 494.410000 508.500000 495.590000 ;
      RECT 466.500000 494.410000 499.500000 495.590000 ;
      RECT 457.500000 494.410000 458.500000 495.590000 ;
      RECT 416.500000 494.410000 449.500000 495.590000 ;
      RECT 407.500000 494.410000 408.500000 495.590000 ;
      RECT 372.500000 494.410000 373.500000 495.590000 ;
      RECT 357.500000 494.410000 358.500000 495.590000 ;
      RECT 316.500000 494.410000 349.500000 495.590000 ;
      RECT 307.500000 494.410000 308.500000 495.590000 ;
      RECT 266.500000 494.410000 299.500000 495.590000 ;
      RECT 257.500000 494.410000 258.500000 495.590000 ;
      RECT 216.500000 494.410000 249.500000 495.590000 ;
      RECT 207.500000 494.410000 208.500000 495.590000 ;
      RECT 166.500000 494.410000 199.500000 495.590000 ;
      RECT 157.500000 494.410000 158.500000 495.590000 ;
      RECT 116.500000 494.410000 149.500000 495.590000 ;
      RECT 107.500000 494.410000 108.500000 495.590000 ;
      RECT 66.500000 494.410000 99.500000 495.590000 ;
      RECT 57.500000 494.410000 58.500000 495.590000 ;
      RECT 29.500000 494.410000 49.500000 495.590000 ;
      RECT 15.500000 494.410000 16.500000 495.590000 ;
      RECT 1157.500000 493.590000 1186.000000 494.410000 ;
      RECT 707.500000 493.590000 723.500000 494.410000 ;
      RECT 657.500000 493.590000 699.500000 494.410000 ;
      RECT 607.500000 493.590000 649.500000 494.410000 ;
      RECT 557.500000 493.590000 599.500000 494.410000 ;
      RECT 507.500000 493.590000 549.500000 494.410000 ;
      RECT 457.500000 493.590000 499.500000 494.410000 ;
      RECT 407.500000 493.590000 449.500000 494.410000 ;
      RECT 357.500000 493.590000 373.500000 494.410000 ;
      RECT 307.500000 493.590000 349.500000 494.410000 ;
      RECT 257.500000 493.590000 299.500000 494.410000 ;
      RECT 207.500000 493.590000 249.500000 494.410000 ;
      RECT 157.500000 493.590000 199.500000 494.410000 ;
      RECT 107.500000 493.590000 149.500000 494.410000 ;
      RECT 57.500000 493.590000 99.500000 494.410000 ;
      RECT 15.500000 493.590000 49.500000 494.410000 ;
      RECT 1157.500000 492.410000 1158.500000 493.590000 ;
      RECT 1139.000000 492.410000 1149.500000 495.590000 ;
      RECT 736.500000 492.410000 739.000000 495.590000 ;
      RECT 716.500000 492.410000 723.500000 493.590000 ;
      RECT 707.500000 492.410000 708.500000 493.590000 ;
      RECT 666.500000 492.410000 699.500000 493.590000 ;
      RECT 657.500000 492.410000 658.500000 493.590000 ;
      RECT 616.500000 492.410000 649.500000 493.590000 ;
      RECT 607.500000 492.410000 608.500000 493.590000 ;
      RECT 566.500000 492.410000 599.500000 493.590000 ;
      RECT 557.500000 492.410000 558.500000 493.590000 ;
      RECT 516.500000 492.410000 549.500000 493.590000 ;
      RECT 507.500000 492.410000 508.500000 493.590000 ;
      RECT 466.500000 492.410000 499.500000 493.590000 ;
      RECT 457.500000 492.410000 458.500000 493.590000 ;
      RECT 416.500000 492.410000 449.500000 493.590000 ;
      RECT 407.500000 492.410000 408.500000 493.590000 ;
      RECT 386.500000 492.410000 399.500000 495.590000 ;
      RECT 372.500000 492.410000 373.500000 493.590000 ;
      RECT 357.500000 492.410000 358.500000 493.590000 ;
      RECT 316.500000 492.410000 349.500000 493.590000 ;
      RECT 307.500000 492.410000 308.500000 493.590000 ;
      RECT 266.500000 492.410000 299.500000 493.590000 ;
      RECT 257.500000 492.410000 258.500000 493.590000 ;
      RECT 216.500000 492.410000 249.500000 493.590000 ;
      RECT 207.500000 492.410000 208.500000 493.590000 ;
      RECT 166.500000 492.410000 199.500000 493.590000 ;
      RECT 157.500000 492.410000 158.500000 493.590000 ;
      RECT 116.500000 492.410000 149.500000 493.590000 ;
      RECT 107.500000 492.410000 108.500000 493.590000 ;
      RECT 66.500000 492.410000 99.500000 493.590000 ;
      RECT 57.500000 492.410000 58.500000 493.590000 ;
      RECT 29.500000 492.410000 49.500000 493.590000 ;
      RECT 15.500000 492.410000 16.500000 493.590000 ;
      RECT 0.000000 492.410000 2.500000 495.590000 ;
      RECT 1139.000000 491.590000 1158.500000 492.410000 ;
      RECT 716.500000 491.590000 739.000000 492.410000 ;
      RECT 666.500000 491.590000 708.500000 492.410000 ;
      RECT 616.500000 491.590000 658.500000 492.410000 ;
      RECT 566.500000 491.590000 608.500000 492.410000 ;
      RECT 516.500000 491.590000 558.500000 492.410000 ;
      RECT 466.500000 491.590000 508.500000 492.410000 ;
      RECT 416.500000 491.590000 458.500000 492.410000 ;
      RECT 372.500000 491.590000 408.500000 492.410000 ;
      RECT 316.500000 491.590000 358.500000 492.410000 ;
      RECT 266.500000 491.590000 308.500000 492.410000 ;
      RECT 216.500000 491.590000 258.500000 492.410000 ;
      RECT 166.500000 491.590000 208.500000 492.410000 ;
      RECT 116.500000 491.590000 158.500000 492.410000 ;
      RECT 66.500000 491.590000 108.500000 492.410000 ;
      RECT 29.500000 491.590000 58.500000 492.410000 ;
      RECT 0.000000 491.590000 16.500000 492.410000 ;
      RECT 1166.500000 490.410000 1186.000000 493.590000 ;
      RECT 1157.500000 490.410000 1158.500000 491.590000 ;
      RECT 716.500000 490.410000 723.500000 491.590000 ;
      RECT 707.500000 490.410000 708.500000 491.590000 ;
      RECT 666.500000 490.410000 699.500000 491.590000 ;
      RECT 657.500000 490.410000 658.500000 491.590000 ;
      RECT 616.500000 490.410000 649.500000 491.590000 ;
      RECT 607.500000 490.410000 608.500000 491.590000 ;
      RECT 566.500000 490.410000 599.500000 491.590000 ;
      RECT 557.500000 490.410000 558.500000 491.590000 ;
      RECT 516.500000 490.410000 549.500000 491.590000 ;
      RECT 507.500000 490.410000 508.500000 491.590000 ;
      RECT 466.500000 490.410000 499.500000 491.590000 ;
      RECT 457.500000 490.410000 458.500000 491.590000 ;
      RECT 416.500000 490.410000 449.500000 491.590000 ;
      RECT 407.500000 490.410000 408.500000 491.590000 ;
      RECT 372.500000 490.410000 399.500000 491.590000 ;
      RECT 357.500000 490.410000 358.500000 491.590000 ;
      RECT 316.500000 490.410000 349.500000 491.590000 ;
      RECT 307.500000 490.410000 308.500000 491.590000 ;
      RECT 266.500000 490.410000 299.500000 491.590000 ;
      RECT 257.500000 490.410000 258.500000 491.590000 ;
      RECT 216.500000 490.410000 249.500000 491.590000 ;
      RECT 207.500000 490.410000 208.500000 491.590000 ;
      RECT 166.500000 490.410000 199.500000 491.590000 ;
      RECT 157.500000 490.410000 158.500000 491.590000 ;
      RECT 116.500000 490.410000 149.500000 491.590000 ;
      RECT 107.500000 490.410000 108.500000 491.590000 ;
      RECT 66.500000 490.410000 99.500000 491.590000 ;
      RECT 57.500000 490.410000 58.500000 491.590000 ;
      RECT 29.500000 490.410000 49.500000 491.590000 ;
      RECT 15.500000 490.410000 16.500000 491.590000 ;
      RECT 1157.500000 489.590000 1186.000000 490.410000 ;
      RECT 707.500000 489.590000 723.500000 490.410000 ;
      RECT 657.500000 489.590000 699.500000 490.410000 ;
      RECT 607.500000 489.590000 649.500000 490.410000 ;
      RECT 557.500000 489.590000 599.500000 490.410000 ;
      RECT 507.500000 489.590000 549.500000 490.410000 ;
      RECT 457.500000 489.590000 499.500000 490.410000 ;
      RECT 407.500000 489.590000 449.500000 490.410000 ;
      RECT 357.500000 489.590000 399.500000 490.410000 ;
      RECT 307.500000 489.590000 349.500000 490.410000 ;
      RECT 257.500000 489.590000 299.500000 490.410000 ;
      RECT 207.500000 489.590000 249.500000 490.410000 ;
      RECT 157.500000 489.590000 199.500000 490.410000 ;
      RECT 107.500000 489.590000 149.500000 490.410000 ;
      RECT 57.500000 489.590000 99.500000 490.410000 ;
      RECT 15.500000 489.590000 49.500000 490.410000 ;
      RECT 1157.500000 488.410000 1158.500000 489.590000 ;
      RECT 1139.000000 488.410000 1149.500000 491.590000 ;
      RECT 736.500000 488.410000 739.000000 491.590000 ;
      RECT 722.500000 488.410000 723.500000 489.590000 ;
      RECT 707.500000 488.410000 708.500000 489.590000 ;
      RECT 666.500000 488.410000 699.500000 489.590000 ;
      RECT 657.500000 488.410000 658.500000 489.590000 ;
      RECT 616.500000 488.410000 649.500000 489.590000 ;
      RECT 607.500000 488.410000 608.500000 489.590000 ;
      RECT 566.500000 488.410000 599.500000 489.590000 ;
      RECT 557.500000 488.410000 558.500000 489.590000 ;
      RECT 516.500000 488.410000 549.500000 489.590000 ;
      RECT 507.500000 488.410000 508.500000 489.590000 ;
      RECT 466.500000 488.410000 499.500000 489.590000 ;
      RECT 457.500000 488.410000 458.500000 489.590000 ;
      RECT 416.500000 488.410000 449.500000 489.590000 ;
      RECT 407.500000 488.410000 408.500000 489.590000 ;
      RECT 372.500000 488.410000 399.500000 489.590000 ;
      RECT 357.500000 488.410000 359.500000 489.590000 ;
      RECT 316.500000 488.410000 349.500000 489.590000 ;
      RECT 307.500000 488.410000 308.500000 489.590000 ;
      RECT 266.500000 488.410000 299.500000 489.590000 ;
      RECT 257.500000 488.410000 258.500000 489.590000 ;
      RECT 216.500000 488.410000 249.500000 489.590000 ;
      RECT 207.500000 488.410000 208.500000 489.590000 ;
      RECT 166.500000 488.410000 199.500000 489.590000 ;
      RECT 157.500000 488.410000 158.500000 489.590000 ;
      RECT 116.500000 488.410000 149.500000 489.590000 ;
      RECT 107.500000 488.410000 108.500000 489.590000 ;
      RECT 66.500000 488.410000 99.500000 489.590000 ;
      RECT 57.500000 488.410000 58.500000 489.590000 ;
      RECT 29.500000 488.410000 49.500000 489.590000 ;
      RECT 15.500000 488.410000 16.500000 489.590000 ;
      RECT 0.000000 488.410000 2.500000 491.590000 ;
      RECT 1139.000000 487.590000 1158.500000 488.410000 ;
      RECT 722.500000 487.590000 739.000000 488.410000 ;
      RECT 666.500000 487.590000 708.500000 488.410000 ;
      RECT 616.500000 487.590000 658.500000 488.410000 ;
      RECT 566.500000 487.590000 608.500000 488.410000 ;
      RECT 516.500000 487.590000 558.500000 488.410000 ;
      RECT 466.500000 487.590000 508.500000 488.410000 ;
      RECT 416.500000 487.590000 458.500000 488.410000 ;
      RECT 372.500000 487.590000 408.500000 488.410000 ;
      RECT 316.500000 487.590000 359.500000 488.410000 ;
      RECT 266.500000 487.590000 308.500000 488.410000 ;
      RECT 216.500000 487.590000 258.500000 488.410000 ;
      RECT 166.500000 487.590000 208.500000 488.410000 ;
      RECT 116.500000 487.590000 158.500000 488.410000 ;
      RECT 66.500000 487.590000 108.500000 488.410000 ;
      RECT 29.500000 487.590000 58.500000 488.410000 ;
      RECT 0.000000 487.590000 16.500000 488.410000 ;
      RECT 0.000000 487.170000 2.500000 487.590000 ;
      RECT 1166.500000 487.165000 1186.000000 489.590000 ;
      RECT 1166.500000 486.410000 1183.980000 487.165000 ;
      RECT 1157.500000 486.410000 1158.500000 487.590000 ;
      RECT 722.500000 486.410000 723.500000 487.590000 ;
      RECT 707.500000 486.410000 708.500000 487.590000 ;
      RECT 666.500000 486.410000 699.500000 487.590000 ;
      RECT 657.500000 486.410000 658.500000 487.590000 ;
      RECT 616.500000 486.410000 649.500000 487.590000 ;
      RECT 607.500000 486.410000 608.500000 487.590000 ;
      RECT 566.500000 486.410000 599.500000 487.590000 ;
      RECT 557.500000 486.410000 558.500000 487.590000 ;
      RECT 516.500000 486.410000 549.500000 487.590000 ;
      RECT 507.500000 486.410000 508.500000 487.590000 ;
      RECT 466.500000 486.410000 499.500000 487.590000 ;
      RECT 457.500000 486.410000 458.500000 487.590000 ;
      RECT 416.500000 486.410000 449.500000 487.590000 ;
      RECT 407.500000 486.410000 408.500000 487.590000 ;
      RECT 372.500000 486.410000 399.500000 487.590000 ;
      RECT 357.500000 486.410000 359.500000 487.590000 ;
      RECT 316.500000 486.410000 349.500000 487.590000 ;
      RECT 307.500000 486.410000 308.500000 487.590000 ;
      RECT 266.500000 486.410000 299.500000 487.590000 ;
      RECT 257.500000 486.410000 258.500000 487.590000 ;
      RECT 216.500000 486.410000 249.500000 487.590000 ;
      RECT 207.500000 486.410000 208.500000 487.590000 ;
      RECT 166.500000 486.410000 199.500000 487.590000 ;
      RECT 157.500000 486.410000 158.500000 487.590000 ;
      RECT 116.500000 486.410000 149.500000 487.590000 ;
      RECT 107.500000 486.410000 108.500000 487.590000 ;
      RECT 66.500000 486.410000 99.500000 487.590000 ;
      RECT 57.500000 486.410000 58.500000 487.590000 ;
      RECT 29.500000 486.410000 49.500000 487.590000 ;
      RECT 15.500000 486.410000 16.500000 487.590000 ;
      RECT 1157.500000 485.590000 1183.980000 486.410000 ;
      RECT 707.500000 485.590000 723.500000 486.410000 ;
      RECT 657.500000 485.590000 699.500000 486.410000 ;
      RECT 607.500000 485.590000 649.500000 486.410000 ;
      RECT 557.500000 485.590000 599.500000 486.410000 ;
      RECT 507.500000 485.590000 549.500000 486.410000 ;
      RECT 457.500000 485.590000 499.500000 486.410000 ;
      RECT 407.500000 485.590000 449.500000 486.410000 ;
      RECT 357.500000 485.590000 399.500000 486.410000 ;
      RECT 307.500000 485.590000 349.500000 486.410000 ;
      RECT 257.500000 485.590000 299.500000 486.410000 ;
      RECT 207.500000 485.590000 249.500000 486.410000 ;
      RECT 157.500000 485.590000 199.500000 486.410000 ;
      RECT 107.500000 485.590000 149.500000 486.410000 ;
      RECT 57.500000 485.590000 99.500000 486.410000 ;
      RECT 15.500000 485.590000 49.500000 486.410000 ;
      RECT 1157.500000 484.410000 1158.500000 485.590000 ;
      RECT 1139.000000 484.410000 1149.500000 487.590000 ;
      RECT 736.500000 484.410000 739.000000 487.590000 ;
      RECT 722.500000 484.410000 723.500000 485.590000 ;
      RECT 707.500000 484.410000 708.500000 485.590000 ;
      RECT 666.500000 484.410000 699.500000 485.590000 ;
      RECT 657.500000 484.410000 658.500000 485.590000 ;
      RECT 616.500000 484.410000 649.500000 485.590000 ;
      RECT 607.500000 484.410000 608.500000 485.590000 ;
      RECT 566.500000 484.410000 599.500000 485.590000 ;
      RECT 557.500000 484.410000 558.500000 485.590000 ;
      RECT 516.500000 484.410000 549.500000 485.590000 ;
      RECT 507.500000 484.410000 508.500000 485.590000 ;
      RECT 466.500000 484.410000 499.500000 485.590000 ;
      RECT 457.500000 484.410000 458.500000 485.590000 ;
      RECT 416.500000 484.410000 449.500000 485.590000 ;
      RECT 407.500000 484.410000 408.500000 485.590000 ;
      RECT 372.500000 484.410000 399.500000 485.590000 ;
      RECT 357.500000 484.410000 359.500000 485.590000 ;
      RECT 316.500000 484.410000 349.500000 485.590000 ;
      RECT 307.500000 484.410000 308.500000 485.590000 ;
      RECT 266.500000 484.410000 299.500000 485.590000 ;
      RECT 257.500000 484.410000 258.500000 485.590000 ;
      RECT 216.500000 484.410000 249.500000 485.590000 ;
      RECT 207.500000 484.410000 208.500000 485.590000 ;
      RECT 166.500000 484.410000 199.500000 485.590000 ;
      RECT 157.500000 484.410000 158.500000 485.590000 ;
      RECT 116.500000 484.410000 149.500000 485.590000 ;
      RECT 107.500000 484.410000 108.500000 485.590000 ;
      RECT 66.500000 484.410000 99.500000 485.590000 ;
      RECT 57.500000 484.410000 58.500000 485.590000 ;
      RECT 29.500000 484.410000 49.500000 485.590000 ;
      RECT 15.500000 484.410000 16.500000 485.590000 ;
      RECT 2.020000 484.410000 2.500000 487.170000 ;
      RECT 2.020000 484.070000 16.500000 484.410000 ;
      RECT 1166.500000 484.065000 1183.980000 485.590000 ;
      RECT 1139.000000 483.590000 1158.500000 484.410000 ;
      RECT 722.500000 483.590000 739.000000 484.410000 ;
      RECT 666.500000 483.590000 708.500000 484.410000 ;
      RECT 616.500000 483.590000 658.500000 484.410000 ;
      RECT 566.500000 483.590000 608.500000 484.410000 ;
      RECT 516.500000 483.590000 558.500000 484.410000 ;
      RECT 466.500000 483.590000 508.500000 484.410000 ;
      RECT 416.500000 483.590000 458.500000 484.410000 ;
      RECT 372.500000 483.590000 408.500000 484.410000 ;
      RECT 316.500000 483.590000 359.500000 484.410000 ;
      RECT 266.500000 483.590000 308.500000 484.410000 ;
      RECT 216.500000 483.590000 258.500000 484.410000 ;
      RECT 166.500000 483.590000 208.500000 484.410000 ;
      RECT 116.500000 483.590000 158.500000 484.410000 ;
      RECT 66.500000 483.590000 108.500000 484.410000 ;
      RECT 29.500000 483.590000 58.500000 484.410000 ;
      RECT 0.000000 483.590000 16.500000 484.070000 ;
      RECT 1166.500000 482.410000 1186.000000 484.065000 ;
      RECT 1157.500000 482.410000 1158.500000 483.590000 ;
      RECT 722.500000 482.410000 723.500000 483.590000 ;
      RECT 707.500000 482.410000 708.500000 483.590000 ;
      RECT 666.500000 482.410000 699.500000 483.590000 ;
      RECT 657.500000 482.410000 658.500000 483.590000 ;
      RECT 616.500000 482.410000 649.500000 483.590000 ;
      RECT 607.500000 482.410000 608.500000 483.590000 ;
      RECT 566.500000 482.410000 599.500000 483.590000 ;
      RECT 557.500000 482.410000 558.500000 483.590000 ;
      RECT 516.500000 482.410000 549.500000 483.590000 ;
      RECT 507.500000 482.410000 508.500000 483.590000 ;
      RECT 466.500000 482.410000 499.500000 483.590000 ;
      RECT 457.500000 482.410000 458.500000 483.590000 ;
      RECT 416.500000 482.410000 449.500000 483.590000 ;
      RECT 407.500000 482.410000 408.500000 483.590000 ;
      RECT 372.500000 482.410000 399.500000 483.590000 ;
      RECT 357.500000 482.410000 359.500000 483.590000 ;
      RECT 316.500000 482.410000 349.500000 483.590000 ;
      RECT 307.500000 482.410000 308.500000 483.590000 ;
      RECT 266.500000 482.410000 299.500000 483.590000 ;
      RECT 257.500000 482.410000 258.500000 483.590000 ;
      RECT 216.500000 482.410000 249.500000 483.590000 ;
      RECT 207.500000 482.410000 208.500000 483.590000 ;
      RECT 166.500000 482.410000 199.500000 483.590000 ;
      RECT 157.500000 482.410000 158.500000 483.590000 ;
      RECT 116.500000 482.410000 149.500000 483.590000 ;
      RECT 107.500000 482.410000 108.500000 483.590000 ;
      RECT 66.500000 482.410000 99.500000 483.590000 ;
      RECT 57.500000 482.410000 58.500000 483.590000 ;
      RECT 29.500000 482.410000 49.500000 483.590000 ;
      RECT 15.500000 482.410000 16.500000 483.590000 ;
      RECT 1157.500000 481.590000 1186.000000 482.410000 ;
      RECT 707.500000 481.590000 723.500000 482.410000 ;
      RECT 657.500000 481.590000 699.500000 482.410000 ;
      RECT 607.500000 481.590000 649.500000 482.410000 ;
      RECT 557.500000 481.590000 599.500000 482.410000 ;
      RECT 507.500000 481.590000 549.500000 482.410000 ;
      RECT 457.500000 481.590000 499.500000 482.410000 ;
      RECT 407.500000 481.590000 449.500000 482.410000 ;
      RECT 357.500000 481.590000 399.500000 482.410000 ;
      RECT 307.500000 481.590000 349.500000 482.410000 ;
      RECT 257.500000 481.590000 299.500000 482.410000 ;
      RECT 207.500000 481.590000 249.500000 482.410000 ;
      RECT 157.500000 481.590000 199.500000 482.410000 ;
      RECT 107.500000 481.590000 149.500000 482.410000 ;
      RECT 57.500000 481.590000 99.500000 482.410000 ;
      RECT 15.500000 481.590000 49.500000 482.410000 ;
      RECT 1166.500000 481.485000 1186.000000 481.590000 ;
      RECT 1157.500000 480.410000 1158.500000 481.590000 ;
      RECT 1139.000000 480.410000 1149.500000 483.590000 ;
      RECT 736.500000 480.410000 739.000000 483.590000 ;
      RECT 722.500000 480.410000 723.500000 481.590000 ;
      RECT 707.500000 480.410000 708.500000 481.590000 ;
      RECT 666.500000 480.410000 699.500000 481.590000 ;
      RECT 657.500000 480.410000 658.500000 481.590000 ;
      RECT 616.500000 480.410000 649.500000 481.590000 ;
      RECT 607.500000 480.410000 608.500000 481.590000 ;
      RECT 566.500000 480.410000 599.500000 481.590000 ;
      RECT 557.500000 480.410000 558.500000 481.590000 ;
      RECT 516.500000 480.410000 549.500000 481.590000 ;
      RECT 507.500000 480.410000 508.500000 481.590000 ;
      RECT 466.500000 480.410000 499.500000 481.590000 ;
      RECT 457.500000 480.410000 458.500000 481.590000 ;
      RECT 416.500000 480.410000 449.500000 481.590000 ;
      RECT 407.500000 480.410000 408.500000 481.590000 ;
      RECT 372.500000 480.410000 399.500000 481.590000 ;
      RECT 357.500000 480.410000 359.500000 481.590000 ;
      RECT 316.500000 480.410000 349.500000 481.590000 ;
      RECT 307.500000 480.410000 308.500000 481.590000 ;
      RECT 266.500000 480.410000 299.500000 481.590000 ;
      RECT 257.500000 480.410000 258.500000 481.590000 ;
      RECT 216.500000 480.410000 249.500000 481.590000 ;
      RECT 207.500000 480.410000 208.500000 481.590000 ;
      RECT 166.500000 480.410000 199.500000 481.590000 ;
      RECT 157.500000 480.410000 158.500000 481.590000 ;
      RECT 116.500000 480.410000 149.500000 481.590000 ;
      RECT 107.500000 480.410000 108.500000 481.590000 ;
      RECT 66.500000 480.410000 99.500000 481.590000 ;
      RECT 57.500000 480.410000 58.500000 481.590000 ;
      RECT 29.500000 480.410000 49.500000 481.590000 ;
      RECT 15.500000 480.410000 16.500000 481.590000 ;
      RECT 0.000000 480.410000 2.500000 483.590000 ;
      RECT 1139.000000 479.590000 1158.500000 480.410000 ;
      RECT 722.500000 479.590000 739.000000 480.410000 ;
      RECT 666.500000 479.590000 708.500000 480.410000 ;
      RECT 616.500000 479.590000 658.500000 480.410000 ;
      RECT 566.500000 479.590000 608.500000 480.410000 ;
      RECT 516.500000 479.590000 558.500000 480.410000 ;
      RECT 466.500000 479.590000 508.500000 480.410000 ;
      RECT 416.500000 479.590000 458.500000 480.410000 ;
      RECT 372.500000 479.590000 408.500000 480.410000 ;
      RECT 316.500000 479.590000 359.500000 480.410000 ;
      RECT 266.500000 479.590000 308.500000 480.410000 ;
      RECT 216.500000 479.590000 258.500000 480.410000 ;
      RECT 166.500000 479.590000 208.500000 480.410000 ;
      RECT 116.500000 479.590000 158.500000 480.410000 ;
      RECT 66.500000 479.590000 108.500000 480.410000 ;
      RECT 29.500000 479.590000 58.500000 480.410000 ;
      RECT 0.000000 479.590000 16.500000 480.410000 ;
      RECT 1166.500000 478.410000 1183.980000 481.485000 ;
      RECT 1157.500000 478.410000 1158.500000 479.590000 ;
      RECT 722.500000 478.410000 723.500000 479.590000 ;
      RECT 707.500000 478.410000 708.500000 479.590000 ;
      RECT 666.500000 478.410000 699.500000 479.590000 ;
      RECT 657.500000 478.410000 658.500000 479.590000 ;
      RECT 616.500000 478.410000 649.500000 479.590000 ;
      RECT 607.500000 478.410000 608.500000 479.590000 ;
      RECT 566.500000 478.410000 599.500000 479.590000 ;
      RECT 557.500000 478.410000 558.500000 479.590000 ;
      RECT 516.500000 478.410000 549.500000 479.590000 ;
      RECT 507.500000 478.410000 508.500000 479.590000 ;
      RECT 466.500000 478.410000 499.500000 479.590000 ;
      RECT 457.500000 478.410000 458.500000 479.590000 ;
      RECT 416.500000 478.410000 449.500000 479.590000 ;
      RECT 407.500000 478.410000 408.500000 479.590000 ;
      RECT 372.500000 478.410000 399.500000 479.590000 ;
      RECT 357.500000 478.410000 359.500000 479.590000 ;
      RECT 316.500000 478.410000 349.500000 479.590000 ;
      RECT 307.500000 478.410000 308.500000 479.590000 ;
      RECT 266.500000 478.410000 299.500000 479.590000 ;
      RECT 257.500000 478.410000 258.500000 479.590000 ;
      RECT 216.500000 478.410000 249.500000 479.590000 ;
      RECT 207.500000 478.410000 208.500000 479.590000 ;
      RECT 166.500000 478.410000 199.500000 479.590000 ;
      RECT 157.500000 478.410000 158.500000 479.590000 ;
      RECT 116.500000 478.410000 149.500000 479.590000 ;
      RECT 107.500000 478.410000 108.500000 479.590000 ;
      RECT 66.500000 478.410000 99.500000 479.590000 ;
      RECT 57.500000 478.410000 58.500000 479.590000 ;
      RECT 29.500000 478.410000 49.500000 479.590000 ;
      RECT 15.500000 478.410000 16.500000 479.590000 ;
      RECT 1157.500000 478.385000 1183.980000 478.410000 ;
      RECT 1157.500000 477.590000 1186.000000 478.385000 ;
      RECT 707.500000 477.590000 723.500000 478.410000 ;
      RECT 657.500000 477.590000 699.500000 478.410000 ;
      RECT 607.500000 477.590000 649.500000 478.410000 ;
      RECT 557.500000 477.590000 599.500000 478.410000 ;
      RECT 507.500000 477.590000 549.500000 478.410000 ;
      RECT 457.500000 477.590000 499.500000 478.410000 ;
      RECT 407.500000 477.590000 449.500000 478.410000 ;
      RECT 357.500000 477.590000 399.500000 478.410000 ;
      RECT 307.500000 477.590000 349.500000 478.410000 ;
      RECT 257.500000 477.590000 299.500000 478.410000 ;
      RECT 207.500000 477.590000 249.500000 478.410000 ;
      RECT 157.500000 477.590000 199.500000 478.410000 ;
      RECT 107.500000 477.590000 149.500000 478.410000 ;
      RECT 57.500000 477.590000 99.500000 478.410000 ;
      RECT 15.500000 477.590000 49.500000 478.410000 ;
      RECT 1166.500000 477.525000 1186.000000 477.590000 ;
      RECT 0.000000 476.575000 2.500000 479.590000 ;
      RECT 1157.500000 476.410000 1158.500000 477.590000 ;
      RECT 1139.000000 476.410000 1149.500000 479.590000 ;
      RECT 736.500000 476.410000 739.000000 479.590000 ;
      RECT 722.500000 476.410000 723.500000 477.590000 ;
      RECT 707.500000 476.410000 708.500000 477.590000 ;
      RECT 666.500000 476.410000 699.500000 477.590000 ;
      RECT 657.500000 476.410000 658.500000 477.590000 ;
      RECT 616.500000 476.410000 649.500000 477.590000 ;
      RECT 607.500000 476.410000 608.500000 477.590000 ;
      RECT 566.500000 476.410000 599.500000 477.590000 ;
      RECT 557.500000 476.410000 558.500000 477.590000 ;
      RECT 516.500000 476.410000 549.500000 477.590000 ;
      RECT 507.500000 476.410000 508.500000 477.590000 ;
      RECT 466.500000 476.410000 499.500000 477.590000 ;
      RECT 457.500000 476.410000 458.500000 477.590000 ;
      RECT 416.500000 476.410000 449.500000 477.590000 ;
      RECT 407.500000 476.410000 408.500000 477.590000 ;
      RECT 370.000000 476.410000 399.500000 477.590000 ;
      RECT 357.500000 476.410000 362.000000 477.590000 ;
      RECT 316.500000 476.410000 349.500000 477.590000 ;
      RECT 307.500000 476.410000 308.500000 477.590000 ;
      RECT 266.500000 476.410000 299.500000 477.590000 ;
      RECT 257.500000 476.410000 258.500000 477.590000 ;
      RECT 216.500000 476.410000 249.500000 477.590000 ;
      RECT 207.500000 476.410000 208.500000 477.590000 ;
      RECT 166.500000 476.410000 199.500000 477.590000 ;
      RECT 157.500000 476.410000 158.500000 477.590000 ;
      RECT 116.500000 476.410000 149.500000 477.590000 ;
      RECT 107.500000 476.410000 108.500000 477.590000 ;
      RECT 66.500000 476.410000 99.500000 477.590000 ;
      RECT 57.500000 476.410000 58.500000 477.590000 ;
      RECT 29.500000 476.410000 49.500000 477.590000 ;
      RECT 15.500000 476.410000 16.500000 477.590000 ;
      RECT 2.020000 476.410000 2.500000 476.575000 ;
      RECT 1139.000000 475.590000 1158.500000 476.410000 ;
      RECT 722.500000 475.590000 739.000000 476.410000 ;
      RECT 666.500000 475.590000 708.500000 476.410000 ;
      RECT 616.500000 475.590000 658.500000 476.410000 ;
      RECT 566.500000 475.590000 608.500000 476.410000 ;
      RECT 516.500000 475.590000 558.500000 476.410000 ;
      RECT 466.500000 475.590000 508.500000 476.410000 ;
      RECT 416.500000 475.590000 458.500000 476.410000 ;
      RECT 370.000000 475.590000 408.500000 476.410000 ;
      RECT 316.500000 475.590000 362.000000 476.410000 ;
      RECT 266.500000 475.590000 308.500000 476.410000 ;
      RECT 216.500000 475.590000 258.500000 476.410000 ;
      RECT 166.500000 475.590000 208.500000 476.410000 ;
      RECT 116.500000 475.590000 158.500000 476.410000 ;
      RECT 66.500000 475.590000 108.500000 476.410000 ;
      RECT 29.500000 475.590000 58.500000 476.410000 ;
      RECT 2.020000 475.590000 16.500000 476.410000 ;
      RECT 1166.500000 474.425000 1183.980000 477.525000 ;
      RECT 1166.500000 474.410000 1186.000000 474.425000 ;
      RECT 1157.500000 474.410000 1158.500000 475.590000 ;
      RECT 722.500000 474.410000 723.500000 475.590000 ;
      RECT 707.500000 474.410000 708.500000 475.590000 ;
      RECT 666.500000 474.410000 699.500000 475.590000 ;
      RECT 657.500000 474.410000 658.500000 475.590000 ;
      RECT 616.500000 474.410000 649.500000 475.590000 ;
      RECT 607.500000 474.410000 608.500000 475.590000 ;
      RECT 566.500000 474.410000 599.500000 475.590000 ;
      RECT 557.500000 474.410000 558.500000 475.590000 ;
      RECT 516.500000 474.410000 549.500000 475.590000 ;
      RECT 507.500000 474.410000 508.500000 475.590000 ;
      RECT 466.500000 474.410000 499.500000 475.590000 ;
      RECT 457.500000 474.410000 458.500000 475.590000 ;
      RECT 416.500000 474.410000 449.500000 475.590000 ;
      RECT 407.500000 474.410000 408.500000 475.590000 ;
      RECT 370.000000 474.410000 399.500000 475.590000 ;
      RECT 357.500000 474.410000 362.000000 475.590000 ;
      RECT 316.500000 474.410000 349.500000 475.590000 ;
      RECT 307.500000 474.410000 308.500000 475.590000 ;
      RECT 266.500000 474.410000 299.500000 475.590000 ;
      RECT 257.500000 474.410000 258.500000 475.590000 ;
      RECT 216.500000 474.410000 249.500000 475.590000 ;
      RECT 207.500000 474.410000 208.500000 475.590000 ;
      RECT 166.500000 474.410000 199.500000 475.590000 ;
      RECT 157.500000 474.410000 158.500000 475.590000 ;
      RECT 116.500000 474.410000 149.500000 475.590000 ;
      RECT 107.500000 474.410000 108.500000 475.590000 ;
      RECT 66.500000 474.410000 99.500000 475.590000 ;
      RECT 57.500000 474.410000 58.500000 475.590000 ;
      RECT 29.500000 474.410000 49.500000 475.590000 ;
      RECT 15.500000 474.410000 16.500000 475.590000 ;
      RECT 1157.500000 473.590000 1186.000000 474.410000 ;
      RECT 707.500000 473.590000 723.500000 474.410000 ;
      RECT 657.500000 473.590000 699.500000 474.410000 ;
      RECT 607.500000 473.590000 649.500000 474.410000 ;
      RECT 557.500000 473.590000 599.500000 474.410000 ;
      RECT 507.500000 473.590000 549.500000 474.410000 ;
      RECT 457.500000 473.590000 499.500000 474.410000 ;
      RECT 407.500000 473.590000 449.500000 474.410000 ;
      RECT 357.500000 473.590000 399.500000 474.410000 ;
      RECT 307.500000 473.590000 349.500000 474.410000 ;
      RECT 257.500000 473.590000 299.500000 474.410000 ;
      RECT 207.500000 473.590000 249.500000 474.410000 ;
      RECT 157.500000 473.590000 199.500000 474.410000 ;
      RECT 107.500000 473.590000 149.500000 474.410000 ;
      RECT 57.500000 473.590000 99.500000 474.410000 ;
      RECT 15.500000 473.590000 49.500000 474.410000 ;
      RECT 2.020000 473.475000 2.500000 475.590000 ;
      RECT 0.000000 472.615000 2.500000 473.475000 ;
      RECT 1157.500000 472.410000 1158.500000 473.590000 ;
      RECT 1139.000000 472.410000 1149.500000 475.590000 ;
      RECT 736.500000 472.410000 739.000000 475.590000 ;
      RECT 722.500000 472.410000 723.500000 473.590000 ;
      RECT 707.500000 472.410000 708.500000 473.590000 ;
      RECT 666.500000 472.410000 699.500000 473.590000 ;
      RECT 657.500000 472.410000 658.500000 473.590000 ;
      RECT 616.500000 472.410000 649.500000 473.590000 ;
      RECT 607.500000 472.410000 608.500000 473.590000 ;
      RECT 566.500000 472.410000 599.500000 473.590000 ;
      RECT 557.500000 472.410000 558.500000 473.590000 ;
      RECT 516.500000 472.410000 549.500000 473.590000 ;
      RECT 507.500000 472.410000 508.500000 473.590000 ;
      RECT 466.500000 472.410000 499.500000 473.590000 ;
      RECT 457.500000 472.410000 458.500000 473.590000 ;
      RECT 416.500000 472.410000 449.500000 473.590000 ;
      RECT 407.500000 472.410000 408.500000 473.590000 ;
      RECT 370.000000 472.410000 399.500000 473.590000 ;
      RECT 357.500000 472.410000 358.500000 473.590000 ;
      RECT 316.500000 472.410000 349.500000 473.590000 ;
      RECT 307.500000 472.410000 308.500000 473.590000 ;
      RECT 266.500000 472.410000 299.500000 473.590000 ;
      RECT 257.500000 472.410000 258.500000 473.590000 ;
      RECT 216.500000 472.410000 249.500000 473.590000 ;
      RECT 207.500000 472.410000 208.500000 473.590000 ;
      RECT 166.500000 472.410000 199.500000 473.590000 ;
      RECT 157.500000 472.410000 158.500000 473.590000 ;
      RECT 116.500000 472.410000 149.500000 473.590000 ;
      RECT 107.500000 472.410000 108.500000 473.590000 ;
      RECT 66.500000 472.410000 99.500000 473.590000 ;
      RECT 57.500000 472.410000 58.500000 473.590000 ;
      RECT 29.500000 472.410000 49.500000 473.590000 ;
      RECT 15.500000 472.410000 16.500000 473.590000 ;
      RECT 2.020000 472.410000 2.500000 472.615000 ;
      RECT 1139.000000 471.590000 1158.500000 472.410000 ;
      RECT 722.500000 471.590000 739.000000 472.410000 ;
      RECT 666.500000 471.590000 708.500000 472.410000 ;
      RECT 616.500000 471.590000 658.500000 472.410000 ;
      RECT 566.500000 471.590000 608.500000 472.410000 ;
      RECT 516.500000 471.590000 558.500000 472.410000 ;
      RECT 466.500000 471.590000 508.500000 472.410000 ;
      RECT 416.500000 471.590000 458.500000 472.410000 ;
      RECT 370.000000 471.590000 408.500000 472.410000 ;
      RECT 316.500000 471.590000 358.500000 472.410000 ;
      RECT 266.500000 471.590000 308.500000 472.410000 ;
      RECT 216.500000 471.590000 258.500000 472.410000 ;
      RECT 166.500000 471.590000 208.500000 472.410000 ;
      RECT 116.500000 471.590000 158.500000 472.410000 ;
      RECT 66.500000 471.590000 108.500000 472.410000 ;
      RECT 29.500000 471.590000 58.500000 472.410000 ;
      RECT 2.020000 471.590000 16.500000 472.410000 ;
      RECT 1166.500000 470.410000 1186.000000 473.590000 ;
      RECT 1157.500000 470.410000 1158.500000 471.590000 ;
      RECT 722.500000 470.410000 723.500000 471.590000 ;
      RECT 707.500000 470.410000 708.500000 471.590000 ;
      RECT 666.500000 470.410000 699.500000 471.590000 ;
      RECT 657.500000 470.410000 658.500000 471.590000 ;
      RECT 616.500000 470.410000 649.500000 471.590000 ;
      RECT 607.500000 470.410000 608.500000 471.590000 ;
      RECT 566.500000 470.410000 599.500000 471.590000 ;
      RECT 557.500000 470.410000 558.500000 471.590000 ;
      RECT 516.500000 470.410000 549.500000 471.590000 ;
      RECT 507.500000 470.410000 508.500000 471.590000 ;
      RECT 466.500000 470.410000 499.500000 471.590000 ;
      RECT 457.500000 470.410000 458.500000 471.590000 ;
      RECT 416.500000 470.410000 449.500000 471.590000 ;
      RECT 407.500000 470.410000 408.500000 471.590000 ;
      RECT 370.000000 470.410000 399.500000 471.590000 ;
      RECT 357.500000 470.410000 358.500000 471.590000 ;
      RECT 316.500000 470.410000 349.500000 471.590000 ;
      RECT 307.500000 470.410000 308.500000 471.590000 ;
      RECT 266.500000 470.410000 299.500000 471.590000 ;
      RECT 257.500000 470.410000 258.500000 471.590000 ;
      RECT 216.500000 470.410000 249.500000 471.590000 ;
      RECT 207.500000 470.410000 208.500000 471.590000 ;
      RECT 166.500000 470.410000 199.500000 471.590000 ;
      RECT 157.500000 470.410000 158.500000 471.590000 ;
      RECT 116.500000 470.410000 149.500000 471.590000 ;
      RECT 107.500000 470.410000 108.500000 471.590000 ;
      RECT 66.500000 470.410000 99.500000 471.590000 ;
      RECT 57.500000 470.410000 58.500000 471.590000 ;
      RECT 29.500000 470.410000 49.500000 471.590000 ;
      RECT 15.500000 470.410000 16.500000 471.590000 ;
      RECT 1157.500000 469.590000 1186.000000 470.410000 ;
      RECT 707.500000 469.590000 723.500000 470.410000 ;
      RECT 657.500000 469.590000 699.500000 470.410000 ;
      RECT 607.500000 469.590000 649.500000 470.410000 ;
      RECT 557.500000 469.590000 599.500000 470.410000 ;
      RECT 507.500000 469.590000 549.500000 470.410000 ;
      RECT 457.500000 469.590000 499.500000 470.410000 ;
      RECT 407.500000 469.590000 449.500000 470.410000 ;
      RECT 357.500000 469.590000 399.500000 470.410000 ;
      RECT 307.500000 469.590000 349.500000 470.410000 ;
      RECT 257.500000 469.590000 299.500000 470.410000 ;
      RECT 207.500000 469.590000 249.500000 470.410000 ;
      RECT 157.500000 469.590000 199.500000 470.410000 ;
      RECT 107.500000 469.590000 149.500000 470.410000 ;
      RECT 57.500000 469.590000 99.500000 470.410000 ;
      RECT 15.500000 469.590000 49.500000 470.410000 ;
      RECT 2.020000 469.515000 2.500000 471.590000 ;
      RECT 1157.500000 468.410000 1158.500000 469.590000 ;
      RECT 1139.000000 468.410000 1149.500000 471.590000 ;
      RECT 736.500000 468.410000 739.000000 471.590000 ;
      RECT 722.500000 468.410000 723.500000 469.590000 ;
      RECT 707.500000 468.410000 708.500000 469.590000 ;
      RECT 666.500000 468.410000 699.500000 469.590000 ;
      RECT 657.500000 468.410000 658.500000 469.590000 ;
      RECT 616.500000 468.410000 649.500000 469.590000 ;
      RECT 607.500000 468.410000 608.500000 469.590000 ;
      RECT 566.500000 468.410000 599.500000 469.590000 ;
      RECT 557.500000 468.410000 558.500000 469.590000 ;
      RECT 516.500000 468.410000 549.500000 469.590000 ;
      RECT 507.500000 468.410000 508.500000 469.590000 ;
      RECT 466.500000 468.410000 499.500000 469.590000 ;
      RECT 457.500000 468.410000 458.500000 469.590000 ;
      RECT 416.500000 468.410000 449.500000 469.590000 ;
      RECT 407.500000 468.410000 408.500000 469.590000 ;
      RECT 366.500000 468.410000 399.500000 469.590000 ;
      RECT 357.500000 468.410000 358.500000 469.590000 ;
      RECT 316.500000 468.410000 349.500000 469.590000 ;
      RECT 307.500000 468.410000 308.500000 469.590000 ;
      RECT 266.500000 468.410000 299.500000 469.590000 ;
      RECT 257.500000 468.410000 258.500000 469.590000 ;
      RECT 216.500000 468.410000 249.500000 469.590000 ;
      RECT 207.500000 468.410000 208.500000 469.590000 ;
      RECT 166.500000 468.410000 199.500000 469.590000 ;
      RECT 157.500000 468.410000 158.500000 469.590000 ;
      RECT 116.500000 468.410000 149.500000 469.590000 ;
      RECT 107.500000 468.410000 108.500000 469.590000 ;
      RECT 66.500000 468.410000 99.500000 469.590000 ;
      RECT 57.500000 468.410000 58.500000 469.590000 ;
      RECT 29.500000 468.410000 49.500000 469.590000 ;
      RECT 15.500000 468.410000 16.500000 469.590000 ;
      RECT 0.000000 468.410000 2.500000 469.515000 ;
      RECT 1139.000000 467.590000 1158.500000 468.410000 ;
      RECT 722.500000 467.590000 739.000000 468.410000 ;
      RECT 666.500000 467.590000 708.500000 468.410000 ;
      RECT 616.500000 467.590000 658.500000 468.410000 ;
      RECT 566.500000 467.590000 608.500000 468.410000 ;
      RECT 516.500000 467.590000 558.500000 468.410000 ;
      RECT 466.500000 467.590000 508.500000 468.410000 ;
      RECT 416.500000 467.590000 458.500000 468.410000 ;
      RECT 366.500000 467.590000 408.500000 468.410000 ;
      RECT 316.500000 467.590000 358.500000 468.410000 ;
      RECT 266.500000 467.590000 308.500000 468.410000 ;
      RECT 216.500000 467.590000 258.500000 468.410000 ;
      RECT 166.500000 467.590000 208.500000 468.410000 ;
      RECT 116.500000 467.590000 158.500000 468.410000 ;
      RECT 66.500000 467.590000 108.500000 468.410000 ;
      RECT 29.500000 467.590000 58.500000 468.410000 ;
      RECT 0.000000 467.590000 16.500000 468.410000 ;
      RECT 0.000000 466.935000 2.500000 467.590000 ;
      RECT 1166.500000 466.930000 1186.000000 469.590000 ;
      RECT 1166.500000 466.410000 1183.980000 466.930000 ;
      RECT 1157.500000 466.410000 1158.500000 467.590000 ;
      RECT 722.500000 466.410000 723.500000 467.590000 ;
      RECT 707.500000 466.410000 708.500000 467.590000 ;
      RECT 666.500000 466.410000 699.500000 467.590000 ;
      RECT 657.500000 466.410000 658.500000 467.590000 ;
      RECT 616.500000 466.410000 649.500000 467.590000 ;
      RECT 607.500000 466.410000 608.500000 467.590000 ;
      RECT 566.500000 466.410000 599.500000 467.590000 ;
      RECT 557.500000 466.410000 558.500000 467.590000 ;
      RECT 516.500000 466.410000 549.500000 467.590000 ;
      RECT 507.500000 466.410000 508.500000 467.590000 ;
      RECT 466.500000 466.410000 499.500000 467.590000 ;
      RECT 457.500000 466.410000 458.500000 467.590000 ;
      RECT 416.500000 466.410000 449.500000 467.590000 ;
      RECT 407.500000 466.410000 408.500000 467.590000 ;
      RECT 366.500000 466.410000 399.500000 467.590000 ;
      RECT 357.500000 466.410000 358.500000 467.590000 ;
      RECT 316.500000 466.410000 349.500000 467.590000 ;
      RECT 307.500000 466.410000 308.500000 467.590000 ;
      RECT 266.500000 466.410000 299.500000 467.590000 ;
      RECT 257.500000 466.410000 258.500000 467.590000 ;
      RECT 216.500000 466.410000 249.500000 467.590000 ;
      RECT 207.500000 466.410000 208.500000 467.590000 ;
      RECT 166.500000 466.410000 199.500000 467.590000 ;
      RECT 157.500000 466.410000 158.500000 467.590000 ;
      RECT 116.500000 466.410000 149.500000 467.590000 ;
      RECT 107.500000 466.410000 108.500000 467.590000 ;
      RECT 66.500000 466.410000 99.500000 467.590000 ;
      RECT 57.500000 466.410000 58.500000 467.590000 ;
      RECT 29.500000 466.410000 49.500000 467.590000 ;
      RECT 15.500000 466.410000 16.500000 467.590000 ;
      RECT 1157.500000 465.590000 1183.980000 466.410000 ;
      RECT 707.500000 465.590000 723.500000 466.410000 ;
      RECT 657.500000 465.590000 699.500000 466.410000 ;
      RECT 607.500000 465.590000 649.500000 466.410000 ;
      RECT 557.500000 465.590000 599.500000 466.410000 ;
      RECT 507.500000 465.590000 549.500000 466.410000 ;
      RECT 457.500000 465.590000 499.500000 466.410000 ;
      RECT 407.500000 465.590000 449.500000 466.410000 ;
      RECT 357.500000 465.590000 399.500000 466.410000 ;
      RECT 307.500000 465.590000 349.500000 466.410000 ;
      RECT 257.500000 465.590000 299.500000 466.410000 ;
      RECT 207.500000 465.590000 249.500000 466.410000 ;
      RECT 157.500000 465.590000 199.500000 466.410000 ;
      RECT 107.500000 465.590000 149.500000 466.410000 ;
      RECT 57.500000 465.590000 99.500000 466.410000 ;
      RECT 15.500000 465.590000 49.500000 466.410000 ;
      RECT 1157.500000 464.410000 1158.500000 465.590000 ;
      RECT 1139.000000 464.410000 1149.500000 467.590000 ;
      RECT 736.500000 464.410000 739.000000 467.590000 ;
      RECT 722.500000 464.410000 723.500000 465.590000 ;
      RECT 707.500000 464.410000 708.500000 465.590000 ;
      RECT 666.500000 464.410000 699.500000 465.590000 ;
      RECT 657.500000 464.410000 658.500000 465.590000 ;
      RECT 616.500000 464.410000 649.500000 465.590000 ;
      RECT 607.500000 464.410000 608.500000 465.590000 ;
      RECT 566.500000 464.410000 599.500000 465.590000 ;
      RECT 557.500000 464.410000 558.500000 465.590000 ;
      RECT 516.500000 464.410000 549.500000 465.590000 ;
      RECT 507.500000 464.410000 508.500000 465.590000 ;
      RECT 466.500000 464.410000 499.500000 465.590000 ;
      RECT 457.500000 464.410000 458.500000 465.590000 ;
      RECT 416.500000 464.410000 449.500000 465.590000 ;
      RECT 407.500000 464.410000 408.500000 465.590000 ;
      RECT 366.500000 464.410000 399.500000 465.590000 ;
      RECT 357.500000 464.410000 358.500000 465.590000 ;
      RECT 316.500000 464.410000 349.500000 465.590000 ;
      RECT 307.500000 464.410000 308.500000 465.590000 ;
      RECT 266.500000 464.410000 299.500000 465.590000 ;
      RECT 257.500000 464.410000 258.500000 465.590000 ;
      RECT 216.500000 464.410000 249.500000 465.590000 ;
      RECT 207.500000 464.410000 208.500000 465.590000 ;
      RECT 166.500000 464.410000 199.500000 465.590000 ;
      RECT 157.500000 464.410000 158.500000 465.590000 ;
      RECT 116.500000 464.410000 149.500000 465.590000 ;
      RECT 107.500000 464.410000 108.500000 465.590000 ;
      RECT 66.500000 464.410000 99.500000 465.590000 ;
      RECT 57.500000 464.410000 58.500000 465.590000 ;
      RECT 29.500000 464.410000 49.500000 465.590000 ;
      RECT 15.500000 464.410000 16.500000 465.590000 ;
      RECT 2.020000 464.410000 2.500000 466.935000 ;
      RECT 2.020000 463.835000 16.500000 464.410000 ;
      RECT 1166.500000 463.830000 1183.980000 465.590000 ;
      RECT 1139.000000 463.590000 1158.500000 464.410000 ;
      RECT 722.500000 463.590000 739.000000 464.410000 ;
      RECT 666.500000 463.590000 708.500000 464.410000 ;
      RECT 616.500000 463.590000 658.500000 464.410000 ;
      RECT 566.500000 463.590000 608.500000 464.410000 ;
      RECT 516.500000 463.590000 558.500000 464.410000 ;
      RECT 466.500000 463.590000 508.500000 464.410000 ;
      RECT 416.500000 463.590000 458.500000 464.410000 ;
      RECT 366.500000 463.590000 408.500000 464.410000 ;
      RECT 316.500000 463.590000 358.500000 464.410000 ;
      RECT 266.500000 463.590000 308.500000 464.410000 ;
      RECT 216.500000 463.590000 258.500000 464.410000 ;
      RECT 166.500000 463.590000 208.500000 464.410000 ;
      RECT 116.500000 463.590000 158.500000 464.410000 ;
      RECT 66.500000 463.590000 108.500000 464.410000 ;
      RECT 29.500000 463.590000 58.500000 464.410000 ;
      RECT 0.000000 463.590000 16.500000 463.835000 ;
      RECT 1166.500000 462.410000 1186.000000 463.830000 ;
      RECT 1157.500000 462.410000 1158.500000 463.590000 ;
      RECT 722.500000 462.410000 723.500000 463.590000 ;
      RECT 707.500000 462.410000 708.500000 463.590000 ;
      RECT 666.500000 462.410000 699.500000 463.590000 ;
      RECT 657.500000 462.410000 658.500000 463.590000 ;
      RECT 616.500000 462.410000 649.500000 463.590000 ;
      RECT 607.500000 462.410000 608.500000 463.590000 ;
      RECT 566.500000 462.410000 599.500000 463.590000 ;
      RECT 557.500000 462.410000 558.500000 463.590000 ;
      RECT 516.500000 462.410000 549.500000 463.590000 ;
      RECT 507.500000 462.410000 508.500000 463.590000 ;
      RECT 466.500000 462.410000 499.500000 463.590000 ;
      RECT 457.500000 462.410000 458.500000 463.590000 ;
      RECT 416.500000 462.410000 449.500000 463.590000 ;
      RECT 407.500000 462.410000 408.500000 463.590000 ;
      RECT 366.500000 462.410000 399.500000 463.590000 ;
      RECT 357.500000 462.410000 358.500000 463.590000 ;
      RECT 316.500000 462.410000 349.500000 463.590000 ;
      RECT 307.500000 462.410000 308.500000 463.590000 ;
      RECT 266.500000 462.410000 299.500000 463.590000 ;
      RECT 257.500000 462.410000 258.500000 463.590000 ;
      RECT 216.500000 462.410000 249.500000 463.590000 ;
      RECT 207.500000 462.410000 208.500000 463.590000 ;
      RECT 166.500000 462.410000 199.500000 463.590000 ;
      RECT 157.500000 462.410000 158.500000 463.590000 ;
      RECT 116.500000 462.410000 149.500000 463.590000 ;
      RECT 107.500000 462.410000 108.500000 463.590000 ;
      RECT 66.500000 462.410000 99.500000 463.590000 ;
      RECT 57.500000 462.410000 58.500000 463.590000 ;
      RECT 29.500000 462.410000 49.500000 463.590000 ;
      RECT 15.500000 462.410000 16.500000 463.590000 ;
      RECT 1157.500000 461.590000 1186.000000 462.410000 ;
      RECT 707.500000 461.590000 723.500000 462.410000 ;
      RECT 657.500000 461.590000 699.500000 462.410000 ;
      RECT 607.500000 461.590000 649.500000 462.410000 ;
      RECT 557.500000 461.590000 599.500000 462.410000 ;
      RECT 507.500000 461.590000 549.500000 462.410000 ;
      RECT 457.500000 461.590000 499.500000 462.410000 ;
      RECT 407.500000 461.590000 449.500000 462.410000 ;
      RECT 357.500000 461.590000 399.500000 462.410000 ;
      RECT 307.500000 461.590000 349.500000 462.410000 ;
      RECT 207.500000 461.590000 249.500000 462.410000 ;
      RECT 107.500000 461.590000 149.500000 462.410000 ;
      RECT 57.500000 461.590000 99.500000 462.410000 ;
      RECT 15.500000 461.590000 49.500000 462.410000 ;
      RECT 1157.500000 460.410000 1158.500000 461.590000 ;
      RECT 1139.000000 460.410000 1149.500000 463.590000 ;
      RECT 736.500000 460.410000 739.000000 463.590000 ;
      RECT 722.500000 460.410000 723.500000 461.590000 ;
      RECT 707.500000 460.410000 708.500000 461.590000 ;
      RECT 666.500000 460.410000 699.500000 461.590000 ;
      RECT 657.500000 460.410000 658.500000 461.590000 ;
      RECT 616.500000 460.410000 649.500000 461.590000 ;
      RECT 607.500000 460.410000 608.500000 461.590000 ;
      RECT 566.500000 460.410000 599.500000 461.590000 ;
      RECT 557.500000 460.410000 558.500000 461.590000 ;
      RECT 516.500000 460.410000 549.500000 461.590000 ;
      RECT 507.500000 460.410000 508.500000 461.590000 ;
      RECT 466.500000 460.410000 499.500000 461.590000 ;
      RECT 457.500000 460.410000 458.500000 461.590000 ;
      RECT 416.500000 460.410000 449.500000 461.590000 ;
      RECT 407.500000 460.410000 408.500000 461.590000 ;
      RECT 366.500000 460.410000 399.500000 461.590000 ;
      RECT 357.500000 460.410000 358.500000 461.590000 ;
      RECT 316.500000 460.410000 349.500000 461.590000 ;
      RECT 307.500000 460.410000 308.500000 461.590000 ;
      RECT 257.500000 460.410000 299.500000 462.410000 ;
      RECT 216.500000 460.410000 249.500000 461.590000 ;
      RECT 207.500000 460.410000 208.500000 461.590000 ;
      RECT 157.500000 460.410000 199.500000 462.410000 ;
      RECT 116.500000 460.410000 149.500000 461.590000 ;
      RECT 107.500000 460.410000 108.500000 461.590000 ;
      RECT 66.500000 460.410000 99.500000 461.590000 ;
      RECT 57.500000 460.410000 58.500000 461.590000 ;
      RECT 29.500000 460.410000 49.500000 461.590000 ;
      RECT 15.500000 460.410000 16.500000 461.590000 ;
      RECT 0.000000 460.410000 2.500000 463.590000 ;
      RECT 1139.000000 459.590000 1158.500000 460.410000 ;
      RECT 722.500000 459.590000 739.000000 460.410000 ;
      RECT 666.500000 459.590000 708.500000 460.410000 ;
      RECT 616.500000 459.590000 658.500000 460.410000 ;
      RECT 566.500000 459.590000 608.500000 460.410000 ;
      RECT 516.500000 459.590000 558.500000 460.410000 ;
      RECT 466.500000 459.590000 508.500000 460.410000 ;
      RECT 416.500000 459.590000 458.500000 460.410000 ;
      RECT 366.500000 459.590000 408.500000 460.410000 ;
      RECT 316.500000 459.590000 358.500000 460.410000 ;
      RECT 216.500000 459.590000 308.500000 460.410000 ;
      RECT 116.500000 459.590000 208.500000 460.410000 ;
      RECT 66.500000 459.590000 108.500000 460.410000 ;
      RECT 29.500000 459.590000 58.500000 460.410000 ;
      RECT 0.000000 459.590000 16.500000 460.410000 ;
      RECT 1166.500000 458.410000 1186.000000 461.590000 ;
      RECT 1157.500000 458.410000 1158.500000 459.590000 ;
      RECT 722.500000 458.410000 723.500000 459.590000 ;
      RECT 707.500000 458.410000 708.500000 459.590000 ;
      RECT 666.500000 458.410000 699.500000 459.590000 ;
      RECT 657.500000 458.410000 658.500000 459.590000 ;
      RECT 616.500000 458.410000 649.500000 459.590000 ;
      RECT 607.500000 458.410000 608.500000 459.590000 ;
      RECT 566.500000 458.410000 599.500000 459.590000 ;
      RECT 557.500000 458.410000 558.500000 459.590000 ;
      RECT 516.500000 458.410000 549.500000 459.590000 ;
      RECT 507.500000 458.410000 508.500000 459.590000 ;
      RECT 466.500000 458.410000 499.500000 459.590000 ;
      RECT 457.500000 458.410000 458.500000 459.590000 ;
      RECT 416.500000 458.410000 449.500000 459.590000 ;
      RECT 407.500000 458.410000 408.500000 459.590000 ;
      RECT 366.500000 458.410000 399.500000 459.590000 ;
      RECT 357.500000 458.410000 358.500000 459.590000 ;
      RECT 316.500000 458.410000 349.500000 459.590000 ;
      RECT 307.500000 458.410000 308.500000 459.590000 ;
      RECT 216.500000 458.410000 249.500000 459.590000 ;
      RECT 207.500000 458.410000 208.500000 459.590000 ;
      RECT 116.500000 458.410000 149.500000 459.590000 ;
      RECT 107.500000 458.410000 108.500000 459.590000 ;
      RECT 66.500000 458.410000 99.500000 459.590000 ;
      RECT 57.500000 458.410000 58.500000 459.590000 ;
      RECT 29.500000 458.410000 49.500000 459.590000 ;
      RECT 15.500000 458.410000 16.500000 459.590000 ;
      RECT 1157.500000 457.590000 1186.000000 458.410000 ;
      RECT 707.500000 457.590000 723.500000 458.410000 ;
      RECT 657.500000 457.590000 699.500000 458.410000 ;
      RECT 607.500000 457.590000 649.500000 458.410000 ;
      RECT 557.500000 457.590000 599.500000 458.410000 ;
      RECT 507.500000 457.590000 549.500000 458.410000 ;
      RECT 457.500000 457.590000 499.500000 458.410000 ;
      RECT 407.500000 457.590000 449.500000 458.410000 ;
      RECT 357.500000 457.590000 399.500000 458.410000 ;
      RECT 307.500000 457.590000 349.500000 458.410000 ;
      RECT 207.500000 457.590000 249.500000 458.410000 ;
      RECT 107.500000 457.590000 149.500000 458.410000 ;
      RECT 57.500000 457.590000 99.500000 458.410000 ;
      RECT 15.500000 457.590000 49.500000 458.410000 ;
      RECT 1157.500000 456.410000 1158.500000 457.590000 ;
      RECT 1139.000000 456.410000 1149.500000 459.590000 ;
      RECT 736.500000 456.410000 739.000000 459.590000 ;
      RECT 722.500000 456.410000 723.500000 457.590000 ;
      RECT 707.500000 456.410000 708.500000 457.590000 ;
      RECT 666.500000 456.410000 699.500000 457.590000 ;
      RECT 657.500000 456.410000 658.500000 457.590000 ;
      RECT 616.500000 456.410000 649.500000 457.590000 ;
      RECT 607.500000 456.410000 608.500000 457.590000 ;
      RECT 566.500000 456.410000 599.500000 457.590000 ;
      RECT 557.500000 456.410000 558.500000 457.590000 ;
      RECT 516.500000 456.410000 549.500000 457.590000 ;
      RECT 507.500000 456.410000 508.500000 457.590000 ;
      RECT 466.500000 456.410000 499.500000 457.590000 ;
      RECT 457.500000 456.410000 458.500000 457.590000 ;
      RECT 416.500000 456.410000 449.500000 457.590000 ;
      RECT 407.500000 456.410000 408.500000 457.590000 ;
      RECT 366.500000 456.410000 399.500000 457.590000 ;
      RECT 357.500000 456.410000 358.500000 457.590000 ;
      RECT 316.500000 456.410000 349.500000 457.590000 ;
      RECT 307.500000 456.410000 308.500000 457.590000 ;
      RECT 257.500000 456.410000 299.500000 459.590000 ;
      RECT 216.500000 456.410000 249.500000 457.590000 ;
      RECT 207.500000 456.410000 208.500000 457.590000 ;
      RECT 157.500000 456.410000 199.500000 459.590000 ;
      RECT 116.500000 456.410000 149.500000 457.590000 ;
      RECT 107.500000 456.410000 108.500000 457.590000 ;
      RECT 66.500000 456.410000 99.500000 457.590000 ;
      RECT 57.500000 456.410000 58.500000 457.590000 ;
      RECT 29.500000 456.410000 49.500000 457.590000 ;
      RECT 15.500000 456.410000 16.500000 457.590000 ;
      RECT 0.000000 456.410000 2.500000 459.590000 ;
      RECT 1139.000000 455.590000 1158.500000 456.410000 ;
      RECT 722.500000 455.590000 739.000000 456.410000 ;
      RECT 666.500000 455.590000 708.500000 456.410000 ;
      RECT 616.500000 455.590000 658.500000 456.410000 ;
      RECT 566.500000 455.590000 608.500000 456.410000 ;
      RECT 516.500000 455.590000 558.500000 456.410000 ;
      RECT 466.500000 455.590000 508.500000 456.410000 ;
      RECT 416.500000 455.590000 458.500000 456.410000 ;
      RECT 366.500000 455.590000 408.500000 456.410000 ;
      RECT 316.500000 455.590000 358.500000 456.410000 ;
      RECT 216.500000 455.590000 308.500000 456.410000 ;
      RECT 116.500000 455.590000 208.500000 456.410000 ;
      RECT 66.500000 455.590000 108.500000 456.410000 ;
      RECT 29.500000 455.590000 58.500000 456.410000 ;
      RECT 0.000000 455.590000 16.500000 456.410000 ;
      RECT 1166.500000 454.410000 1186.000000 457.590000 ;
      RECT 1157.500000 454.410000 1158.500000 455.590000 ;
      RECT 722.500000 454.410000 723.500000 455.590000 ;
      RECT 707.500000 454.410000 708.500000 455.590000 ;
      RECT 666.500000 454.410000 699.500000 455.590000 ;
      RECT 657.500000 454.410000 658.500000 455.590000 ;
      RECT 616.500000 454.410000 649.500000 455.590000 ;
      RECT 607.500000 454.410000 608.500000 455.590000 ;
      RECT 566.500000 454.410000 599.500000 455.590000 ;
      RECT 557.500000 454.410000 558.500000 455.590000 ;
      RECT 516.500000 454.410000 549.500000 455.590000 ;
      RECT 507.500000 454.410000 508.500000 455.590000 ;
      RECT 466.500000 454.410000 499.500000 455.590000 ;
      RECT 457.500000 454.410000 458.500000 455.590000 ;
      RECT 416.500000 454.410000 449.500000 455.590000 ;
      RECT 407.500000 454.410000 408.500000 455.590000 ;
      RECT 366.500000 454.410000 399.500000 455.590000 ;
      RECT 357.500000 454.410000 358.500000 455.590000 ;
      RECT 316.500000 454.410000 349.500000 455.590000 ;
      RECT 307.500000 454.410000 308.500000 455.590000 ;
      RECT 216.500000 454.410000 249.500000 455.590000 ;
      RECT 207.500000 454.410000 208.500000 455.590000 ;
      RECT 116.500000 454.410000 149.500000 455.590000 ;
      RECT 107.500000 454.410000 108.500000 455.590000 ;
      RECT 66.500000 454.410000 99.500000 455.590000 ;
      RECT 57.500000 454.410000 58.500000 455.590000 ;
      RECT 29.500000 454.410000 49.500000 455.590000 ;
      RECT 15.500000 454.410000 16.500000 455.590000 ;
      RECT 1157.500000 453.590000 1186.000000 454.410000 ;
      RECT 707.500000 453.590000 723.500000 454.410000 ;
      RECT 657.500000 453.590000 699.500000 454.410000 ;
      RECT 607.500000 453.590000 649.500000 454.410000 ;
      RECT 557.500000 453.590000 599.500000 454.410000 ;
      RECT 507.500000 453.590000 549.500000 454.410000 ;
      RECT 457.500000 453.590000 499.500000 454.410000 ;
      RECT 407.500000 453.590000 449.500000 454.410000 ;
      RECT 357.500000 453.590000 399.500000 454.410000 ;
      RECT 307.500000 453.590000 349.500000 454.410000 ;
      RECT 207.500000 453.590000 249.500000 454.410000 ;
      RECT 107.500000 453.590000 149.500000 454.410000 ;
      RECT 57.500000 453.590000 99.500000 454.410000 ;
      RECT 15.500000 453.590000 49.500000 454.410000 ;
      RECT 1157.500000 452.410000 1158.500000 453.590000 ;
      RECT 1139.000000 452.410000 1149.500000 455.590000 ;
      RECT 736.500000 452.410000 739.000000 455.590000 ;
      RECT 722.500000 452.410000 723.500000 453.590000 ;
      RECT 707.500000 452.410000 708.500000 453.590000 ;
      RECT 666.500000 452.410000 699.500000 453.590000 ;
      RECT 657.500000 452.410000 658.500000 453.590000 ;
      RECT 616.500000 452.410000 649.500000 453.590000 ;
      RECT 607.500000 452.410000 608.500000 453.590000 ;
      RECT 566.500000 452.410000 599.500000 453.590000 ;
      RECT 557.500000 452.410000 558.500000 453.590000 ;
      RECT 516.500000 452.410000 549.500000 453.590000 ;
      RECT 507.500000 452.410000 508.500000 453.590000 ;
      RECT 466.500000 452.410000 499.500000 453.590000 ;
      RECT 457.500000 452.410000 458.500000 453.590000 ;
      RECT 416.500000 452.410000 449.500000 453.590000 ;
      RECT 407.500000 452.410000 408.500000 453.590000 ;
      RECT 366.500000 452.410000 399.500000 453.590000 ;
      RECT 357.500000 452.410000 358.500000 453.590000 ;
      RECT 316.500000 452.410000 349.500000 453.590000 ;
      RECT 307.500000 452.410000 308.500000 453.590000 ;
      RECT 257.500000 452.410000 299.500000 455.590000 ;
      RECT 216.500000 452.410000 249.500000 453.590000 ;
      RECT 207.500000 452.410000 208.500000 453.590000 ;
      RECT 157.500000 452.410000 199.500000 455.590000 ;
      RECT 116.500000 452.410000 149.500000 453.590000 ;
      RECT 107.500000 452.410000 108.500000 453.590000 ;
      RECT 66.500000 452.410000 99.500000 453.590000 ;
      RECT 57.500000 452.410000 58.500000 453.590000 ;
      RECT 29.500000 452.410000 49.500000 453.590000 ;
      RECT 15.500000 452.410000 16.500000 453.590000 ;
      RECT 0.000000 452.410000 2.500000 455.590000 ;
      RECT 1139.000000 451.590000 1158.500000 452.410000 ;
      RECT 722.500000 451.590000 739.000000 452.410000 ;
      RECT 666.500000 451.590000 708.500000 452.410000 ;
      RECT 616.500000 451.590000 658.500000 452.410000 ;
      RECT 566.500000 451.590000 608.500000 452.410000 ;
      RECT 516.500000 451.590000 558.500000 452.410000 ;
      RECT 466.500000 451.590000 508.500000 452.410000 ;
      RECT 416.500000 451.590000 458.500000 452.410000 ;
      RECT 366.500000 451.590000 408.500000 452.410000 ;
      RECT 316.500000 451.590000 358.500000 452.410000 ;
      RECT 216.500000 451.590000 308.500000 452.410000 ;
      RECT 116.500000 451.590000 208.500000 452.410000 ;
      RECT 66.500000 451.590000 108.500000 452.410000 ;
      RECT 29.500000 451.590000 58.500000 452.410000 ;
      RECT 0.000000 451.590000 16.500000 452.410000 ;
      RECT 1166.500000 450.410000 1186.000000 453.590000 ;
      RECT 1157.500000 450.410000 1158.500000 451.590000 ;
      RECT 722.500000 450.410000 723.500000 451.590000 ;
      RECT 707.500000 450.410000 708.500000 451.590000 ;
      RECT 666.500000 450.410000 699.500000 451.590000 ;
      RECT 657.500000 450.410000 658.500000 451.590000 ;
      RECT 616.500000 450.410000 649.500000 451.590000 ;
      RECT 607.500000 450.410000 608.500000 451.590000 ;
      RECT 566.500000 450.410000 599.500000 451.590000 ;
      RECT 557.500000 450.410000 558.500000 451.590000 ;
      RECT 516.500000 450.410000 549.500000 451.590000 ;
      RECT 507.500000 450.410000 508.500000 451.590000 ;
      RECT 466.500000 450.410000 499.500000 451.590000 ;
      RECT 457.500000 450.410000 458.500000 451.590000 ;
      RECT 416.500000 450.410000 449.500000 451.590000 ;
      RECT 407.500000 450.410000 408.500000 451.590000 ;
      RECT 366.500000 450.410000 399.500000 451.590000 ;
      RECT 357.500000 450.410000 358.500000 451.590000 ;
      RECT 316.500000 450.410000 349.500000 451.590000 ;
      RECT 307.500000 450.410000 308.500000 451.590000 ;
      RECT 216.500000 450.410000 299.500000 451.590000 ;
      RECT 207.500000 450.410000 208.500000 451.590000 ;
      RECT 116.500000 450.410000 199.500000 451.590000 ;
      RECT 107.500000 450.410000 108.500000 451.590000 ;
      RECT 66.500000 450.410000 99.500000 451.590000 ;
      RECT 57.500000 450.410000 58.500000 451.590000 ;
      RECT 29.500000 450.410000 49.500000 451.590000 ;
      RECT 15.500000 450.410000 16.500000 451.590000 ;
      RECT 1157.500000 449.590000 1186.000000 450.410000 ;
      RECT 707.500000 449.590000 723.500000 450.410000 ;
      RECT 657.500000 449.590000 699.500000 450.410000 ;
      RECT 607.500000 449.590000 649.500000 450.410000 ;
      RECT 557.500000 449.590000 599.500000 450.410000 ;
      RECT 507.500000 449.590000 549.500000 450.410000 ;
      RECT 457.500000 449.590000 499.500000 450.410000 ;
      RECT 407.500000 449.590000 449.500000 450.410000 ;
      RECT 357.500000 449.590000 399.500000 450.410000 ;
      RECT 307.500000 449.590000 349.500000 450.410000 ;
      RECT 207.500000 449.590000 299.500000 450.410000 ;
      RECT 107.500000 449.590000 199.500000 450.410000 ;
      RECT 57.500000 449.590000 99.500000 450.410000 ;
      RECT 15.500000 449.590000 49.500000 450.410000 ;
      RECT 1157.500000 448.410000 1158.500000 449.590000 ;
      RECT 1139.000000 448.410000 1149.500000 451.590000 ;
      RECT 736.500000 448.410000 739.000000 451.590000 ;
      RECT 722.500000 448.410000 723.500000 449.590000 ;
      RECT 707.500000 448.410000 708.500000 449.590000 ;
      RECT 666.500000 448.410000 699.500000 449.590000 ;
      RECT 657.500000 448.410000 658.500000 449.590000 ;
      RECT 616.500000 448.410000 649.500000 449.590000 ;
      RECT 607.500000 448.410000 608.500000 449.590000 ;
      RECT 566.500000 448.410000 599.500000 449.590000 ;
      RECT 557.500000 448.410000 558.500000 449.590000 ;
      RECT 516.500000 448.410000 549.500000 449.590000 ;
      RECT 507.500000 448.410000 508.500000 449.590000 ;
      RECT 466.500000 448.410000 499.500000 449.590000 ;
      RECT 457.500000 448.410000 458.500000 449.590000 ;
      RECT 416.500000 448.410000 449.500000 449.590000 ;
      RECT 407.500000 448.410000 408.500000 449.590000 ;
      RECT 366.500000 448.410000 399.500000 449.590000 ;
      RECT 357.500000 448.410000 358.500000 449.590000 ;
      RECT 316.500000 448.410000 349.500000 449.590000 ;
      RECT 307.500000 448.410000 308.500000 449.590000 ;
      RECT 216.500000 448.410000 299.500000 449.590000 ;
      RECT 207.500000 448.410000 208.500000 449.590000 ;
      RECT 116.500000 448.410000 199.500000 449.590000 ;
      RECT 107.500000 448.410000 108.500000 449.590000 ;
      RECT 66.500000 448.410000 99.500000 449.590000 ;
      RECT 57.500000 448.410000 58.500000 449.590000 ;
      RECT 29.500000 448.410000 49.500000 449.590000 ;
      RECT 15.500000 448.410000 16.500000 449.590000 ;
      RECT 0.000000 448.410000 2.500000 451.590000 ;
      RECT 1139.000000 447.590000 1158.500000 448.410000 ;
      RECT 722.500000 447.590000 739.000000 448.410000 ;
      RECT 666.500000 447.590000 708.500000 448.410000 ;
      RECT 616.500000 447.590000 658.500000 448.410000 ;
      RECT 566.500000 447.590000 608.500000 448.410000 ;
      RECT 516.500000 447.590000 558.500000 448.410000 ;
      RECT 466.500000 447.590000 508.500000 448.410000 ;
      RECT 416.500000 447.590000 458.500000 448.410000 ;
      RECT 366.500000 447.590000 408.500000 448.410000 ;
      RECT 316.500000 447.590000 358.500000 448.410000 ;
      RECT 216.500000 447.590000 308.500000 448.410000 ;
      RECT 116.500000 447.590000 208.500000 448.410000 ;
      RECT 66.500000 447.590000 108.500000 448.410000 ;
      RECT 29.500000 447.590000 58.500000 448.410000 ;
      RECT 0.000000 447.590000 16.500000 448.410000 ;
      RECT 1166.500000 446.410000 1186.000000 449.590000 ;
      RECT 1157.500000 446.410000 1158.500000 447.590000 ;
      RECT 722.500000 446.410000 723.500000 447.590000 ;
      RECT 707.500000 446.410000 708.500000 447.590000 ;
      RECT 666.500000 446.410000 699.500000 447.590000 ;
      RECT 657.500000 446.410000 658.500000 447.590000 ;
      RECT 616.500000 446.410000 649.500000 447.590000 ;
      RECT 607.500000 446.410000 608.500000 447.590000 ;
      RECT 566.500000 446.410000 599.500000 447.590000 ;
      RECT 557.500000 446.410000 558.500000 447.590000 ;
      RECT 516.500000 446.410000 549.500000 447.590000 ;
      RECT 507.500000 446.410000 508.500000 447.590000 ;
      RECT 466.500000 446.410000 499.500000 447.590000 ;
      RECT 457.500000 446.410000 458.500000 447.590000 ;
      RECT 416.500000 446.410000 449.500000 447.590000 ;
      RECT 407.500000 446.410000 408.500000 447.590000 ;
      RECT 366.500000 446.410000 399.500000 447.590000 ;
      RECT 357.500000 446.410000 358.500000 447.590000 ;
      RECT 316.500000 446.410000 349.500000 447.590000 ;
      RECT 307.500000 446.410000 308.500000 447.590000 ;
      RECT 216.500000 446.410000 299.500000 447.590000 ;
      RECT 207.500000 446.410000 208.500000 447.590000 ;
      RECT 116.500000 446.410000 199.500000 447.590000 ;
      RECT 107.500000 446.410000 108.500000 447.590000 ;
      RECT 66.500000 446.410000 99.500000 447.590000 ;
      RECT 57.500000 446.410000 58.500000 447.590000 ;
      RECT 29.500000 446.410000 49.500000 447.590000 ;
      RECT 15.500000 446.410000 16.500000 447.590000 ;
      RECT 1139.000000 446.000000 1149.500000 447.590000 ;
      RECT 736.500000 446.000000 739.000000 447.590000 ;
      RECT 1157.500000 445.590000 1186.000000 446.410000 ;
      RECT 1060.750000 445.590000 1149.500000 446.000000 ;
      RECT 999.630000 445.590000 1009.115000 446.000000 ;
      RECT 876.205000 445.590000 996.530000 446.000000 ;
      RECT 736.500000 445.590000 868.305000 446.000000 ;
      RECT 707.500000 445.590000 723.500000 446.410000 ;
      RECT 657.500000 445.590000 699.500000 446.410000 ;
      RECT 607.500000 445.590000 649.500000 446.410000 ;
      RECT 557.500000 445.590000 599.500000 446.410000 ;
      RECT 507.500000 445.590000 549.500000 446.410000 ;
      RECT 457.500000 445.590000 499.500000 446.410000 ;
      RECT 407.500000 445.590000 449.500000 446.410000 ;
      RECT 357.500000 445.590000 399.500000 446.410000 ;
      RECT 307.500000 445.590000 349.500000 446.410000 ;
      RECT 207.500000 445.590000 299.500000 446.410000 ;
      RECT 107.500000 445.590000 199.500000 446.410000 ;
      RECT 57.500000 445.590000 99.500000 446.410000 ;
      RECT 15.500000 445.590000 49.500000 446.410000 ;
      RECT 1157.500000 444.410000 1158.500000 445.590000 ;
      RECT 1116.500000 444.410000 1149.500000 445.590000 ;
      RECT 736.500000 444.410000 758.500000 445.590000 ;
      RECT 722.500000 444.410000 723.500000 445.590000 ;
      RECT 707.500000 444.410000 708.500000 445.590000 ;
      RECT 666.500000 444.410000 699.500000 445.590000 ;
      RECT 657.500000 444.410000 658.500000 445.590000 ;
      RECT 616.500000 444.410000 649.500000 445.590000 ;
      RECT 607.500000 444.410000 608.500000 445.590000 ;
      RECT 566.500000 444.410000 599.500000 445.590000 ;
      RECT 557.500000 444.410000 558.500000 445.590000 ;
      RECT 516.500000 444.410000 549.500000 445.590000 ;
      RECT 507.500000 444.410000 508.500000 445.590000 ;
      RECT 466.500000 444.410000 499.500000 445.590000 ;
      RECT 457.500000 444.410000 458.500000 445.590000 ;
      RECT 416.500000 444.410000 449.500000 445.590000 ;
      RECT 407.500000 444.410000 408.500000 445.590000 ;
      RECT 366.500000 444.410000 399.500000 445.590000 ;
      RECT 357.500000 444.410000 358.500000 445.590000 ;
      RECT 316.500000 444.410000 349.500000 445.590000 ;
      RECT 307.500000 444.410000 308.500000 445.590000 ;
      RECT 216.500000 444.410000 299.500000 445.590000 ;
      RECT 207.500000 444.410000 208.500000 445.590000 ;
      RECT 116.500000 444.410000 199.500000 445.590000 ;
      RECT 107.500000 444.410000 108.500000 445.590000 ;
      RECT 66.500000 444.410000 99.500000 445.590000 ;
      RECT 57.500000 444.410000 58.500000 445.590000 ;
      RECT 29.500000 444.410000 49.500000 445.590000 ;
      RECT 15.500000 444.410000 16.500000 445.590000 ;
      RECT 0.000000 444.410000 2.500000 447.590000 ;
      RECT 1029.110000 443.980000 1040.755000 446.000000 ;
      RECT 999.630000 443.980000 1008.500000 445.590000 ;
      RECT 966.500000 443.980000 996.530000 445.590000 ;
      RECT 876.205000 443.980000 908.500000 445.590000 ;
      RECT 866.500000 443.980000 868.305000 445.590000 ;
      RECT 1166.500000 443.590000 1186.000000 445.590000 ;
      RECT 1116.500000 443.590000 1158.500000 444.410000 ;
      RECT 1066.500000 443.590000 1108.500000 445.590000 ;
      RECT 1016.500000 443.590000 1058.500000 443.980000 ;
      RECT 966.500000 443.590000 1008.500000 443.980000 ;
      RECT 916.500000 443.590000 958.500000 445.590000 ;
      RECT 866.500000 443.590000 908.500000 443.980000 ;
      RECT 816.500000 443.590000 858.500000 445.590000 ;
      RECT 766.500000 443.590000 808.500000 445.590000 ;
      RECT 722.500000 443.590000 758.500000 444.410000 ;
      RECT 666.500000 443.590000 708.500000 444.410000 ;
      RECT 616.500000 443.590000 658.500000 444.410000 ;
      RECT 566.500000 443.590000 608.500000 444.410000 ;
      RECT 516.500000 443.590000 558.500000 444.410000 ;
      RECT 466.500000 443.590000 508.500000 444.410000 ;
      RECT 416.500000 443.590000 458.500000 444.410000 ;
      RECT 366.500000 443.590000 408.500000 444.410000 ;
      RECT 316.500000 443.590000 358.500000 444.410000 ;
      RECT 216.500000 443.590000 308.500000 444.410000 ;
      RECT 116.500000 443.590000 208.500000 444.410000 ;
      RECT 66.500000 443.590000 108.500000 444.410000 ;
      RECT 29.500000 443.590000 58.500000 444.410000 ;
      RECT 0.000000 443.590000 16.500000 444.410000 ;
      RECT 1166.500000 442.410000 1170.500000 443.590000 ;
      RECT 1157.500000 442.410000 1158.500000 443.590000 ;
      RECT 1116.500000 442.410000 1149.500000 443.590000 ;
      RECT 1107.500000 442.410000 1108.500000 443.590000 ;
      RECT 1066.500000 442.410000 1099.500000 443.590000 ;
      RECT 1057.500000 442.410000 1058.500000 443.590000 ;
      RECT 1016.500000 442.410000 1049.500000 443.590000 ;
      RECT 1007.500000 442.410000 1008.500000 443.590000 ;
      RECT 966.500000 442.410000 999.500000 443.590000 ;
      RECT 957.500000 442.410000 958.500000 443.590000 ;
      RECT 916.500000 442.410000 949.500000 443.590000 ;
      RECT 907.500000 442.410000 908.500000 443.590000 ;
      RECT 866.500000 442.410000 899.500000 443.590000 ;
      RECT 857.500000 442.410000 858.500000 443.590000 ;
      RECT 816.500000 442.410000 849.500000 443.590000 ;
      RECT 807.500000 442.410000 808.500000 443.590000 ;
      RECT 766.500000 442.410000 799.500000 443.590000 ;
      RECT 757.500000 442.410000 758.500000 443.590000 ;
      RECT 722.500000 442.410000 723.500000 443.590000 ;
      RECT 707.500000 442.410000 708.500000 443.590000 ;
      RECT 666.500000 442.410000 699.500000 443.590000 ;
      RECT 657.500000 442.410000 658.500000 443.590000 ;
      RECT 616.500000 442.410000 649.500000 443.590000 ;
      RECT 607.500000 442.410000 608.500000 443.590000 ;
      RECT 566.500000 442.410000 599.500000 443.590000 ;
      RECT 557.500000 442.410000 558.500000 443.590000 ;
      RECT 516.500000 442.410000 549.500000 443.590000 ;
      RECT 507.500000 442.410000 508.500000 443.590000 ;
      RECT 466.500000 442.410000 499.500000 443.590000 ;
      RECT 457.500000 442.410000 458.500000 443.590000 ;
      RECT 416.500000 442.410000 449.500000 443.590000 ;
      RECT 407.500000 442.410000 408.500000 443.590000 ;
      RECT 366.500000 442.410000 399.500000 443.590000 ;
      RECT 357.500000 442.410000 358.500000 443.590000 ;
      RECT 316.500000 442.410000 349.500000 443.590000 ;
      RECT 307.500000 442.410000 308.500000 443.590000 ;
      RECT 216.500000 442.410000 299.500000 443.590000 ;
      RECT 207.500000 442.410000 208.500000 443.590000 ;
      RECT 116.500000 442.410000 199.500000 443.590000 ;
      RECT 107.500000 442.410000 108.500000 443.590000 ;
      RECT 66.500000 442.410000 99.500000 443.590000 ;
      RECT 57.500000 442.410000 58.500000 443.590000 ;
      RECT 29.500000 442.410000 49.500000 443.590000 ;
      RECT 15.500000 442.410000 16.500000 443.590000 ;
      RECT 1157.500000 441.590000 1170.500000 442.410000 ;
      RECT 1107.500000 441.590000 1149.500000 442.410000 ;
      RECT 1057.500000 441.590000 1099.500000 442.410000 ;
      RECT 1007.500000 441.590000 1049.500000 442.410000 ;
      RECT 957.500000 441.590000 999.500000 442.410000 ;
      RECT 907.500000 441.590000 949.500000 442.410000 ;
      RECT 857.500000 441.590000 899.500000 442.410000 ;
      RECT 807.500000 441.590000 849.500000 442.410000 ;
      RECT 757.500000 441.590000 799.500000 442.410000 ;
      RECT 707.500000 441.590000 723.500000 442.410000 ;
      RECT 657.500000 441.590000 699.500000 442.410000 ;
      RECT 607.500000 441.590000 649.500000 442.410000 ;
      RECT 557.500000 441.590000 599.500000 442.410000 ;
      RECT 507.500000 441.590000 549.500000 442.410000 ;
      RECT 457.500000 441.590000 499.500000 442.410000 ;
      RECT 407.500000 441.590000 449.500000 442.410000 ;
      RECT 357.500000 441.590000 399.500000 442.410000 ;
      RECT 307.500000 441.590000 349.500000 442.410000 ;
      RECT 207.500000 441.590000 299.500000 442.410000 ;
      RECT 107.500000 441.590000 199.500000 442.410000 ;
      RECT 57.500000 441.590000 99.500000 442.410000 ;
      RECT 15.500000 441.590000 49.500000 442.410000 ;
      RECT 1183.500000 440.410000 1186.000000 443.590000 ;
      RECT 1166.500000 440.410000 1170.500000 441.590000 ;
      RECT 1157.500000 440.410000 1158.500000 441.590000 ;
      RECT 1116.500000 440.410000 1149.500000 441.590000 ;
      RECT 1107.500000 440.410000 1108.500000 441.590000 ;
      RECT 1066.500000 440.410000 1099.500000 441.590000 ;
      RECT 1057.500000 440.410000 1058.500000 441.590000 ;
      RECT 1016.500000 440.410000 1049.500000 441.590000 ;
      RECT 1007.500000 440.410000 1008.500000 441.590000 ;
      RECT 966.500000 440.410000 999.500000 441.590000 ;
      RECT 957.500000 440.410000 958.500000 441.590000 ;
      RECT 916.500000 440.410000 949.500000 441.590000 ;
      RECT 907.500000 440.410000 908.500000 441.590000 ;
      RECT 866.500000 440.410000 899.500000 441.590000 ;
      RECT 857.500000 440.410000 858.500000 441.590000 ;
      RECT 816.500000 440.410000 849.500000 441.590000 ;
      RECT 807.500000 440.410000 808.500000 441.590000 ;
      RECT 766.500000 440.410000 799.500000 441.590000 ;
      RECT 757.500000 440.410000 758.500000 441.590000 ;
      RECT 736.500000 440.410000 749.500000 443.590000 ;
      RECT 722.500000 440.410000 723.500000 441.590000 ;
      RECT 707.500000 440.410000 708.500000 441.590000 ;
      RECT 666.500000 440.410000 699.500000 441.590000 ;
      RECT 657.500000 440.410000 658.500000 441.590000 ;
      RECT 616.500000 440.410000 649.500000 441.590000 ;
      RECT 607.500000 440.410000 608.500000 441.590000 ;
      RECT 566.500000 440.410000 599.500000 441.590000 ;
      RECT 557.500000 440.410000 558.500000 441.590000 ;
      RECT 516.500000 440.410000 549.500000 441.590000 ;
      RECT 507.500000 440.410000 508.500000 441.590000 ;
      RECT 466.500000 440.410000 499.500000 441.590000 ;
      RECT 457.500000 440.410000 458.500000 441.590000 ;
      RECT 416.500000 440.410000 449.500000 441.590000 ;
      RECT 407.500000 440.410000 408.500000 441.590000 ;
      RECT 366.500000 440.410000 399.500000 441.590000 ;
      RECT 357.500000 440.410000 358.500000 441.590000 ;
      RECT 316.500000 440.410000 349.500000 441.590000 ;
      RECT 307.500000 440.410000 308.500000 441.590000 ;
      RECT 216.500000 440.410000 299.500000 441.590000 ;
      RECT 207.500000 440.410000 208.500000 441.590000 ;
      RECT 116.500000 440.410000 199.500000 441.590000 ;
      RECT 107.500000 440.410000 108.500000 441.590000 ;
      RECT 66.500000 440.410000 99.500000 441.590000 ;
      RECT 57.500000 440.410000 58.500000 441.590000 ;
      RECT 29.500000 440.410000 49.500000 441.590000 ;
      RECT 15.500000 440.410000 16.500000 441.590000 ;
      RECT 0.000000 440.410000 2.500000 443.590000 ;
      RECT 1166.500000 439.590000 1186.000000 440.410000 ;
      RECT 1116.500000 439.590000 1158.500000 440.410000 ;
      RECT 1066.500000 439.590000 1108.500000 440.410000 ;
      RECT 1016.500000 439.590000 1058.500000 440.410000 ;
      RECT 966.500000 439.590000 1008.500000 440.410000 ;
      RECT 916.500000 439.590000 958.500000 440.410000 ;
      RECT 866.500000 439.590000 908.500000 440.410000 ;
      RECT 816.500000 439.590000 858.500000 440.410000 ;
      RECT 766.500000 439.590000 808.500000 440.410000 ;
      RECT 722.500000 439.590000 758.500000 440.410000 ;
      RECT 666.500000 439.590000 708.500000 440.410000 ;
      RECT 616.500000 439.590000 658.500000 440.410000 ;
      RECT 566.500000 439.590000 608.500000 440.410000 ;
      RECT 516.500000 439.590000 558.500000 440.410000 ;
      RECT 466.500000 439.590000 508.500000 440.410000 ;
      RECT 416.500000 439.590000 458.500000 440.410000 ;
      RECT 366.500000 439.590000 408.500000 440.410000 ;
      RECT 316.500000 439.590000 358.500000 440.410000 ;
      RECT 216.500000 439.590000 308.500000 440.410000 ;
      RECT 116.500000 439.590000 208.500000 440.410000 ;
      RECT 66.500000 439.590000 108.500000 440.410000 ;
      RECT 29.500000 439.590000 58.500000 440.410000 ;
      RECT 0.000000 439.590000 16.500000 440.410000 ;
      RECT 1166.500000 438.410000 1170.500000 439.590000 ;
      RECT 1157.500000 438.410000 1158.500000 439.590000 ;
      RECT 1116.500000 438.410000 1149.500000 439.590000 ;
      RECT 1107.500000 438.410000 1108.500000 439.590000 ;
      RECT 1066.500000 438.410000 1099.500000 439.590000 ;
      RECT 1057.500000 438.410000 1058.500000 439.590000 ;
      RECT 1016.500000 438.410000 1049.500000 439.590000 ;
      RECT 1007.500000 438.410000 1008.500000 439.590000 ;
      RECT 966.500000 438.410000 999.500000 439.590000 ;
      RECT 957.500000 438.410000 958.500000 439.590000 ;
      RECT 916.500000 438.410000 949.500000 439.590000 ;
      RECT 907.500000 438.410000 908.500000 439.590000 ;
      RECT 866.500000 438.410000 899.500000 439.590000 ;
      RECT 857.500000 438.410000 858.500000 439.590000 ;
      RECT 816.500000 438.410000 849.500000 439.590000 ;
      RECT 807.500000 438.410000 808.500000 439.590000 ;
      RECT 766.500000 438.410000 799.500000 439.590000 ;
      RECT 757.500000 438.410000 758.500000 439.590000 ;
      RECT 722.500000 438.410000 723.500000 439.590000 ;
      RECT 707.500000 438.410000 708.500000 439.590000 ;
      RECT 666.500000 438.410000 699.500000 439.590000 ;
      RECT 657.500000 438.410000 658.500000 439.590000 ;
      RECT 616.500000 438.410000 649.500000 439.590000 ;
      RECT 607.500000 438.410000 608.500000 439.590000 ;
      RECT 566.500000 438.410000 599.500000 439.590000 ;
      RECT 557.500000 438.410000 558.500000 439.590000 ;
      RECT 516.500000 438.410000 549.500000 439.590000 ;
      RECT 507.500000 438.410000 508.500000 439.590000 ;
      RECT 466.500000 438.410000 499.500000 439.590000 ;
      RECT 457.500000 438.410000 458.500000 439.590000 ;
      RECT 416.500000 438.410000 449.500000 439.590000 ;
      RECT 407.500000 438.410000 408.500000 439.590000 ;
      RECT 366.500000 438.410000 399.500000 439.590000 ;
      RECT 357.500000 438.410000 358.500000 439.590000 ;
      RECT 316.500000 438.410000 349.500000 439.590000 ;
      RECT 307.500000 438.410000 308.500000 439.590000 ;
      RECT 216.500000 438.410000 299.500000 439.590000 ;
      RECT 207.500000 438.410000 208.500000 439.590000 ;
      RECT 116.500000 438.410000 199.500000 439.590000 ;
      RECT 107.500000 438.410000 108.500000 439.590000 ;
      RECT 66.500000 438.410000 99.500000 439.590000 ;
      RECT 57.500000 438.410000 58.500000 439.590000 ;
      RECT 29.500000 438.410000 49.500000 439.590000 ;
      RECT 15.500000 438.410000 16.500000 439.590000 ;
      RECT 1157.500000 437.590000 1170.500000 438.410000 ;
      RECT 1107.500000 437.590000 1149.500000 438.410000 ;
      RECT 1057.500000 437.590000 1099.500000 438.410000 ;
      RECT 1007.500000 437.590000 1049.500000 438.410000 ;
      RECT 957.500000 437.590000 999.500000 438.410000 ;
      RECT 907.500000 437.590000 949.500000 438.410000 ;
      RECT 857.500000 437.590000 899.500000 438.410000 ;
      RECT 807.500000 437.590000 849.500000 438.410000 ;
      RECT 757.500000 437.590000 799.500000 438.410000 ;
      RECT 707.500000 437.590000 723.500000 438.410000 ;
      RECT 657.500000 437.590000 699.500000 438.410000 ;
      RECT 607.500000 437.590000 649.500000 438.410000 ;
      RECT 557.500000 437.590000 599.500000 438.410000 ;
      RECT 507.500000 437.590000 549.500000 438.410000 ;
      RECT 457.500000 437.590000 499.500000 438.410000 ;
      RECT 407.500000 437.590000 449.500000 438.410000 ;
      RECT 357.500000 437.590000 399.500000 438.410000 ;
      RECT 307.500000 437.590000 349.500000 438.410000 ;
      RECT 207.500000 437.590000 299.500000 438.410000 ;
      RECT 107.500000 437.590000 199.500000 438.410000 ;
      RECT 57.500000 437.590000 99.500000 438.410000 ;
      RECT 15.500000 437.590000 49.500000 438.410000 ;
      RECT 1183.500000 436.410000 1186.000000 439.590000 ;
      RECT 1166.500000 436.410000 1170.500000 437.590000 ;
      RECT 1157.500000 436.410000 1158.500000 437.590000 ;
      RECT 1116.500000 436.410000 1149.500000 437.590000 ;
      RECT 1107.500000 436.410000 1108.500000 437.590000 ;
      RECT 1066.500000 436.410000 1099.500000 437.590000 ;
      RECT 1057.500000 436.410000 1058.500000 437.590000 ;
      RECT 1016.500000 436.410000 1049.500000 437.590000 ;
      RECT 1007.500000 436.410000 1008.500000 437.590000 ;
      RECT 966.500000 436.410000 999.500000 437.590000 ;
      RECT 957.500000 436.410000 958.500000 437.590000 ;
      RECT 916.500000 436.410000 949.500000 437.590000 ;
      RECT 907.500000 436.410000 908.500000 437.590000 ;
      RECT 866.500000 436.410000 899.500000 437.590000 ;
      RECT 857.500000 436.410000 858.500000 437.590000 ;
      RECT 816.500000 436.410000 849.500000 437.590000 ;
      RECT 807.500000 436.410000 808.500000 437.590000 ;
      RECT 766.500000 436.410000 799.500000 437.590000 ;
      RECT 757.500000 436.410000 758.500000 437.590000 ;
      RECT 736.500000 436.410000 749.500000 439.590000 ;
      RECT 722.500000 436.410000 723.500000 437.590000 ;
      RECT 707.500000 436.410000 708.500000 437.590000 ;
      RECT 666.500000 436.410000 699.500000 437.590000 ;
      RECT 657.500000 436.410000 658.500000 437.590000 ;
      RECT 616.500000 436.410000 649.500000 437.590000 ;
      RECT 607.500000 436.410000 608.500000 437.590000 ;
      RECT 566.500000 436.410000 599.500000 437.590000 ;
      RECT 557.500000 436.410000 558.500000 437.590000 ;
      RECT 516.500000 436.410000 549.500000 437.590000 ;
      RECT 507.500000 436.410000 508.500000 437.590000 ;
      RECT 466.500000 436.410000 499.500000 437.590000 ;
      RECT 457.500000 436.410000 458.500000 437.590000 ;
      RECT 416.500000 436.410000 449.500000 437.590000 ;
      RECT 407.500000 436.410000 408.500000 437.590000 ;
      RECT 366.500000 436.410000 399.500000 437.590000 ;
      RECT 357.500000 436.410000 358.500000 437.590000 ;
      RECT 316.500000 436.410000 349.500000 437.590000 ;
      RECT 307.500000 436.410000 308.500000 437.590000 ;
      RECT 216.500000 436.410000 299.500000 437.590000 ;
      RECT 207.500000 436.410000 208.500000 437.590000 ;
      RECT 116.500000 436.410000 199.500000 437.590000 ;
      RECT 107.500000 436.410000 108.500000 437.590000 ;
      RECT 66.500000 436.410000 99.500000 437.590000 ;
      RECT 57.500000 436.410000 58.500000 437.590000 ;
      RECT 29.500000 436.410000 49.500000 437.590000 ;
      RECT 15.500000 436.410000 16.500000 437.590000 ;
      RECT 0.000000 436.410000 2.500000 439.590000 ;
      RECT 1166.500000 435.590000 1186.000000 436.410000 ;
      RECT 1116.500000 435.590000 1158.500000 436.410000 ;
      RECT 1066.500000 435.590000 1108.500000 436.410000 ;
      RECT 1016.500000 435.590000 1058.500000 436.410000 ;
      RECT 966.500000 435.590000 1008.500000 436.410000 ;
      RECT 916.500000 435.590000 958.500000 436.410000 ;
      RECT 866.500000 435.590000 908.500000 436.410000 ;
      RECT 816.500000 435.590000 858.500000 436.410000 ;
      RECT 766.500000 435.590000 808.500000 436.410000 ;
      RECT 722.500000 435.590000 758.500000 436.410000 ;
      RECT 666.500000 435.590000 708.500000 436.410000 ;
      RECT 616.500000 435.590000 658.500000 436.410000 ;
      RECT 566.500000 435.590000 608.500000 436.410000 ;
      RECT 516.500000 435.590000 558.500000 436.410000 ;
      RECT 466.500000 435.590000 508.500000 436.410000 ;
      RECT 416.500000 435.590000 458.500000 436.410000 ;
      RECT 366.500000 435.590000 408.500000 436.410000 ;
      RECT 316.500000 435.590000 358.500000 436.410000 ;
      RECT 216.500000 435.590000 308.500000 436.410000 ;
      RECT 116.500000 435.590000 208.500000 436.410000 ;
      RECT 66.500000 435.590000 108.500000 436.410000 ;
      RECT 29.500000 435.590000 58.500000 436.410000 ;
      RECT 0.000000 435.590000 16.500000 436.410000 ;
      RECT 1166.500000 434.410000 1170.500000 435.590000 ;
      RECT 1157.500000 434.410000 1158.500000 435.590000 ;
      RECT 1116.500000 434.410000 1149.500000 435.590000 ;
      RECT 1107.500000 434.410000 1108.500000 435.590000 ;
      RECT 1066.500000 434.410000 1099.500000 435.590000 ;
      RECT 1057.500000 434.410000 1058.500000 435.590000 ;
      RECT 1016.500000 434.410000 1049.500000 435.590000 ;
      RECT 1007.500000 434.410000 1008.500000 435.590000 ;
      RECT 966.500000 434.410000 999.500000 435.590000 ;
      RECT 957.500000 434.410000 958.500000 435.590000 ;
      RECT 916.500000 434.410000 949.500000 435.590000 ;
      RECT 907.500000 434.410000 908.500000 435.590000 ;
      RECT 866.500000 434.410000 899.500000 435.590000 ;
      RECT 857.500000 434.410000 858.500000 435.590000 ;
      RECT 816.500000 434.410000 849.500000 435.590000 ;
      RECT 807.500000 434.410000 808.500000 435.590000 ;
      RECT 766.500000 434.410000 799.500000 435.590000 ;
      RECT 757.500000 434.410000 758.500000 435.590000 ;
      RECT 722.500000 434.410000 723.500000 435.590000 ;
      RECT 707.500000 434.410000 708.500000 435.590000 ;
      RECT 666.500000 434.410000 699.500000 435.590000 ;
      RECT 657.500000 434.410000 658.500000 435.590000 ;
      RECT 616.500000 434.410000 649.500000 435.590000 ;
      RECT 607.500000 434.410000 608.500000 435.590000 ;
      RECT 566.500000 434.410000 599.500000 435.590000 ;
      RECT 557.500000 434.410000 558.500000 435.590000 ;
      RECT 516.500000 434.410000 549.500000 435.590000 ;
      RECT 507.500000 434.410000 508.500000 435.590000 ;
      RECT 466.500000 434.410000 499.500000 435.590000 ;
      RECT 457.500000 434.410000 458.500000 435.590000 ;
      RECT 416.500000 434.410000 449.500000 435.590000 ;
      RECT 407.500000 434.410000 408.500000 435.590000 ;
      RECT 366.500000 434.410000 399.500000 435.590000 ;
      RECT 357.500000 434.410000 358.500000 435.590000 ;
      RECT 316.500000 434.410000 349.500000 435.590000 ;
      RECT 307.500000 434.410000 308.500000 435.590000 ;
      RECT 216.500000 434.410000 299.500000 435.590000 ;
      RECT 207.500000 434.410000 208.500000 435.590000 ;
      RECT 116.500000 434.410000 199.500000 435.590000 ;
      RECT 107.500000 434.410000 108.500000 435.590000 ;
      RECT 66.500000 434.410000 99.500000 435.590000 ;
      RECT 57.500000 434.410000 58.500000 435.590000 ;
      RECT 29.500000 434.410000 49.500000 435.590000 ;
      RECT 15.500000 434.410000 16.500000 435.590000 ;
      RECT 1157.500000 433.590000 1170.500000 434.410000 ;
      RECT 1107.500000 433.590000 1149.500000 434.410000 ;
      RECT 1057.500000 433.590000 1099.500000 434.410000 ;
      RECT 1007.500000 433.590000 1049.500000 434.410000 ;
      RECT 957.500000 433.590000 999.500000 434.410000 ;
      RECT 907.500000 433.590000 949.500000 434.410000 ;
      RECT 857.500000 433.590000 899.500000 434.410000 ;
      RECT 807.500000 433.590000 849.500000 434.410000 ;
      RECT 757.500000 433.590000 799.500000 434.410000 ;
      RECT 707.500000 433.590000 723.500000 434.410000 ;
      RECT 657.500000 433.590000 699.500000 434.410000 ;
      RECT 607.500000 433.590000 649.500000 434.410000 ;
      RECT 557.500000 433.590000 599.500000 434.410000 ;
      RECT 507.500000 433.590000 549.500000 434.410000 ;
      RECT 457.500000 433.590000 499.500000 434.410000 ;
      RECT 407.500000 433.590000 449.500000 434.410000 ;
      RECT 357.500000 433.590000 399.500000 434.410000 ;
      RECT 307.500000 433.590000 349.500000 434.410000 ;
      RECT 207.500000 433.590000 299.500000 434.410000 ;
      RECT 107.500000 433.590000 199.500000 434.410000 ;
      RECT 57.500000 433.590000 99.500000 434.410000 ;
      RECT 15.500000 433.590000 49.500000 434.410000 ;
      RECT 1183.500000 432.410000 1186.000000 435.590000 ;
      RECT 1166.500000 432.410000 1170.500000 433.590000 ;
      RECT 1157.500000 432.410000 1158.500000 433.590000 ;
      RECT 1116.500000 432.410000 1149.500000 433.590000 ;
      RECT 1107.500000 432.410000 1108.500000 433.590000 ;
      RECT 1066.500000 432.410000 1099.500000 433.590000 ;
      RECT 1057.500000 432.410000 1058.500000 433.590000 ;
      RECT 1016.500000 432.410000 1049.500000 433.590000 ;
      RECT 1007.500000 432.410000 1008.500000 433.590000 ;
      RECT 966.500000 432.410000 999.500000 433.590000 ;
      RECT 957.500000 432.410000 958.500000 433.590000 ;
      RECT 916.500000 432.410000 949.500000 433.590000 ;
      RECT 907.500000 432.410000 908.500000 433.590000 ;
      RECT 866.500000 432.410000 899.500000 433.590000 ;
      RECT 857.500000 432.410000 858.500000 433.590000 ;
      RECT 816.500000 432.410000 849.500000 433.590000 ;
      RECT 807.500000 432.410000 808.500000 433.590000 ;
      RECT 766.500000 432.410000 799.500000 433.590000 ;
      RECT 757.500000 432.410000 758.500000 433.590000 ;
      RECT 736.500000 432.410000 749.500000 435.590000 ;
      RECT 722.500000 432.410000 723.500000 433.590000 ;
      RECT 707.500000 432.410000 708.500000 433.590000 ;
      RECT 666.500000 432.410000 699.500000 433.590000 ;
      RECT 657.500000 432.410000 658.500000 433.590000 ;
      RECT 616.500000 432.410000 649.500000 433.590000 ;
      RECT 607.500000 432.410000 608.500000 433.590000 ;
      RECT 566.500000 432.410000 599.500000 433.590000 ;
      RECT 557.500000 432.410000 558.500000 433.590000 ;
      RECT 516.500000 432.410000 549.500000 433.590000 ;
      RECT 507.500000 432.410000 508.500000 433.590000 ;
      RECT 466.500000 432.410000 499.500000 433.590000 ;
      RECT 457.500000 432.410000 458.500000 433.590000 ;
      RECT 416.500000 432.410000 449.500000 433.590000 ;
      RECT 407.500000 432.410000 408.500000 433.590000 ;
      RECT 366.500000 432.410000 399.500000 433.590000 ;
      RECT 357.500000 432.410000 358.500000 433.590000 ;
      RECT 316.500000 432.410000 349.500000 433.590000 ;
      RECT 307.500000 432.410000 308.500000 433.590000 ;
      RECT 216.500000 432.410000 299.500000 433.590000 ;
      RECT 207.500000 432.410000 208.500000 433.590000 ;
      RECT 116.500000 432.410000 199.500000 433.590000 ;
      RECT 107.500000 432.410000 108.500000 433.590000 ;
      RECT 66.500000 432.410000 99.500000 433.590000 ;
      RECT 57.500000 432.410000 58.500000 433.590000 ;
      RECT 29.500000 432.410000 49.500000 433.590000 ;
      RECT 15.500000 432.410000 16.500000 433.590000 ;
      RECT 0.000000 432.410000 2.500000 435.590000 ;
      RECT 1166.500000 431.590000 1186.000000 432.410000 ;
      RECT 1116.500000 431.590000 1158.500000 432.410000 ;
      RECT 1066.500000 431.590000 1108.500000 432.410000 ;
      RECT 1016.500000 431.590000 1058.500000 432.410000 ;
      RECT 966.500000 431.590000 1008.500000 432.410000 ;
      RECT 916.500000 431.590000 958.500000 432.410000 ;
      RECT 866.500000 431.590000 908.500000 432.410000 ;
      RECT 816.500000 431.590000 858.500000 432.410000 ;
      RECT 766.500000 431.590000 808.500000 432.410000 ;
      RECT 722.500000 431.590000 758.500000 432.410000 ;
      RECT 666.500000 431.590000 708.500000 432.410000 ;
      RECT 616.500000 431.590000 658.500000 432.410000 ;
      RECT 566.500000 431.590000 608.500000 432.410000 ;
      RECT 516.500000 431.590000 558.500000 432.410000 ;
      RECT 466.500000 431.590000 508.500000 432.410000 ;
      RECT 416.500000 431.590000 458.500000 432.410000 ;
      RECT 366.500000 431.590000 408.500000 432.410000 ;
      RECT 316.500000 431.590000 358.500000 432.410000 ;
      RECT 216.500000 431.590000 308.500000 432.410000 ;
      RECT 116.500000 431.590000 208.500000 432.410000 ;
      RECT 66.500000 431.590000 108.500000 432.410000 ;
      RECT 29.500000 431.590000 58.500000 432.410000 ;
      RECT 0.000000 431.590000 16.500000 432.410000 ;
      RECT 1166.500000 430.410000 1170.500000 431.590000 ;
      RECT 1157.500000 430.410000 1158.500000 431.590000 ;
      RECT 1116.500000 430.410000 1149.500000 431.590000 ;
      RECT 1107.500000 430.410000 1108.500000 431.590000 ;
      RECT 1066.500000 430.410000 1099.500000 431.590000 ;
      RECT 1057.500000 430.410000 1058.500000 431.590000 ;
      RECT 1016.500000 430.410000 1049.500000 431.590000 ;
      RECT 1007.500000 430.410000 1008.500000 431.590000 ;
      RECT 966.500000 430.410000 999.500000 431.590000 ;
      RECT 957.500000 430.410000 958.500000 431.590000 ;
      RECT 916.500000 430.410000 949.500000 431.590000 ;
      RECT 907.500000 430.410000 908.500000 431.590000 ;
      RECT 866.500000 430.410000 899.500000 431.590000 ;
      RECT 857.500000 430.410000 858.500000 431.590000 ;
      RECT 816.500000 430.410000 849.500000 431.590000 ;
      RECT 807.500000 430.410000 808.500000 431.590000 ;
      RECT 766.500000 430.410000 799.500000 431.590000 ;
      RECT 757.500000 430.410000 758.500000 431.590000 ;
      RECT 722.500000 430.410000 749.500000 431.590000 ;
      RECT 707.500000 430.410000 708.500000 431.590000 ;
      RECT 666.500000 430.410000 699.500000 431.590000 ;
      RECT 657.500000 430.410000 658.500000 431.590000 ;
      RECT 616.500000 430.410000 649.500000 431.590000 ;
      RECT 607.500000 430.410000 608.500000 431.590000 ;
      RECT 566.500000 430.410000 599.500000 431.590000 ;
      RECT 557.500000 430.410000 558.500000 431.590000 ;
      RECT 516.500000 430.410000 549.500000 431.590000 ;
      RECT 507.500000 430.410000 508.500000 431.590000 ;
      RECT 466.500000 430.410000 499.500000 431.590000 ;
      RECT 457.500000 430.410000 458.500000 431.590000 ;
      RECT 416.500000 430.410000 449.500000 431.590000 ;
      RECT 407.500000 430.410000 408.500000 431.590000 ;
      RECT 366.500000 430.410000 399.500000 431.590000 ;
      RECT 357.500000 430.410000 358.500000 431.590000 ;
      RECT 316.500000 430.410000 349.500000 431.590000 ;
      RECT 307.500000 430.410000 308.500000 431.590000 ;
      RECT 216.500000 430.410000 299.500000 431.590000 ;
      RECT 207.500000 430.410000 208.500000 431.590000 ;
      RECT 116.500000 430.410000 199.500000 431.590000 ;
      RECT 107.500000 430.410000 108.500000 431.590000 ;
      RECT 66.500000 430.410000 99.500000 431.590000 ;
      RECT 57.500000 430.410000 58.500000 431.590000 ;
      RECT 29.500000 430.410000 49.500000 431.590000 ;
      RECT 15.500000 430.410000 16.500000 431.590000 ;
      RECT 1157.500000 429.590000 1170.500000 430.410000 ;
      RECT 1107.500000 429.590000 1149.500000 430.410000 ;
      RECT 1057.500000 429.590000 1099.500000 430.410000 ;
      RECT 1007.500000 429.590000 1049.500000 430.410000 ;
      RECT 957.500000 429.590000 999.500000 430.410000 ;
      RECT 907.500000 429.590000 949.500000 430.410000 ;
      RECT 857.500000 429.590000 899.500000 430.410000 ;
      RECT 807.500000 429.590000 849.500000 430.410000 ;
      RECT 757.500000 429.590000 799.500000 430.410000 ;
      RECT 707.500000 429.590000 749.500000 430.410000 ;
      RECT 657.500000 429.590000 699.500000 430.410000 ;
      RECT 607.500000 429.590000 649.500000 430.410000 ;
      RECT 557.500000 429.590000 599.500000 430.410000 ;
      RECT 507.500000 429.590000 549.500000 430.410000 ;
      RECT 457.500000 429.590000 499.500000 430.410000 ;
      RECT 407.500000 429.590000 449.500000 430.410000 ;
      RECT 357.500000 429.590000 399.500000 430.410000 ;
      RECT 307.500000 429.590000 349.500000 430.410000 ;
      RECT 207.500000 429.590000 299.500000 430.410000 ;
      RECT 107.500000 429.590000 199.500000 430.410000 ;
      RECT 57.500000 429.590000 99.500000 430.410000 ;
      RECT 15.500000 429.590000 49.500000 430.410000 ;
      RECT 1183.500000 428.410000 1186.000000 431.590000 ;
      RECT 1169.500000 428.410000 1170.500000 429.590000 ;
      RECT 1116.500000 428.410000 1149.500000 429.590000 ;
      RECT 1107.500000 428.410000 1108.500000 429.590000 ;
      RECT 1066.500000 428.410000 1099.500000 429.590000 ;
      RECT 1057.500000 428.410000 1058.500000 429.590000 ;
      RECT 1016.500000 428.410000 1049.500000 429.590000 ;
      RECT 1007.500000 428.410000 1008.500000 429.590000 ;
      RECT 966.500000 428.410000 999.500000 429.590000 ;
      RECT 957.500000 428.410000 958.500000 429.590000 ;
      RECT 916.500000 428.410000 949.500000 429.590000 ;
      RECT 907.500000 428.410000 908.500000 429.590000 ;
      RECT 866.500000 428.410000 899.500000 429.590000 ;
      RECT 857.500000 428.410000 858.500000 429.590000 ;
      RECT 816.500000 428.410000 849.500000 429.590000 ;
      RECT 807.500000 428.410000 808.500000 429.590000 ;
      RECT 766.500000 428.410000 799.500000 429.590000 ;
      RECT 757.500000 428.410000 758.500000 429.590000 ;
      RECT 722.500000 428.410000 749.500000 429.590000 ;
      RECT 707.500000 428.410000 709.500000 429.590000 ;
      RECT 666.500000 428.410000 699.500000 429.590000 ;
      RECT 657.500000 428.410000 658.500000 429.590000 ;
      RECT 616.500000 428.410000 649.500000 429.590000 ;
      RECT 607.500000 428.410000 608.500000 429.590000 ;
      RECT 566.500000 428.410000 599.500000 429.590000 ;
      RECT 557.500000 428.410000 558.500000 429.590000 ;
      RECT 516.500000 428.410000 549.500000 429.590000 ;
      RECT 507.500000 428.410000 508.500000 429.590000 ;
      RECT 466.500000 428.410000 499.500000 429.590000 ;
      RECT 457.500000 428.410000 458.500000 429.590000 ;
      RECT 416.500000 428.410000 449.500000 429.590000 ;
      RECT 407.500000 428.410000 408.500000 429.590000 ;
      RECT 366.500000 428.410000 399.500000 429.590000 ;
      RECT 357.500000 428.410000 358.500000 429.590000 ;
      RECT 316.500000 428.410000 349.500000 429.590000 ;
      RECT 307.500000 428.410000 308.500000 429.590000 ;
      RECT 216.500000 428.410000 299.500000 429.590000 ;
      RECT 207.500000 428.410000 208.500000 429.590000 ;
      RECT 116.500000 428.410000 199.500000 429.590000 ;
      RECT 107.500000 428.410000 108.500000 429.590000 ;
      RECT 66.500000 428.410000 99.500000 429.590000 ;
      RECT 57.500000 428.410000 58.500000 429.590000 ;
      RECT 29.500000 428.410000 49.500000 429.590000 ;
      RECT 15.500000 428.410000 16.500000 429.590000 ;
      RECT 0.000000 428.410000 2.500000 431.590000 ;
      RECT 1169.500000 427.590000 1186.000000 428.410000 ;
      RECT 1116.500000 427.590000 1156.500000 428.410000 ;
      RECT 1066.500000 427.590000 1108.500000 428.410000 ;
      RECT 1016.500000 427.590000 1058.500000 428.410000 ;
      RECT 966.500000 427.590000 1008.500000 428.410000 ;
      RECT 916.500000 427.590000 958.500000 428.410000 ;
      RECT 866.500000 427.590000 908.500000 428.410000 ;
      RECT 816.500000 427.590000 858.500000 428.410000 ;
      RECT 766.500000 427.590000 808.500000 428.410000 ;
      RECT 722.500000 427.590000 758.500000 428.410000 ;
      RECT 666.500000 427.590000 709.500000 428.410000 ;
      RECT 616.500000 427.590000 658.500000 428.410000 ;
      RECT 566.500000 427.590000 608.500000 428.410000 ;
      RECT 516.500000 427.590000 558.500000 428.410000 ;
      RECT 466.500000 427.590000 508.500000 428.410000 ;
      RECT 416.500000 427.590000 458.500000 428.410000 ;
      RECT 366.500000 427.590000 408.500000 428.410000 ;
      RECT 316.500000 427.590000 358.500000 428.410000 ;
      RECT 216.500000 427.590000 308.500000 428.410000 ;
      RECT 116.500000 427.590000 208.500000 428.410000 ;
      RECT 66.500000 427.590000 108.500000 428.410000 ;
      RECT 29.500000 427.590000 58.500000 428.410000 ;
      RECT 0.000000 427.590000 16.500000 428.410000 ;
      RECT 1169.500000 426.410000 1170.500000 427.590000 ;
      RECT 1116.500000 426.410000 1149.500000 427.590000 ;
      RECT 1107.500000 426.410000 1108.500000 427.590000 ;
      RECT 1066.500000 426.410000 1099.500000 427.590000 ;
      RECT 1057.500000 426.410000 1058.500000 427.590000 ;
      RECT 1016.500000 426.410000 1049.500000 427.590000 ;
      RECT 1007.500000 426.410000 1008.500000 427.590000 ;
      RECT 966.500000 426.410000 999.500000 427.590000 ;
      RECT 957.500000 426.410000 958.500000 427.590000 ;
      RECT 916.500000 426.410000 949.500000 427.590000 ;
      RECT 907.500000 426.410000 908.500000 427.590000 ;
      RECT 866.500000 426.410000 899.500000 427.590000 ;
      RECT 857.500000 426.410000 858.500000 427.590000 ;
      RECT 816.500000 426.410000 849.500000 427.590000 ;
      RECT 807.500000 426.410000 808.500000 427.590000 ;
      RECT 766.500000 426.410000 799.500000 427.590000 ;
      RECT 757.500000 426.410000 758.500000 427.590000 ;
      RECT 722.500000 426.410000 749.500000 427.590000 ;
      RECT 707.500000 426.410000 709.500000 427.590000 ;
      RECT 666.500000 426.410000 699.500000 427.590000 ;
      RECT 657.500000 426.410000 658.500000 427.590000 ;
      RECT 616.500000 426.410000 649.500000 427.590000 ;
      RECT 607.500000 426.410000 608.500000 427.590000 ;
      RECT 566.500000 426.410000 599.500000 427.590000 ;
      RECT 557.500000 426.410000 558.500000 427.590000 ;
      RECT 516.500000 426.410000 549.500000 427.590000 ;
      RECT 507.500000 426.410000 508.500000 427.590000 ;
      RECT 466.500000 426.410000 499.500000 427.590000 ;
      RECT 457.500000 426.410000 458.500000 427.590000 ;
      RECT 416.500000 426.410000 449.500000 427.590000 ;
      RECT 407.500000 426.410000 408.500000 427.590000 ;
      RECT 366.500000 426.410000 399.500000 427.590000 ;
      RECT 357.500000 426.410000 358.500000 427.590000 ;
      RECT 316.500000 426.410000 349.500000 427.590000 ;
      RECT 307.500000 426.410000 308.500000 427.590000 ;
      RECT 216.500000 426.410000 299.500000 427.590000 ;
      RECT 207.500000 426.410000 208.500000 427.590000 ;
      RECT 116.500000 426.410000 199.500000 427.590000 ;
      RECT 107.500000 426.410000 108.500000 427.590000 ;
      RECT 66.500000 426.410000 99.500000 427.590000 ;
      RECT 57.500000 426.410000 58.500000 427.590000 ;
      RECT 29.500000 426.410000 49.500000 427.590000 ;
      RECT 15.500000 426.410000 16.500000 427.590000 ;
      RECT 1157.500000 425.590000 1170.500000 426.410000 ;
      RECT 1107.500000 425.590000 1149.500000 426.410000 ;
      RECT 1057.500000 425.590000 1099.500000 426.410000 ;
      RECT 1007.500000 425.590000 1049.500000 426.410000 ;
      RECT 957.500000 425.590000 999.500000 426.410000 ;
      RECT 907.500000 425.590000 949.500000 426.410000 ;
      RECT 857.500000 425.590000 899.500000 426.410000 ;
      RECT 807.500000 425.590000 849.500000 426.410000 ;
      RECT 757.500000 425.590000 799.500000 426.410000 ;
      RECT 707.500000 425.590000 749.500000 426.410000 ;
      RECT 657.500000 425.590000 699.500000 426.410000 ;
      RECT 607.500000 425.590000 649.500000 426.410000 ;
      RECT 557.500000 425.590000 599.500000 426.410000 ;
      RECT 507.500000 425.590000 549.500000 426.410000 ;
      RECT 457.500000 425.590000 499.500000 426.410000 ;
      RECT 407.500000 425.590000 449.500000 426.410000 ;
      RECT 357.500000 425.590000 399.500000 426.410000 ;
      RECT 307.500000 425.590000 349.500000 426.410000 ;
      RECT 207.500000 425.590000 299.500000 426.410000 ;
      RECT 107.500000 425.590000 199.500000 426.410000 ;
      RECT 57.500000 425.590000 99.500000 426.410000 ;
      RECT 15.500000 425.590000 49.500000 426.410000 ;
      RECT 1183.500000 424.410000 1186.000000 427.590000 ;
      RECT 1169.500000 424.410000 1170.500000 425.590000 ;
      RECT 1116.500000 424.410000 1149.500000 425.590000 ;
      RECT 1107.500000 424.410000 1108.500000 425.590000 ;
      RECT 1066.500000 424.410000 1099.500000 425.590000 ;
      RECT 1057.500000 424.410000 1058.500000 425.590000 ;
      RECT 1016.500000 424.410000 1049.500000 425.590000 ;
      RECT 1007.500000 424.410000 1008.500000 425.590000 ;
      RECT 966.500000 424.410000 999.500000 425.590000 ;
      RECT 957.500000 424.410000 958.500000 425.590000 ;
      RECT 916.500000 424.410000 949.500000 425.590000 ;
      RECT 907.500000 424.410000 908.500000 425.590000 ;
      RECT 866.500000 424.410000 899.500000 425.590000 ;
      RECT 857.500000 424.410000 858.500000 425.590000 ;
      RECT 816.500000 424.410000 849.500000 425.590000 ;
      RECT 807.500000 424.410000 808.500000 425.590000 ;
      RECT 766.500000 424.410000 799.500000 425.590000 ;
      RECT 757.500000 424.410000 758.500000 425.590000 ;
      RECT 722.500000 424.410000 749.500000 425.590000 ;
      RECT 707.500000 424.410000 709.500000 425.590000 ;
      RECT 666.500000 424.410000 699.500000 425.590000 ;
      RECT 657.500000 424.410000 658.500000 425.590000 ;
      RECT 616.500000 424.410000 649.500000 425.590000 ;
      RECT 607.500000 424.410000 608.500000 425.590000 ;
      RECT 566.500000 424.410000 599.500000 425.590000 ;
      RECT 557.500000 424.410000 558.500000 425.590000 ;
      RECT 516.500000 424.410000 549.500000 425.590000 ;
      RECT 507.500000 424.410000 508.500000 425.590000 ;
      RECT 466.500000 424.410000 499.500000 425.590000 ;
      RECT 457.500000 424.410000 458.500000 425.590000 ;
      RECT 416.500000 424.410000 449.500000 425.590000 ;
      RECT 407.500000 424.410000 408.500000 425.590000 ;
      RECT 366.500000 424.410000 399.500000 425.590000 ;
      RECT 357.500000 424.410000 358.500000 425.590000 ;
      RECT 316.500000 424.410000 349.500000 425.590000 ;
      RECT 307.500000 424.410000 308.500000 425.590000 ;
      RECT 216.500000 424.410000 299.500000 425.590000 ;
      RECT 207.500000 424.410000 208.500000 425.590000 ;
      RECT 116.500000 424.410000 199.500000 425.590000 ;
      RECT 107.500000 424.410000 108.500000 425.590000 ;
      RECT 66.500000 424.410000 99.500000 425.590000 ;
      RECT 57.500000 424.410000 58.500000 425.590000 ;
      RECT 29.500000 424.410000 49.500000 425.590000 ;
      RECT 15.500000 424.410000 16.500000 425.590000 ;
      RECT 0.000000 424.410000 2.500000 427.590000 ;
      RECT 1169.500000 423.590000 1186.000000 424.410000 ;
      RECT 1116.500000 423.590000 1156.500000 424.410000 ;
      RECT 1066.500000 423.590000 1108.500000 424.410000 ;
      RECT 1016.500000 423.590000 1058.500000 424.410000 ;
      RECT 966.500000 423.590000 1008.500000 424.410000 ;
      RECT 916.500000 423.590000 958.500000 424.410000 ;
      RECT 866.500000 423.590000 908.500000 424.410000 ;
      RECT 816.500000 423.590000 858.500000 424.410000 ;
      RECT 766.500000 423.590000 808.500000 424.410000 ;
      RECT 722.500000 423.590000 758.500000 424.410000 ;
      RECT 666.500000 423.590000 709.500000 424.410000 ;
      RECT 616.500000 423.590000 658.500000 424.410000 ;
      RECT 566.500000 423.590000 608.500000 424.410000 ;
      RECT 516.500000 423.590000 558.500000 424.410000 ;
      RECT 466.500000 423.590000 508.500000 424.410000 ;
      RECT 416.500000 423.590000 458.500000 424.410000 ;
      RECT 366.500000 423.590000 408.500000 424.410000 ;
      RECT 316.500000 423.590000 358.500000 424.410000 ;
      RECT 216.500000 423.590000 308.500000 424.410000 ;
      RECT 116.500000 423.590000 208.500000 424.410000 ;
      RECT 66.500000 423.590000 108.500000 424.410000 ;
      RECT 29.500000 423.590000 58.500000 424.410000 ;
      RECT 0.000000 423.590000 16.500000 424.410000 ;
      RECT 1169.500000 422.410000 1170.500000 423.590000 ;
      RECT 1116.500000 422.410000 1149.500000 423.590000 ;
      RECT 1107.500000 422.410000 1108.500000 423.590000 ;
      RECT 1066.500000 422.410000 1099.500000 423.590000 ;
      RECT 1057.500000 422.410000 1058.500000 423.590000 ;
      RECT 1016.500000 422.410000 1049.500000 423.590000 ;
      RECT 1007.500000 422.410000 1008.500000 423.590000 ;
      RECT 966.500000 422.410000 999.500000 423.590000 ;
      RECT 957.500000 422.410000 958.500000 423.590000 ;
      RECT 916.500000 422.410000 949.500000 423.590000 ;
      RECT 907.500000 422.410000 908.500000 423.590000 ;
      RECT 866.500000 422.410000 899.500000 423.590000 ;
      RECT 857.500000 422.410000 858.500000 423.590000 ;
      RECT 816.500000 422.410000 849.500000 423.590000 ;
      RECT 807.500000 422.410000 808.500000 423.590000 ;
      RECT 766.500000 422.410000 799.500000 423.590000 ;
      RECT 757.500000 422.410000 758.500000 423.590000 ;
      RECT 722.500000 422.410000 749.500000 423.590000 ;
      RECT 707.500000 422.410000 709.500000 423.590000 ;
      RECT 666.500000 422.410000 699.500000 423.590000 ;
      RECT 657.500000 422.410000 658.500000 423.590000 ;
      RECT 616.500000 422.410000 649.500000 423.590000 ;
      RECT 607.500000 422.410000 608.500000 423.590000 ;
      RECT 566.500000 422.410000 599.500000 423.590000 ;
      RECT 557.500000 422.410000 558.500000 423.590000 ;
      RECT 516.500000 422.410000 549.500000 423.590000 ;
      RECT 507.500000 422.410000 508.500000 423.590000 ;
      RECT 466.500000 422.410000 499.500000 423.590000 ;
      RECT 457.500000 422.410000 458.500000 423.590000 ;
      RECT 416.500000 422.410000 449.500000 423.590000 ;
      RECT 407.500000 422.410000 408.500000 423.590000 ;
      RECT 366.500000 422.410000 399.500000 423.590000 ;
      RECT 357.500000 422.410000 358.500000 423.590000 ;
      RECT 316.500000 422.410000 349.500000 423.590000 ;
      RECT 307.500000 422.410000 308.500000 423.590000 ;
      RECT 216.500000 422.410000 299.500000 423.590000 ;
      RECT 207.500000 422.410000 208.500000 423.590000 ;
      RECT 116.500000 422.410000 199.500000 423.590000 ;
      RECT 107.500000 422.410000 108.500000 423.590000 ;
      RECT 66.500000 422.410000 99.500000 423.590000 ;
      RECT 57.500000 422.410000 58.500000 423.590000 ;
      RECT 29.500000 422.410000 49.500000 423.590000 ;
      RECT 15.500000 422.410000 16.500000 423.590000 ;
      RECT 1157.500000 421.590000 1170.500000 422.410000 ;
      RECT 1107.500000 421.590000 1149.500000 422.410000 ;
      RECT 1057.500000 421.590000 1099.500000 422.410000 ;
      RECT 1007.500000 421.590000 1049.500000 422.410000 ;
      RECT 957.500000 421.590000 999.500000 422.410000 ;
      RECT 907.500000 421.590000 949.500000 422.410000 ;
      RECT 857.500000 421.590000 899.500000 422.410000 ;
      RECT 807.500000 421.590000 849.500000 422.410000 ;
      RECT 757.500000 421.590000 799.500000 422.410000 ;
      RECT 707.500000 421.590000 749.500000 422.410000 ;
      RECT 657.500000 421.590000 699.500000 422.410000 ;
      RECT 607.500000 421.590000 649.500000 422.410000 ;
      RECT 557.500000 421.590000 599.500000 422.410000 ;
      RECT 507.500000 421.590000 549.500000 422.410000 ;
      RECT 457.500000 421.590000 499.500000 422.410000 ;
      RECT 407.500000 421.590000 449.500000 422.410000 ;
      RECT 357.500000 421.590000 399.500000 422.410000 ;
      RECT 307.500000 421.590000 349.500000 422.410000 ;
      RECT 207.500000 421.590000 299.500000 422.410000 ;
      RECT 107.500000 421.590000 199.500000 422.410000 ;
      RECT 57.500000 421.590000 99.500000 422.410000 ;
      RECT 15.500000 421.590000 49.500000 422.410000 ;
      RECT 1183.500000 420.410000 1186.000000 423.590000 ;
      RECT 1169.500000 420.410000 1170.500000 421.590000 ;
      RECT 1116.500000 420.410000 1149.500000 421.590000 ;
      RECT 1107.500000 420.410000 1108.500000 421.590000 ;
      RECT 1066.500000 420.410000 1099.500000 421.590000 ;
      RECT 1057.500000 420.410000 1058.500000 421.590000 ;
      RECT 1016.500000 420.410000 1049.500000 421.590000 ;
      RECT 1007.500000 420.410000 1008.500000 421.590000 ;
      RECT 966.500000 420.410000 999.500000 421.590000 ;
      RECT 957.500000 420.410000 958.500000 421.590000 ;
      RECT 916.500000 420.410000 949.500000 421.590000 ;
      RECT 907.500000 420.410000 908.500000 421.590000 ;
      RECT 866.500000 420.410000 899.500000 421.590000 ;
      RECT 857.500000 420.410000 858.500000 421.590000 ;
      RECT 816.500000 420.410000 849.500000 421.590000 ;
      RECT 807.500000 420.410000 808.500000 421.590000 ;
      RECT 766.500000 420.410000 799.500000 421.590000 ;
      RECT 757.500000 420.410000 758.500000 421.590000 ;
      RECT 722.500000 420.410000 749.500000 421.590000 ;
      RECT 707.500000 420.410000 709.500000 421.590000 ;
      RECT 666.500000 420.410000 699.500000 421.590000 ;
      RECT 657.500000 420.410000 658.500000 421.590000 ;
      RECT 616.500000 420.410000 649.500000 421.590000 ;
      RECT 607.500000 420.410000 608.500000 421.590000 ;
      RECT 566.500000 420.410000 599.500000 421.590000 ;
      RECT 557.500000 420.410000 558.500000 421.590000 ;
      RECT 516.500000 420.410000 549.500000 421.590000 ;
      RECT 507.500000 420.410000 508.500000 421.590000 ;
      RECT 466.500000 420.410000 499.500000 421.590000 ;
      RECT 457.500000 420.410000 458.500000 421.590000 ;
      RECT 416.500000 420.410000 449.500000 421.590000 ;
      RECT 407.500000 420.410000 408.500000 421.590000 ;
      RECT 366.500000 420.410000 399.500000 421.590000 ;
      RECT 357.500000 420.410000 358.500000 421.590000 ;
      RECT 316.500000 420.410000 349.500000 421.590000 ;
      RECT 307.500000 420.410000 308.500000 421.590000 ;
      RECT 216.500000 420.410000 299.500000 421.590000 ;
      RECT 207.500000 420.410000 208.500000 421.590000 ;
      RECT 116.500000 420.410000 199.500000 421.590000 ;
      RECT 107.500000 420.410000 108.500000 421.590000 ;
      RECT 66.500000 420.410000 99.500000 421.590000 ;
      RECT 57.500000 420.410000 58.500000 421.590000 ;
      RECT 29.500000 420.410000 49.500000 421.590000 ;
      RECT 15.500000 420.410000 16.500000 421.590000 ;
      RECT 0.000000 420.410000 2.500000 423.590000 ;
      RECT 1169.500000 419.590000 1186.000000 420.410000 ;
      RECT 1116.500000 419.590000 1156.500000 420.410000 ;
      RECT 1066.500000 419.590000 1108.500000 420.410000 ;
      RECT 1016.500000 419.590000 1058.500000 420.410000 ;
      RECT 966.500000 419.590000 1008.500000 420.410000 ;
      RECT 916.500000 419.590000 958.500000 420.410000 ;
      RECT 866.500000 419.590000 908.500000 420.410000 ;
      RECT 816.500000 419.590000 858.500000 420.410000 ;
      RECT 766.500000 419.590000 808.500000 420.410000 ;
      RECT 722.500000 419.590000 758.500000 420.410000 ;
      RECT 666.500000 419.590000 709.500000 420.410000 ;
      RECT 616.500000 419.590000 658.500000 420.410000 ;
      RECT 566.500000 419.590000 608.500000 420.410000 ;
      RECT 516.500000 419.590000 558.500000 420.410000 ;
      RECT 466.500000 419.590000 508.500000 420.410000 ;
      RECT 366.500000 419.590000 408.500000 420.410000 ;
      RECT 316.500000 419.590000 358.500000 420.410000 ;
      RECT 216.500000 419.590000 308.500000 420.410000 ;
      RECT 116.500000 419.590000 208.500000 420.410000 ;
      RECT 66.500000 419.590000 108.500000 420.410000 ;
      RECT 29.500000 419.590000 58.500000 420.410000 ;
      RECT 0.000000 419.590000 16.500000 420.410000 ;
      RECT 1169.500000 418.410000 1170.500000 419.590000 ;
      RECT 1116.500000 418.410000 1149.500000 419.590000 ;
      RECT 1107.500000 418.410000 1108.500000 419.590000 ;
      RECT 1066.500000 418.410000 1099.500000 419.590000 ;
      RECT 1057.500000 418.410000 1058.500000 419.590000 ;
      RECT 1016.500000 418.410000 1049.500000 419.590000 ;
      RECT 1007.500000 418.410000 1008.500000 419.590000 ;
      RECT 966.500000 418.410000 999.500000 419.590000 ;
      RECT 957.500000 418.410000 958.500000 419.590000 ;
      RECT 916.500000 418.410000 949.500000 419.590000 ;
      RECT 907.500000 418.410000 908.500000 419.590000 ;
      RECT 866.500000 418.410000 899.500000 419.590000 ;
      RECT 857.500000 418.410000 858.500000 419.590000 ;
      RECT 816.500000 418.410000 849.500000 419.590000 ;
      RECT 807.500000 418.410000 808.500000 419.590000 ;
      RECT 766.500000 418.410000 799.500000 419.590000 ;
      RECT 757.500000 418.410000 758.500000 419.590000 ;
      RECT 722.500000 418.410000 749.500000 419.590000 ;
      RECT 707.500000 418.410000 709.500000 419.590000 ;
      RECT 666.500000 418.410000 699.500000 419.590000 ;
      RECT 657.500000 418.410000 658.500000 419.590000 ;
      RECT 616.500000 418.410000 649.500000 419.590000 ;
      RECT 607.500000 418.410000 608.500000 419.590000 ;
      RECT 566.500000 418.410000 599.500000 419.590000 ;
      RECT 557.500000 418.410000 558.500000 419.590000 ;
      RECT 516.500000 418.410000 549.500000 419.590000 ;
      RECT 507.500000 418.410000 508.500000 419.590000 ;
      RECT 466.500000 418.410000 499.500000 419.590000 ;
      RECT 416.500000 418.410000 458.500000 420.410000 ;
      RECT 407.500000 418.410000 408.500000 419.590000 ;
      RECT 366.500000 418.410000 399.500000 419.590000 ;
      RECT 357.500000 418.410000 358.500000 419.590000 ;
      RECT 316.500000 418.410000 349.500000 419.590000 ;
      RECT 307.500000 418.410000 308.500000 419.590000 ;
      RECT 216.500000 418.410000 299.500000 419.590000 ;
      RECT 207.500000 418.410000 208.500000 419.590000 ;
      RECT 116.500000 418.410000 199.500000 419.590000 ;
      RECT 107.500000 418.410000 108.500000 419.590000 ;
      RECT 66.500000 418.410000 99.500000 419.590000 ;
      RECT 57.500000 418.410000 58.500000 419.590000 ;
      RECT 29.500000 418.410000 49.500000 419.590000 ;
      RECT 15.500000 418.410000 16.500000 419.590000 ;
      RECT 1157.500000 417.590000 1170.500000 418.410000 ;
      RECT 1107.500000 417.590000 1149.500000 418.410000 ;
      RECT 1057.500000 417.590000 1099.500000 418.410000 ;
      RECT 1007.500000 417.590000 1049.500000 418.410000 ;
      RECT 957.500000 417.590000 999.500000 418.410000 ;
      RECT 907.500000 417.590000 949.500000 418.410000 ;
      RECT 857.500000 417.590000 899.500000 418.410000 ;
      RECT 807.500000 417.590000 849.500000 418.410000 ;
      RECT 757.500000 417.590000 799.500000 418.410000 ;
      RECT 707.500000 417.590000 749.500000 418.410000 ;
      RECT 657.500000 417.590000 699.500000 418.410000 ;
      RECT 607.500000 417.590000 649.500000 418.410000 ;
      RECT 557.500000 417.590000 599.500000 418.410000 ;
      RECT 507.500000 417.590000 549.500000 418.410000 ;
      RECT 407.500000 417.590000 499.500000 418.410000 ;
      RECT 357.500000 417.590000 399.500000 418.410000 ;
      RECT 307.500000 417.590000 349.500000 418.410000 ;
      RECT 207.500000 417.590000 299.500000 418.410000 ;
      RECT 107.500000 417.590000 199.500000 418.410000 ;
      RECT 57.500000 417.590000 99.500000 418.410000 ;
      RECT 15.500000 417.590000 49.500000 418.410000 ;
      RECT 1183.500000 416.410000 1186.000000 419.590000 ;
      RECT 1169.500000 416.410000 1170.500000 417.590000 ;
      RECT 1116.500000 416.410000 1149.500000 417.590000 ;
      RECT 1107.500000 416.410000 1108.500000 417.590000 ;
      RECT 1066.500000 416.410000 1099.500000 417.590000 ;
      RECT 1057.500000 416.410000 1058.500000 417.590000 ;
      RECT 1016.500000 416.410000 1049.500000 417.590000 ;
      RECT 1007.500000 416.410000 1008.500000 417.590000 ;
      RECT 966.500000 416.410000 999.500000 417.590000 ;
      RECT 957.500000 416.410000 958.500000 417.590000 ;
      RECT 916.500000 416.410000 949.500000 417.590000 ;
      RECT 907.500000 416.410000 908.500000 417.590000 ;
      RECT 866.500000 416.410000 899.500000 417.590000 ;
      RECT 857.500000 416.410000 858.500000 417.590000 ;
      RECT 816.500000 416.410000 849.500000 417.590000 ;
      RECT 807.500000 416.410000 808.500000 417.590000 ;
      RECT 766.500000 416.410000 799.500000 417.590000 ;
      RECT 757.500000 416.410000 758.500000 417.590000 ;
      RECT 720.000000 416.410000 749.500000 417.590000 ;
      RECT 707.500000 416.410000 712.000000 417.590000 ;
      RECT 666.500000 416.410000 699.500000 417.590000 ;
      RECT 657.500000 416.410000 658.500000 417.590000 ;
      RECT 616.500000 416.410000 649.500000 417.590000 ;
      RECT 607.500000 416.410000 608.500000 417.590000 ;
      RECT 566.500000 416.410000 599.500000 417.590000 ;
      RECT 557.500000 416.410000 558.500000 417.590000 ;
      RECT 516.500000 416.410000 549.500000 417.590000 ;
      RECT 507.500000 416.410000 508.500000 417.590000 ;
      RECT 416.500000 416.410000 499.500000 417.590000 ;
      RECT 407.500000 416.410000 408.500000 417.590000 ;
      RECT 366.500000 416.410000 399.500000 417.590000 ;
      RECT 357.500000 416.410000 358.500000 417.590000 ;
      RECT 316.500000 416.410000 349.500000 417.590000 ;
      RECT 307.500000 416.410000 308.500000 417.590000 ;
      RECT 216.500000 416.410000 299.500000 417.590000 ;
      RECT 207.500000 416.410000 208.500000 417.590000 ;
      RECT 116.500000 416.410000 199.500000 417.590000 ;
      RECT 107.500000 416.410000 108.500000 417.590000 ;
      RECT 66.500000 416.410000 99.500000 417.590000 ;
      RECT 57.500000 416.410000 58.500000 417.590000 ;
      RECT 29.500000 416.410000 49.500000 417.590000 ;
      RECT 15.500000 416.410000 16.500000 417.590000 ;
      RECT 0.000000 416.410000 2.500000 419.590000 ;
      RECT 1169.500000 415.590000 1186.000000 416.410000 ;
      RECT 1116.500000 415.590000 1156.500000 416.410000 ;
      RECT 1066.500000 415.590000 1108.500000 416.410000 ;
      RECT 1016.500000 415.590000 1058.500000 416.410000 ;
      RECT 966.500000 415.590000 1008.500000 416.410000 ;
      RECT 916.500000 415.590000 958.500000 416.410000 ;
      RECT 866.500000 415.590000 908.500000 416.410000 ;
      RECT 816.500000 415.590000 858.500000 416.410000 ;
      RECT 766.500000 415.590000 808.500000 416.410000 ;
      RECT 720.000000 415.590000 758.500000 416.410000 ;
      RECT 666.500000 415.590000 712.000000 416.410000 ;
      RECT 616.500000 415.590000 658.500000 416.410000 ;
      RECT 566.500000 415.590000 608.500000 416.410000 ;
      RECT 516.500000 415.590000 558.500000 416.410000 ;
      RECT 416.500000 415.590000 508.500000 416.410000 ;
      RECT 366.500000 415.590000 408.500000 416.410000 ;
      RECT 316.500000 415.590000 358.500000 416.410000 ;
      RECT 216.500000 415.590000 308.500000 416.410000 ;
      RECT 116.500000 415.590000 208.500000 416.410000 ;
      RECT 66.500000 415.590000 108.500000 416.410000 ;
      RECT 29.500000 415.590000 58.500000 416.410000 ;
      RECT 0.000000 415.590000 16.500000 416.410000 ;
      RECT 1169.500000 414.410000 1170.500000 415.590000 ;
      RECT 1116.500000 414.410000 1149.500000 415.590000 ;
      RECT 1107.500000 414.410000 1108.500000 415.590000 ;
      RECT 1066.500000 414.410000 1099.500000 415.590000 ;
      RECT 1057.500000 414.410000 1058.500000 415.590000 ;
      RECT 1016.500000 414.410000 1049.500000 415.590000 ;
      RECT 1007.500000 414.410000 1008.500000 415.590000 ;
      RECT 966.500000 414.410000 999.500000 415.590000 ;
      RECT 957.500000 414.410000 958.500000 415.590000 ;
      RECT 916.500000 414.410000 949.500000 415.590000 ;
      RECT 907.500000 414.410000 908.500000 415.590000 ;
      RECT 866.500000 414.410000 899.500000 415.590000 ;
      RECT 857.500000 414.410000 858.500000 415.590000 ;
      RECT 816.500000 414.410000 849.500000 415.590000 ;
      RECT 807.500000 414.410000 808.500000 415.590000 ;
      RECT 766.500000 414.410000 799.500000 415.590000 ;
      RECT 757.500000 414.410000 758.500000 415.590000 ;
      RECT 720.000000 414.410000 749.500000 415.590000 ;
      RECT 707.500000 414.410000 712.000000 415.590000 ;
      RECT 666.500000 414.410000 699.500000 415.590000 ;
      RECT 657.500000 414.410000 658.500000 415.590000 ;
      RECT 616.500000 414.410000 649.500000 415.590000 ;
      RECT 607.500000 414.410000 608.500000 415.590000 ;
      RECT 566.500000 414.410000 599.500000 415.590000 ;
      RECT 557.500000 414.410000 558.500000 415.590000 ;
      RECT 516.500000 414.410000 549.500000 415.590000 ;
      RECT 507.500000 414.410000 508.500000 415.590000 ;
      RECT 416.500000 414.410000 499.500000 415.590000 ;
      RECT 407.500000 414.410000 408.500000 415.590000 ;
      RECT 366.500000 414.410000 399.500000 415.590000 ;
      RECT 357.500000 414.410000 358.500000 415.590000 ;
      RECT 316.500000 414.410000 349.500000 415.590000 ;
      RECT 307.500000 414.410000 308.500000 415.590000 ;
      RECT 216.500000 414.410000 299.500000 415.590000 ;
      RECT 207.500000 414.410000 208.500000 415.590000 ;
      RECT 116.500000 414.410000 199.500000 415.590000 ;
      RECT 107.500000 414.410000 108.500000 415.590000 ;
      RECT 66.500000 414.410000 99.500000 415.590000 ;
      RECT 57.500000 414.410000 58.500000 415.590000 ;
      RECT 29.500000 414.410000 49.500000 415.590000 ;
      RECT 15.500000 414.410000 16.500000 415.590000 ;
      RECT 1157.500000 413.590000 1170.500000 414.410000 ;
      RECT 1107.500000 413.590000 1149.500000 414.410000 ;
      RECT 1057.500000 413.590000 1099.500000 414.410000 ;
      RECT 1007.500000 413.590000 1049.500000 414.410000 ;
      RECT 957.500000 413.590000 999.500000 414.410000 ;
      RECT 907.500000 413.590000 949.500000 414.410000 ;
      RECT 857.500000 413.590000 899.500000 414.410000 ;
      RECT 807.500000 413.590000 849.500000 414.410000 ;
      RECT 757.500000 413.590000 799.500000 414.410000 ;
      RECT 707.500000 413.590000 749.500000 414.410000 ;
      RECT 657.500000 413.590000 699.500000 414.410000 ;
      RECT 607.500000 413.590000 649.500000 414.410000 ;
      RECT 557.500000 413.590000 599.500000 414.410000 ;
      RECT 507.500000 413.590000 549.500000 414.410000 ;
      RECT 407.500000 413.590000 499.500000 414.410000 ;
      RECT 357.500000 413.590000 399.500000 414.410000 ;
      RECT 307.500000 413.590000 349.500000 414.410000 ;
      RECT 207.500000 413.590000 299.500000 414.410000 ;
      RECT 107.500000 413.590000 199.500000 414.410000 ;
      RECT 57.500000 413.590000 99.500000 414.410000 ;
      RECT 15.500000 413.590000 49.500000 414.410000 ;
      RECT 1183.500000 412.410000 1186.000000 415.590000 ;
      RECT 1169.500000 412.410000 1170.500000 413.590000 ;
      RECT 1116.500000 412.410000 1149.500000 413.590000 ;
      RECT 1107.500000 412.410000 1108.500000 413.590000 ;
      RECT 1066.500000 412.410000 1099.500000 413.590000 ;
      RECT 1057.500000 412.410000 1058.500000 413.590000 ;
      RECT 1016.500000 412.410000 1049.500000 413.590000 ;
      RECT 1007.500000 412.410000 1008.500000 413.590000 ;
      RECT 966.500000 412.410000 999.500000 413.590000 ;
      RECT 957.500000 412.410000 958.500000 413.590000 ;
      RECT 916.500000 412.410000 949.500000 413.590000 ;
      RECT 907.500000 412.410000 908.500000 413.590000 ;
      RECT 866.500000 412.410000 899.500000 413.590000 ;
      RECT 857.500000 412.410000 858.500000 413.590000 ;
      RECT 816.500000 412.410000 849.500000 413.590000 ;
      RECT 807.500000 412.410000 808.500000 413.590000 ;
      RECT 766.500000 412.410000 799.500000 413.590000 ;
      RECT 757.500000 412.410000 758.500000 413.590000 ;
      RECT 720.000000 412.410000 749.500000 413.590000 ;
      RECT 707.500000 412.410000 708.500000 413.590000 ;
      RECT 666.500000 412.410000 699.500000 413.590000 ;
      RECT 657.500000 412.410000 658.500000 413.590000 ;
      RECT 616.500000 412.410000 649.500000 413.590000 ;
      RECT 607.500000 412.410000 608.500000 413.590000 ;
      RECT 566.500000 412.410000 599.500000 413.590000 ;
      RECT 557.500000 412.410000 558.500000 413.590000 ;
      RECT 516.500000 412.410000 549.500000 413.590000 ;
      RECT 507.500000 412.410000 508.500000 413.590000 ;
      RECT 416.500000 412.410000 499.500000 413.590000 ;
      RECT 407.500000 412.410000 408.500000 413.590000 ;
      RECT 366.500000 412.410000 399.500000 413.590000 ;
      RECT 357.500000 412.410000 358.500000 413.590000 ;
      RECT 316.500000 412.410000 349.500000 413.590000 ;
      RECT 307.500000 412.410000 308.500000 413.590000 ;
      RECT 216.500000 412.410000 299.500000 413.590000 ;
      RECT 207.500000 412.410000 208.500000 413.590000 ;
      RECT 116.500000 412.410000 199.500000 413.590000 ;
      RECT 107.500000 412.410000 108.500000 413.590000 ;
      RECT 66.500000 412.410000 99.500000 413.590000 ;
      RECT 57.500000 412.410000 58.500000 413.590000 ;
      RECT 29.500000 412.410000 49.500000 413.590000 ;
      RECT 15.500000 412.410000 16.500000 413.590000 ;
      RECT 0.000000 412.410000 2.500000 415.590000 ;
      RECT 1169.500000 411.590000 1186.000000 412.410000 ;
      RECT 1116.500000 411.590000 1156.500000 412.410000 ;
      RECT 1066.500000 411.590000 1108.500000 412.410000 ;
      RECT 1016.500000 411.590000 1058.500000 412.410000 ;
      RECT 966.500000 411.590000 1008.500000 412.410000 ;
      RECT 916.500000 411.590000 958.500000 412.410000 ;
      RECT 866.500000 411.590000 908.500000 412.410000 ;
      RECT 816.500000 411.590000 858.500000 412.410000 ;
      RECT 766.500000 411.590000 808.500000 412.410000 ;
      RECT 720.000000 411.590000 758.500000 412.410000 ;
      RECT 666.500000 411.590000 708.500000 412.410000 ;
      RECT 616.500000 411.590000 658.500000 412.410000 ;
      RECT 566.500000 411.590000 608.500000 412.410000 ;
      RECT 516.500000 411.590000 558.500000 412.410000 ;
      RECT 416.500000 411.590000 508.500000 412.410000 ;
      RECT 366.500000 411.590000 408.500000 412.410000 ;
      RECT 316.500000 411.590000 358.500000 412.410000 ;
      RECT 216.500000 411.590000 308.500000 412.410000 ;
      RECT 116.500000 411.590000 208.500000 412.410000 ;
      RECT 66.500000 411.590000 108.500000 412.410000 ;
      RECT 29.500000 411.590000 58.500000 412.410000 ;
      RECT 0.000000 411.590000 16.500000 412.410000 ;
      RECT 1169.500000 410.410000 1170.500000 411.590000 ;
      RECT 1116.500000 410.410000 1149.500000 411.590000 ;
      RECT 1107.500000 410.410000 1108.500000 411.590000 ;
      RECT 1066.500000 410.410000 1099.500000 411.590000 ;
      RECT 1057.500000 410.410000 1058.500000 411.590000 ;
      RECT 1016.500000 410.410000 1049.500000 411.590000 ;
      RECT 1007.500000 410.410000 1008.500000 411.590000 ;
      RECT 966.500000 410.410000 999.500000 411.590000 ;
      RECT 957.500000 410.410000 958.500000 411.590000 ;
      RECT 916.500000 410.410000 949.500000 411.590000 ;
      RECT 907.500000 410.410000 908.500000 411.590000 ;
      RECT 866.500000 410.410000 899.500000 411.590000 ;
      RECT 857.500000 410.410000 858.500000 411.590000 ;
      RECT 816.500000 410.410000 849.500000 411.590000 ;
      RECT 807.500000 410.410000 808.500000 411.590000 ;
      RECT 766.500000 410.410000 799.500000 411.590000 ;
      RECT 757.500000 410.410000 758.500000 411.590000 ;
      RECT 720.000000 410.410000 749.500000 411.590000 ;
      RECT 707.500000 410.410000 708.500000 411.590000 ;
      RECT 666.500000 410.410000 699.500000 411.590000 ;
      RECT 657.500000 410.410000 658.500000 411.590000 ;
      RECT 616.500000 410.410000 649.500000 411.590000 ;
      RECT 607.500000 410.410000 608.500000 411.590000 ;
      RECT 566.500000 410.410000 599.500000 411.590000 ;
      RECT 557.500000 410.410000 558.500000 411.590000 ;
      RECT 516.500000 410.410000 549.500000 411.590000 ;
      RECT 507.500000 410.410000 508.500000 411.590000 ;
      RECT 416.500000 410.410000 499.500000 411.590000 ;
      RECT 407.500000 410.410000 408.500000 411.590000 ;
      RECT 366.500000 410.410000 399.500000 411.590000 ;
      RECT 357.500000 410.410000 358.500000 411.590000 ;
      RECT 316.500000 410.410000 349.500000 411.590000 ;
      RECT 307.500000 410.410000 308.500000 411.590000 ;
      RECT 216.500000 410.410000 299.500000 411.590000 ;
      RECT 207.500000 410.410000 208.500000 411.590000 ;
      RECT 116.500000 410.410000 199.500000 411.590000 ;
      RECT 107.500000 410.410000 108.500000 411.590000 ;
      RECT 66.500000 410.410000 99.500000 411.590000 ;
      RECT 57.500000 410.410000 58.500000 411.590000 ;
      RECT 29.500000 410.410000 49.500000 411.590000 ;
      RECT 15.500000 410.410000 16.500000 411.590000 ;
      RECT 1157.500000 409.590000 1170.500000 410.410000 ;
      RECT 1107.500000 409.590000 1149.500000 410.410000 ;
      RECT 1057.500000 409.590000 1099.500000 410.410000 ;
      RECT 1007.500000 409.590000 1049.500000 410.410000 ;
      RECT 957.500000 409.590000 999.500000 410.410000 ;
      RECT 907.500000 409.590000 949.500000 410.410000 ;
      RECT 857.500000 409.590000 899.500000 410.410000 ;
      RECT 807.500000 409.590000 849.500000 410.410000 ;
      RECT 757.500000 409.590000 799.500000 410.410000 ;
      RECT 707.500000 409.590000 749.500000 410.410000 ;
      RECT 657.500000 409.590000 699.500000 410.410000 ;
      RECT 607.500000 409.590000 649.500000 410.410000 ;
      RECT 557.500000 409.590000 599.500000 410.410000 ;
      RECT 507.500000 409.590000 549.500000 410.410000 ;
      RECT 407.500000 409.590000 499.500000 410.410000 ;
      RECT 357.500000 409.590000 399.500000 410.410000 ;
      RECT 307.500000 409.590000 349.500000 410.410000 ;
      RECT 207.500000 409.590000 299.500000 410.410000 ;
      RECT 107.500000 409.590000 199.500000 410.410000 ;
      RECT 57.500000 409.590000 99.500000 410.410000 ;
      RECT 15.500000 409.590000 49.500000 410.410000 ;
      RECT 1183.500000 408.410000 1186.000000 411.590000 ;
      RECT 1169.500000 408.410000 1170.500000 409.590000 ;
      RECT 1116.500000 408.410000 1149.500000 409.590000 ;
      RECT 1107.500000 408.410000 1108.500000 409.590000 ;
      RECT 1066.500000 408.410000 1099.500000 409.590000 ;
      RECT 1057.500000 408.410000 1058.500000 409.590000 ;
      RECT 1016.500000 408.410000 1049.500000 409.590000 ;
      RECT 1007.500000 408.410000 1008.500000 409.590000 ;
      RECT 966.500000 408.410000 999.500000 409.590000 ;
      RECT 957.500000 408.410000 958.500000 409.590000 ;
      RECT 916.500000 408.410000 949.500000 409.590000 ;
      RECT 907.500000 408.410000 908.500000 409.590000 ;
      RECT 866.500000 408.410000 899.500000 409.590000 ;
      RECT 857.500000 408.410000 858.500000 409.590000 ;
      RECT 816.500000 408.410000 849.500000 409.590000 ;
      RECT 807.500000 408.410000 808.500000 409.590000 ;
      RECT 766.500000 408.410000 799.500000 409.590000 ;
      RECT 757.500000 408.410000 758.500000 409.590000 ;
      RECT 716.500000 408.410000 749.500000 409.590000 ;
      RECT 707.500000 408.410000 708.500000 409.590000 ;
      RECT 666.500000 408.410000 699.500000 409.590000 ;
      RECT 657.500000 408.410000 658.500000 409.590000 ;
      RECT 616.500000 408.410000 649.500000 409.590000 ;
      RECT 607.500000 408.410000 608.500000 409.590000 ;
      RECT 566.500000 408.410000 599.500000 409.590000 ;
      RECT 557.500000 408.410000 558.500000 409.590000 ;
      RECT 516.500000 408.410000 549.500000 409.590000 ;
      RECT 507.500000 408.410000 508.500000 409.590000 ;
      RECT 416.500000 408.410000 499.500000 409.590000 ;
      RECT 407.500000 408.410000 408.500000 409.590000 ;
      RECT 366.500000 408.410000 399.500000 409.590000 ;
      RECT 357.500000 408.410000 358.500000 409.590000 ;
      RECT 316.500000 408.410000 349.500000 409.590000 ;
      RECT 307.500000 408.410000 308.500000 409.590000 ;
      RECT 266.500000 408.410000 299.500000 409.590000 ;
      RECT 207.500000 408.410000 208.500000 409.590000 ;
      RECT 166.500000 408.410000 199.500000 409.590000 ;
      RECT 107.500000 408.410000 108.500000 409.590000 ;
      RECT 66.500000 408.410000 99.500000 409.590000 ;
      RECT 57.500000 408.410000 58.500000 409.590000 ;
      RECT 29.500000 408.410000 49.500000 409.590000 ;
      RECT 15.500000 408.410000 16.500000 409.590000 ;
      RECT 0.000000 408.410000 2.500000 411.590000 ;
      RECT 1169.500000 407.590000 1186.000000 408.410000 ;
      RECT 1116.500000 407.590000 1156.500000 408.410000 ;
      RECT 1066.500000 407.590000 1108.500000 408.410000 ;
      RECT 1016.500000 407.590000 1058.500000 408.410000 ;
      RECT 966.500000 407.590000 1008.500000 408.410000 ;
      RECT 916.500000 407.590000 958.500000 408.410000 ;
      RECT 866.500000 407.590000 908.500000 408.410000 ;
      RECT 816.500000 407.590000 858.500000 408.410000 ;
      RECT 766.500000 407.590000 808.500000 408.410000 ;
      RECT 716.500000 407.590000 758.500000 408.410000 ;
      RECT 666.500000 407.590000 708.500000 408.410000 ;
      RECT 616.500000 407.590000 658.500000 408.410000 ;
      RECT 566.500000 407.590000 608.500000 408.410000 ;
      RECT 516.500000 407.590000 558.500000 408.410000 ;
      RECT 416.500000 407.590000 508.500000 408.410000 ;
      RECT 366.500000 407.590000 408.500000 408.410000 ;
      RECT 316.500000 407.590000 358.500000 408.410000 ;
      RECT 266.500000 407.590000 308.500000 408.410000 ;
      RECT 216.500000 407.590000 258.500000 409.590000 ;
      RECT 166.500000 407.590000 208.500000 408.410000 ;
      RECT 116.500000 407.590000 158.500000 409.590000 ;
      RECT 66.500000 407.590000 108.500000 408.410000 ;
      RECT 29.500000 407.590000 58.500000 408.410000 ;
      RECT 0.000000 407.590000 16.500000 408.410000 ;
      RECT 1169.500000 406.410000 1170.500000 407.590000 ;
      RECT 1116.500000 406.410000 1149.500000 407.590000 ;
      RECT 1107.500000 406.410000 1108.500000 407.590000 ;
      RECT 1066.500000 406.410000 1099.500000 407.590000 ;
      RECT 1057.500000 406.410000 1058.500000 407.590000 ;
      RECT 1016.500000 406.410000 1049.500000 407.590000 ;
      RECT 1007.500000 406.410000 1008.500000 407.590000 ;
      RECT 966.500000 406.410000 999.500000 407.590000 ;
      RECT 957.500000 406.410000 958.500000 407.590000 ;
      RECT 916.500000 406.410000 949.500000 407.590000 ;
      RECT 907.500000 406.410000 908.500000 407.590000 ;
      RECT 866.500000 406.410000 899.500000 407.590000 ;
      RECT 857.500000 406.410000 858.500000 407.590000 ;
      RECT 816.500000 406.410000 849.500000 407.590000 ;
      RECT 807.500000 406.410000 808.500000 407.590000 ;
      RECT 766.500000 406.410000 799.500000 407.590000 ;
      RECT 757.500000 406.410000 758.500000 407.590000 ;
      RECT 716.500000 406.410000 749.500000 407.590000 ;
      RECT 707.500000 406.410000 708.500000 407.590000 ;
      RECT 666.500000 406.410000 699.500000 407.590000 ;
      RECT 657.500000 406.410000 658.500000 407.590000 ;
      RECT 616.500000 406.410000 649.500000 407.590000 ;
      RECT 607.500000 406.410000 608.500000 407.590000 ;
      RECT 566.500000 406.410000 599.500000 407.590000 ;
      RECT 557.500000 406.410000 558.500000 407.590000 ;
      RECT 516.500000 406.410000 549.500000 407.590000 ;
      RECT 507.500000 406.410000 508.500000 407.590000 ;
      RECT 416.500000 406.410000 499.500000 407.590000 ;
      RECT 407.500000 406.410000 408.500000 407.590000 ;
      RECT 366.500000 406.410000 399.500000 407.590000 ;
      RECT 357.500000 406.410000 358.500000 407.590000 ;
      RECT 316.500000 406.410000 349.500000 407.590000 ;
      RECT 307.500000 406.410000 308.500000 407.590000 ;
      RECT 266.500000 406.410000 299.500000 407.590000 ;
      RECT 257.500000 406.410000 258.500000 407.590000 ;
      RECT 216.500000 406.410000 249.500000 407.590000 ;
      RECT 207.500000 406.410000 208.500000 407.590000 ;
      RECT 166.500000 406.410000 199.500000 407.590000 ;
      RECT 157.500000 406.410000 158.500000 407.590000 ;
      RECT 116.500000 406.410000 149.500000 407.590000 ;
      RECT 107.500000 406.410000 108.500000 407.590000 ;
      RECT 66.500000 406.410000 99.500000 407.590000 ;
      RECT 57.500000 406.410000 58.500000 407.590000 ;
      RECT 29.500000 406.410000 49.500000 407.590000 ;
      RECT 15.500000 406.410000 16.500000 407.590000 ;
      RECT 1157.500000 405.590000 1170.500000 406.410000 ;
      RECT 1107.500000 405.590000 1149.500000 406.410000 ;
      RECT 1057.500000 405.590000 1099.500000 406.410000 ;
      RECT 1007.500000 405.590000 1049.500000 406.410000 ;
      RECT 957.500000 405.590000 999.500000 406.410000 ;
      RECT 907.500000 405.590000 949.500000 406.410000 ;
      RECT 857.500000 405.590000 899.500000 406.410000 ;
      RECT 807.500000 405.590000 849.500000 406.410000 ;
      RECT 757.500000 405.590000 799.500000 406.410000 ;
      RECT 707.500000 405.590000 749.500000 406.410000 ;
      RECT 657.500000 405.590000 699.500000 406.410000 ;
      RECT 607.500000 405.590000 649.500000 406.410000 ;
      RECT 557.500000 405.590000 599.500000 406.410000 ;
      RECT 507.500000 405.590000 549.500000 406.410000 ;
      RECT 407.500000 405.590000 499.500000 406.410000 ;
      RECT 357.500000 405.590000 399.500000 406.410000 ;
      RECT 307.500000 405.590000 349.500000 406.410000 ;
      RECT 257.500000 405.590000 299.500000 406.410000 ;
      RECT 207.500000 405.590000 249.500000 406.410000 ;
      RECT 157.500000 405.590000 199.500000 406.410000 ;
      RECT 107.500000 405.590000 149.500000 406.410000 ;
      RECT 57.500000 405.590000 99.500000 406.410000 ;
      RECT 15.500000 405.590000 49.500000 406.410000 ;
      RECT 1183.500000 404.410000 1186.000000 407.590000 ;
      RECT 1169.500000 404.410000 1170.500000 405.590000 ;
      RECT 1116.500000 404.410000 1149.500000 405.590000 ;
      RECT 1107.500000 404.410000 1108.500000 405.590000 ;
      RECT 1066.500000 404.410000 1099.500000 405.590000 ;
      RECT 1057.500000 404.410000 1058.500000 405.590000 ;
      RECT 1016.500000 404.410000 1049.500000 405.590000 ;
      RECT 1007.500000 404.410000 1008.500000 405.590000 ;
      RECT 966.500000 404.410000 999.500000 405.590000 ;
      RECT 957.500000 404.410000 958.500000 405.590000 ;
      RECT 916.500000 404.410000 949.500000 405.590000 ;
      RECT 907.500000 404.410000 908.500000 405.590000 ;
      RECT 866.500000 404.410000 899.500000 405.590000 ;
      RECT 857.500000 404.410000 858.500000 405.590000 ;
      RECT 816.500000 404.410000 849.500000 405.590000 ;
      RECT 807.500000 404.410000 808.500000 405.590000 ;
      RECT 766.500000 404.410000 799.500000 405.590000 ;
      RECT 757.500000 404.410000 758.500000 405.590000 ;
      RECT 716.500000 404.410000 749.500000 405.590000 ;
      RECT 707.500000 404.410000 708.500000 405.590000 ;
      RECT 666.500000 404.410000 699.500000 405.590000 ;
      RECT 657.500000 404.410000 658.500000 405.590000 ;
      RECT 616.500000 404.410000 649.500000 405.590000 ;
      RECT 607.500000 404.410000 608.500000 405.590000 ;
      RECT 566.500000 404.410000 599.500000 405.590000 ;
      RECT 557.500000 404.410000 558.500000 405.590000 ;
      RECT 516.500000 404.410000 549.500000 405.590000 ;
      RECT 507.500000 404.410000 508.500000 405.590000 ;
      RECT 416.500000 404.410000 499.500000 405.590000 ;
      RECT 407.500000 404.410000 408.500000 405.590000 ;
      RECT 366.500000 404.410000 399.500000 405.590000 ;
      RECT 357.500000 404.410000 358.500000 405.590000 ;
      RECT 316.500000 404.410000 349.500000 405.590000 ;
      RECT 307.500000 404.410000 308.500000 405.590000 ;
      RECT 266.500000 404.410000 299.500000 405.590000 ;
      RECT 257.500000 404.410000 258.500000 405.590000 ;
      RECT 216.500000 404.410000 249.500000 405.590000 ;
      RECT 207.500000 404.410000 208.500000 405.590000 ;
      RECT 166.500000 404.410000 199.500000 405.590000 ;
      RECT 157.500000 404.410000 158.500000 405.590000 ;
      RECT 116.500000 404.410000 149.500000 405.590000 ;
      RECT 107.500000 404.410000 108.500000 405.590000 ;
      RECT 66.500000 404.410000 99.500000 405.590000 ;
      RECT 57.500000 404.410000 58.500000 405.590000 ;
      RECT 29.500000 404.410000 49.500000 405.590000 ;
      RECT 15.500000 404.410000 16.500000 405.590000 ;
      RECT 0.000000 404.410000 2.500000 407.590000 ;
      RECT 1169.500000 403.590000 1186.000000 404.410000 ;
      RECT 1116.500000 403.590000 1156.500000 404.410000 ;
      RECT 1066.500000 403.590000 1108.500000 404.410000 ;
      RECT 1016.500000 403.590000 1058.500000 404.410000 ;
      RECT 966.500000 403.590000 1008.500000 404.410000 ;
      RECT 916.500000 403.590000 958.500000 404.410000 ;
      RECT 866.500000 403.590000 908.500000 404.410000 ;
      RECT 816.500000 403.590000 858.500000 404.410000 ;
      RECT 766.500000 403.590000 808.500000 404.410000 ;
      RECT 716.500000 403.590000 758.500000 404.410000 ;
      RECT 666.500000 403.590000 708.500000 404.410000 ;
      RECT 616.500000 403.590000 658.500000 404.410000 ;
      RECT 566.500000 403.590000 608.500000 404.410000 ;
      RECT 516.500000 403.590000 558.500000 404.410000 ;
      RECT 416.500000 403.590000 508.500000 404.410000 ;
      RECT 366.500000 403.590000 408.500000 404.410000 ;
      RECT 316.500000 403.590000 358.500000 404.410000 ;
      RECT 266.500000 403.590000 308.500000 404.410000 ;
      RECT 216.500000 403.590000 258.500000 404.410000 ;
      RECT 166.500000 403.590000 208.500000 404.410000 ;
      RECT 116.500000 403.590000 158.500000 404.410000 ;
      RECT 66.500000 403.590000 108.500000 404.410000 ;
      RECT 29.500000 403.590000 58.500000 404.410000 ;
      RECT 0.000000 403.590000 16.500000 404.410000 ;
      RECT 1169.500000 402.410000 1170.500000 403.590000 ;
      RECT 1116.500000 402.410000 1149.500000 403.590000 ;
      RECT 1107.500000 402.410000 1108.500000 403.590000 ;
      RECT 1066.500000 402.410000 1099.500000 403.590000 ;
      RECT 1057.500000 402.410000 1058.500000 403.590000 ;
      RECT 1016.500000 402.410000 1049.500000 403.590000 ;
      RECT 1007.500000 402.410000 1008.500000 403.590000 ;
      RECT 966.500000 402.410000 999.500000 403.590000 ;
      RECT 957.500000 402.410000 958.500000 403.590000 ;
      RECT 916.500000 402.410000 949.500000 403.590000 ;
      RECT 907.500000 402.410000 908.500000 403.590000 ;
      RECT 866.500000 402.410000 899.500000 403.590000 ;
      RECT 857.500000 402.410000 858.500000 403.590000 ;
      RECT 816.500000 402.410000 849.500000 403.590000 ;
      RECT 807.500000 402.410000 808.500000 403.590000 ;
      RECT 766.500000 402.410000 799.500000 403.590000 ;
      RECT 757.500000 402.410000 758.500000 403.590000 ;
      RECT 716.500000 402.410000 749.500000 403.590000 ;
      RECT 707.500000 402.410000 708.500000 403.590000 ;
      RECT 666.500000 402.410000 699.500000 403.590000 ;
      RECT 657.500000 402.410000 658.500000 403.590000 ;
      RECT 616.500000 402.410000 649.500000 403.590000 ;
      RECT 607.500000 402.410000 608.500000 403.590000 ;
      RECT 566.500000 402.410000 599.500000 403.590000 ;
      RECT 557.500000 402.410000 558.500000 403.590000 ;
      RECT 516.500000 402.410000 549.500000 403.590000 ;
      RECT 507.500000 402.410000 508.500000 403.590000 ;
      RECT 416.500000 402.410000 499.500000 403.590000 ;
      RECT 407.500000 402.410000 408.500000 403.590000 ;
      RECT 366.500000 402.410000 399.500000 403.590000 ;
      RECT 357.500000 402.410000 358.500000 403.590000 ;
      RECT 316.500000 402.410000 349.500000 403.590000 ;
      RECT 307.500000 402.410000 308.500000 403.590000 ;
      RECT 266.500000 402.410000 299.500000 403.590000 ;
      RECT 257.500000 402.410000 258.500000 403.590000 ;
      RECT 216.500000 402.410000 249.500000 403.590000 ;
      RECT 207.500000 402.410000 208.500000 403.590000 ;
      RECT 166.500000 402.410000 199.500000 403.590000 ;
      RECT 157.500000 402.410000 158.500000 403.590000 ;
      RECT 116.500000 402.410000 149.500000 403.590000 ;
      RECT 107.500000 402.410000 108.500000 403.590000 ;
      RECT 66.500000 402.410000 99.500000 403.590000 ;
      RECT 57.500000 402.410000 58.500000 403.590000 ;
      RECT 29.500000 402.410000 49.500000 403.590000 ;
      RECT 15.500000 402.410000 16.500000 403.590000 ;
      RECT 1157.500000 401.590000 1170.500000 402.410000 ;
      RECT 1107.500000 401.590000 1149.500000 402.410000 ;
      RECT 1057.500000 401.590000 1099.500000 402.410000 ;
      RECT 1007.500000 401.590000 1049.500000 402.410000 ;
      RECT 957.500000 401.590000 999.500000 402.410000 ;
      RECT 907.500000 401.590000 949.500000 402.410000 ;
      RECT 857.500000 401.590000 899.500000 402.410000 ;
      RECT 807.500000 401.590000 849.500000 402.410000 ;
      RECT 757.500000 401.590000 799.500000 402.410000 ;
      RECT 707.500000 401.590000 749.500000 402.410000 ;
      RECT 657.500000 401.590000 699.500000 402.410000 ;
      RECT 607.500000 401.590000 649.500000 402.410000 ;
      RECT 557.500000 401.590000 599.500000 402.410000 ;
      RECT 507.500000 401.590000 549.500000 402.410000 ;
      RECT 407.500000 401.590000 499.500000 402.410000 ;
      RECT 357.500000 401.590000 399.500000 402.410000 ;
      RECT 307.500000 401.590000 349.500000 402.410000 ;
      RECT 257.500000 401.590000 299.500000 402.410000 ;
      RECT 207.500000 401.590000 249.500000 402.410000 ;
      RECT 157.500000 401.590000 199.500000 402.410000 ;
      RECT 107.500000 401.590000 149.500000 402.410000 ;
      RECT 57.500000 401.590000 99.500000 402.410000 ;
      RECT 15.500000 401.590000 49.500000 402.410000 ;
      RECT 1183.500000 400.410000 1186.000000 403.590000 ;
      RECT 1169.500000 400.410000 1170.500000 401.590000 ;
      RECT 1116.500000 400.410000 1149.500000 401.590000 ;
      RECT 1107.500000 400.410000 1108.500000 401.590000 ;
      RECT 1066.500000 400.410000 1099.500000 401.590000 ;
      RECT 1057.500000 400.410000 1058.500000 401.590000 ;
      RECT 1016.500000 400.410000 1049.500000 401.590000 ;
      RECT 1007.500000 400.410000 1008.500000 401.590000 ;
      RECT 966.500000 400.410000 999.500000 401.590000 ;
      RECT 957.500000 400.410000 958.500000 401.590000 ;
      RECT 916.500000 400.410000 949.500000 401.590000 ;
      RECT 907.500000 400.410000 908.500000 401.590000 ;
      RECT 866.500000 400.410000 899.500000 401.590000 ;
      RECT 857.500000 400.410000 858.500000 401.590000 ;
      RECT 816.500000 400.410000 849.500000 401.590000 ;
      RECT 807.500000 400.410000 808.500000 401.590000 ;
      RECT 766.500000 400.410000 799.500000 401.590000 ;
      RECT 757.500000 400.410000 758.500000 401.590000 ;
      RECT 716.500000 400.410000 749.500000 401.590000 ;
      RECT 707.500000 400.410000 708.500000 401.590000 ;
      RECT 666.500000 400.410000 699.500000 401.590000 ;
      RECT 657.500000 400.410000 658.500000 401.590000 ;
      RECT 616.500000 400.410000 649.500000 401.590000 ;
      RECT 607.500000 400.410000 608.500000 401.590000 ;
      RECT 566.500000 400.410000 599.500000 401.590000 ;
      RECT 557.500000 400.410000 558.500000 401.590000 ;
      RECT 516.500000 400.410000 549.500000 401.590000 ;
      RECT 507.500000 400.410000 508.500000 401.590000 ;
      RECT 416.500000 400.410000 499.500000 401.590000 ;
      RECT 407.500000 400.410000 408.500000 401.590000 ;
      RECT 366.500000 400.410000 399.500000 401.590000 ;
      RECT 357.500000 400.410000 358.500000 401.590000 ;
      RECT 316.500000 400.410000 349.500000 401.590000 ;
      RECT 307.500000 400.410000 308.500000 401.590000 ;
      RECT 266.500000 400.410000 299.500000 401.590000 ;
      RECT 257.500000 400.410000 258.500000 401.590000 ;
      RECT 216.500000 400.410000 249.500000 401.590000 ;
      RECT 207.500000 400.410000 208.500000 401.590000 ;
      RECT 166.500000 400.410000 199.500000 401.590000 ;
      RECT 157.500000 400.410000 158.500000 401.590000 ;
      RECT 116.500000 400.410000 149.500000 401.590000 ;
      RECT 107.500000 400.410000 108.500000 401.590000 ;
      RECT 66.500000 400.410000 99.500000 401.590000 ;
      RECT 57.500000 400.410000 58.500000 401.590000 ;
      RECT 29.500000 400.410000 49.500000 401.590000 ;
      RECT 15.500000 400.410000 16.500000 401.590000 ;
      RECT 0.000000 400.410000 2.500000 403.590000 ;
      RECT 1169.500000 399.590000 1186.000000 400.410000 ;
      RECT 1116.500000 399.590000 1156.500000 400.410000 ;
      RECT 1066.500000 399.590000 1108.500000 400.410000 ;
      RECT 1016.500000 399.590000 1058.500000 400.410000 ;
      RECT 966.500000 399.590000 1008.500000 400.410000 ;
      RECT 916.500000 399.590000 958.500000 400.410000 ;
      RECT 866.500000 399.590000 908.500000 400.410000 ;
      RECT 816.500000 399.590000 858.500000 400.410000 ;
      RECT 766.500000 399.590000 808.500000 400.410000 ;
      RECT 716.500000 399.590000 758.500000 400.410000 ;
      RECT 666.500000 399.590000 708.500000 400.410000 ;
      RECT 616.500000 399.590000 658.500000 400.410000 ;
      RECT 566.500000 399.590000 608.500000 400.410000 ;
      RECT 516.500000 399.590000 558.500000 400.410000 ;
      RECT 416.500000 399.590000 508.500000 400.410000 ;
      RECT 366.500000 399.590000 408.500000 400.410000 ;
      RECT 316.500000 399.590000 358.500000 400.410000 ;
      RECT 266.500000 399.590000 308.500000 400.410000 ;
      RECT 216.500000 399.590000 258.500000 400.410000 ;
      RECT 166.500000 399.590000 208.500000 400.410000 ;
      RECT 116.500000 399.590000 158.500000 400.410000 ;
      RECT 66.500000 399.590000 108.500000 400.410000 ;
      RECT 29.500000 399.590000 58.500000 400.410000 ;
      RECT 0.000000 399.590000 16.500000 400.410000 ;
      RECT 0.000000 399.170000 2.500000 399.590000 ;
      RECT 1183.500000 399.165000 1186.000000 399.590000 ;
      RECT 1169.500000 398.410000 1170.500000 399.590000 ;
      RECT 1116.500000 398.410000 1149.500000 399.590000 ;
      RECT 1107.500000 398.410000 1108.500000 399.590000 ;
      RECT 1066.500000 398.410000 1099.500000 399.590000 ;
      RECT 1057.500000 398.410000 1058.500000 399.590000 ;
      RECT 1016.500000 398.410000 1049.500000 399.590000 ;
      RECT 1007.500000 398.410000 1008.500000 399.590000 ;
      RECT 966.500000 398.410000 999.500000 399.590000 ;
      RECT 957.500000 398.410000 958.500000 399.590000 ;
      RECT 916.500000 398.410000 949.500000 399.590000 ;
      RECT 907.500000 398.410000 908.500000 399.590000 ;
      RECT 866.500000 398.410000 899.500000 399.590000 ;
      RECT 857.500000 398.410000 858.500000 399.590000 ;
      RECT 816.500000 398.410000 849.500000 399.590000 ;
      RECT 807.500000 398.410000 808.500000 399.590000 ;
      RECT 766.500000 398.410000 799.500000 399.590000 ;
      RECT 757.500000 398.410000 758.500000 399.590000 ;
      RECT 716.500000 398.410000 749.500000 399.590000 ;
      RECT 707.500000 398.410000 708.500000 399.590000 ;
      RECT 666.500000 398.410000 699.500000 399.590000 ;
      RECT 657.500000 398.410000 658.500000 399.590000 ;
      RECT 616.500000 398.410000 649.500000 399.590000 ;
      RECT 607.500000 398.410000 608.500000 399.590000 ;
      RECT 566.500000 398.410000 599.500000 399.590000 ;
      RECT 557.500000 398.410000 558.500000 399.590000 ;
      RECT 516.500000 398.410000 549.500000 399.590000 ;
      RECT 507.500000 398.410000 508.500000 399.590000 ;
      RECT 416.500000 398.410000 449.500000 399.590000 ;
      RECT 407.500000 398.410000 408.500000 399.590000 ;
      RECT 366.500000 398.410000 399.500000 399.590000 ;
      RECT 357.500000 398.410000 358.500000 399.590000 ;
      RECT 316.500000 398.410000 349.500000 399.590000 ;
      RECT 307.500000 398.410000 308.500000 399.590000 ;
      RECT 266.500000 398.410000 299.500000 399.590000 ;
      RECT 257.500000 398.410000 258.500000 399.590000 ;
      RECT 216.500000 398.410000 249.500000 399.590000 ;
      RECT 207.500000 398.410000 208.500000 399.590000 ;
      RECT 166.500000 398.410000 199.500000 399.590000 ;
      RECT 157.500000 398.410000 158.500000 399.590000 ;
      RECT 116.500000 398.410000 149.500000 399.590000 ;
      RECT 107.500000 398.410000 108.500000 399.590000 ;
      RECT 66.500000 398.410000 99.500000 399.590000 ;
      RECT 57.500000 398.410000 58.500000 399.590000 ;
      RECT 29.500000 398.410000 49.500000 399.590000 ;
      RECT 15.500000 398.410000 16.500000 399.590000 ;
      RECT 1157.500000 397.590000 1170.500000 398.410000 ;
      RECT 1107.500000 397.590000 1149.500000 398.410000 ;
      RECT 1057.500000 397.590000 1099.500000 398.410000 ;
      RECT 1007.500000 397.590000 1049.500000 398.410000 ;
      RECT 957.500000 397.590000 999.500000 398.410000 ;
      RECT 907.500000 397.590000 949.500000 398.410000 ;
      RECT 857.500000 397.590000 899.500000 398.410000 ;
      RECT 807.500000 397.590000 849.500000 398.410000 ;
      RECT 757.500000 397.590000 799.500000 398.410000 ;
      RECT 707.500000 397.590000 749.500000 398.410000 ;
      RECT 657.500000 397.590000 699.500000 398.410000 ;
      RECT 607.500000 397.590000 649.500000 398.410000 ;
      RECT 557.500000 397.590000 599.500000 398.410000 ;
      RECT 507.500000 397.590000 549.500000 398.410000 ;
      RECT 457.500000 397.590000 499.500000 399.590000 ;
      RECT 407.500000 397.590000 449.500000 398.410000 ;
      RECT 357.500000 397.590000 399.500000 398.410000 ;
      RECT 307.500000 397.590000 349.500000 398.410000 ;
      RECT 257.500000 397.590000 299.500000 398.410000 ;
      RECT 207.500000 397.590000 249.500000 398.410000 ;
      RECT 157.500000 397.590000 199.500000 398.410000 ;
      RECT 107.500000 397.590000 149.500000 398.410000 ;
      RECT 57.500000 397.590000 99.500000 398.410000 ;
      RECT 15.500000 397.590000 49.500000 398.410000 ;
      RECT 1183.500000 396.410000 1183.980000 399.165000 ;
      RECT 1169.500000 396.410000 1170.500000 397.590000 ;
      RECT 1116.500000 396.410000 1149.500000 397.590000 ;
      RECT 1107.500000 396.410000 1108.500000 397.590000 ;
      RECT 1066.500000 396.410000 1099.500000 397.590000 ;
      RECT 1057.500000 396.410000 1058.500000 397.590000 ;
      RECT 1016.500000 396.410000 1049.500000 397.590000 ;
      RECT 1007.500000 396.410000 1008.500000 397.590000 ;
      RECT 966.500000 396.410000 999.500000 397.590000 ;
      RECT 957.500000 396.410000 958.500000 397.590000 ;
      RECT 916.500000 396.410000 949.500000 397.590000 ;
      RECT 907.500000 396.410000 908.500000 397.590000 ;
      RECT 866.500000 396.410000 899.500000 397.590000 ;
      RECT 857.500000 396.410000 858.500000 397.590000 ;
      RECT 816.500000 396.410000 849.500000 397.590000 ;
      RECT 807.500000 396.410000 808.500000 397.590000 ;
      RECT 766.500000 396.410000 799.500000 397.590000 ;
      RECT 757.500000 396.410000 758.500000 397.590000 ;
      RECT 716.500000 396.410000 749.500000 397.590000 ;
      RECT 707.500000 396.410000 708.500000 397.590000 ;
      RECT 666.500000 396.410000 699.500000 397.590000 ;
      RECT 657.500000 396.410000 658.500000 397.590000 ;
      RECT 616.500000 396.410000 649.500000 397.590000 ;
      RECT 607.500000 396.410000 608.500000 397.590000 ;
      RECT 566.500000 396.410000 599.500000 397.590000 ;
      RECT 557.500000 396.410000 558.500000 397.590000 ;
      RECT 516.500000 396.410000 549.500000 397.590000 ;
      RECT 507.500000 396.410000 508.500000 397.590000 ;
      RECT 466.500000 396.410000 499.500000 397.590000 ;
      RECT 457.500000 396.410000 458.500000 397.590000 ;
      RECT 416.500000 396.410000 449.500000 397.590000 ;
      RECT 407.500000 396.410000 408.500000 397.590000 ;
      RECT 366.500000 396.410000 399.500000 397.590000 ;
      RECT 357.500000 396.410000 358.500000 397.590000 ;
      RECT 316.500000 396.410000 349.500000 397.590000 ;
      RECT 307.500000 396.410000 308.500000 397.590000 ;
      RECT 266.500000 396.410000 299.500000 397.590000 ;
      RECT 257.500000 396.410000 258.500000 397.590000 ;
      RECT 216.500000 396.410000 249.500000 397.590000 ;
      RECT 207.500000 396.410000 208.500000 397.590000 ;
      RECT 166.500000 396.410000 199.500000 397.590000 ;
      RECT 157.500000 396.410000 158.500000 397.590000 ;
      RECT 116.500000 396.410000 149.500000 397.590000 ;
      RECT 107.500000 396.410000 108.500000 397.590000 ;
      RECT 66.500000 396.410000 99.500000 397.590000 ;
      RECT 57.500000 396.410000 58.500000 397.590000 ;
      RECT 29.500000 396.410000 49.500000 397.590000 ;
      RECT 15.500000 396.410000 16.500000 397.590000 ;
      RECT 2.020000 396.410000 2.500000 399.170000 ;
      RECT 2.020000 396.070000 16.500000 396.410000 ;
      RECT 1169.500000 396.065000 1183.980000 396.410000 ;
      RECT 1169.500000 395.590000 1186.000000 396.065000 ;
      RECT 1116.500000 395.590000 1156.500000 396.410000 ;
      RECT 1066.500000 395.590000 1108.500000 396.410000 ;
      RECT 1016.500000 395.590000 1058.500000 396.410000 ;
      RECT 966.500000 395.590000 1008.500000 396.410000 ;
      RECT 916.500000 395.590000 958.500000 396.410000 ;
      RECT 866.500000 395.590000 908.500000 396.410000 ;
      RECT 816.500000 395.590000 858.500000 396.410000 ;
      RECT 766.500000 395.590000 808.500000 396.410000 ;
      RECT 716.500000 395.590000 758.500000 396.410000 ;
      RECT 666.500000 395.590000 708.500000 396.410000 ;
      RECT 616.500000 395.590000 658.500000 396.410000 ;
      RECT 566.500000 395.590000 608.500000 396.410000 ;
      RECT 516.500000 395.590000 558.500000 396.410000 ;
      RECT 466.500000 395.590000 508.500000 396.410000 ;
      RECT 416.500000 395.590000 458.500000 396.410000 ;
      RECT 366.500000 395.590000 408.500000 396.410000 ;
      RECT 316.500000 395.590000 358.500000 396.410000 ;
      RECT 266.500000 395.590000 308.500000 396.410000 ;
      RECT 216.500000 395.590000 258.500000 396.410000 ;
      RECT 166.500000 395.590000 208.500000 396.410000 ;
      RECT 116.500000 395.590000 158.500000 396.410000 ;
      RECT 66.500000 395.590000 108.500000 396.410000 ;
      RECT 29.500000 395.590000 58.500000 396.410000 ;
      RECT 0.000000 395.590000 16.500000 396.070000 ;
      RECT 1169.500000 394.410000 1170.500000 395.590000 ;
      RECT 1116.500000 394.410000 1149.500000 395.590000 ;
      RECT 1107.500000 394.410000 1108.500000 395.590000 ;
      RECT 1066.500000 394.410000 1099.500000 395.590000 ;
      RECT 1057.500000 394.410000 1058.500000 395.590000 ;
      RECT 1016.500000 394.410000 1049.500000 395.590000 ;
      RECT 1007.500000 394.410000 1008.500000 395.590000 ;
      RECT 966.500000 394.410000 999.500000 395.590000 ;
      RECT 957.500000 394.410000 958.500000 395.590000 ;
      RECT 916.500000 394.410000 949.500000 395.590000 ;
      RECT 907.500000 394.410000 908.500000 395.590000 ;
      RECT 866.500000 394.410000 899.500000 395.590000 ;
      RECT 857.500000 394.410000 858.500000 395.590000 ;
      RECT 816.500000 394.410000 849.500000 395.590000 ;
      RECT 807.500000 394.410000 808.500000 395.590000 ;
      RECT 766.500000 394.410000 799.500000 395.590000 ;
      RECT 757.500000 394.410000 758.500000 395.590000 ;
      RECT 716.500000 394.410000 749.500000 395.590000 ;
      RECT 707.500000 394.410000 708.500000 395.590000 ;
      RECT 666.500000 394.410000 699.500000 395.590000 ;
      RECT 657.500000 394.410000 658.500000 395.590000 ;
      RECT 616.500000 394.410000 649.500000 395.590000 ;
      RECT 607.500000 394.410000 608.500000 395.590000 ;
      RECT 566.500000 394.410000 599.500000 395.590000 ;
      RECT 557.500000 394.410000 558.500000 395.590000 ;
      RECT 516.500000 394.410000 549.500000 395.590000 ;
      RECT 507.500000 394.410000 508.500000 395.590000 ;
      RECT 466.500000 394.410000 499.500000 395.590000 ;
      RECT 457.500000 394.410000 458.500000 395.590000 ;
      RECT 416.500000 394.410000 449.500000 395.590000 ;
      RECT 407.500000 394.410000 408.500000 395.590000 ;
      RECT 366.500000 394.410000 399.500000 395.590000 ;
      RECT 357.500000 394.410000 358.500000 395.590000 ;
      RECT 316.500000 394.410000 349.500000 395.590000 ;
      RECT 307.500000 394.410000 308.500000 395.590000 ;
      RECT 266.500000 394.410000 299.500000 395.590000 ;
      RECT 257.500000 394.410000 258.500000 395.590000 ;
      RECT 216.500000 394.410000 249.500000 395.590000 ;
      RECT 207.500000 394.410000 208.500000 395.590000 ;
      RECT 166.500000 394.410000 199.500000 395.590000 ;
      RECT 157.500000 394.410000 158.500000 395.590000 ;
      RECT 116.500000 394.410000 149.500000 395.590000 ;
      RECT 107.500000 394.410000 108.500000 395.590000 ;
      RECT 66.500000 394.410000 99.500000 395.590000 ;
      RECT 57.500000 394.410000 58.500000 395.590000 ;
      RECT 29.500000 394.410000 49.500000 395.590000 ;
      RECT 15.500000 394.410000 16.500000 395.590000 ;
      RECT 1157.500000 393.590000 1170.500000 394.410000 ;
      RECT 1107.500000 393.590000 1149.500000 394.410000 ;
      RECT 1057.500000 393.590000 1099.500000 394.410000 ;
      RECT 1007.500000 393.590000 1049.500000 394.410000 ;
      RECT 957.500000 393.590000 999.500000 394.410000 ;
      RECT 907.500000 393.590000 949.500000 394.410000 ;
      RECT 857.500000 393.590000 899.500000 394.410000 ;
      RECT 807.500000 393.590000 849.500000 394.410000 ;
      RECT 757.500000 393.590000 799.500000 394.410000 ;
      RECT 707.500000 393.590000 749.500000 394.410000 ;
      RECT 657.500000 393.590000 699.500000 394.410000 ;
      RECT 607.500000 393.590000 649.500000 394.410000 ;
      RECT 557.500000 393.590000 599.500000 394.410000 ;
      RECT 507.500000 393.590000 549.500000 394.410000 ;
      RECT 457.500000 393.590000 499.500000 394.410000 ;
      RECT 407.500000 393.590000 449.500000 394.410000 ;
      RECT 357.500000 393.590000 399.500000 394.410000 ;
      RECT 307.500000 393.590000 349.500000 394.410000 ;
      RECT 257.500000 393.590000 299.500000 394.410000 ;
      RECT 207.500000 393.590000 249.500000 394.410000 ;
      RECT 157.500000 393.590000 199.500000 394.410000 ;
      RECT 107.500000 393.590000 149.500000 394.410000 ;
      RECT 57.500000 393.590000 99.500000 394.410000 ;
      RECT 15.500000 393.590000 49.500000 394.410000 ;
      RECT 1183.500000 393.485000 1186.000000 395.590000 ;
      RECT 1183.500000 392.410000 1183.980000 393.485000 ;
      RECT 1169.500000 392.410000 1170.500000 393.590000 ;
      RECT 1116.500000 392.410000 1149.500000 393.590000 ;
      RECT 1107.500000 392.410000 1108.500000 393.590000 ;
      RECT 1066.500000 392.410000 1099.500000 393.590000 ;
      RECT 1057.500000 392.410000 1058.500000 393.590000 ;
      RECT 1016.500000 392.410000 1049.500000 393.590000 ;
      RECT 1007.500000 392.410000 1008.500000 393.590000 ;
      RECT 966.500000 392.410000 999.500000 393.590000 ;
      RECT 957.500000 392.410000 958.500000 393.590000 ;
      RECT 916.500000 392.410000 949.500000 393.590000 ;
      RECT 907.500000 392.410000 908.500000 393.590000 ;
      RECT 866.500000 392.410000 899.500000 393.590000 ;
      RECT 857.500000 392.410000 858.500000 393.590000 ;
      RECT 816.500000 392.410000 849.500000 393.590000 ;
      RECT 807.500000 392.410000 808.500000 393.590000 ;
      RECT 766.500000 392.410000 799.500000 393.590000 ;
      RECT 757.500000 392.410000 758.500000 393.590000 ;
      RECT 716.500000 392.410000 749.500000 393.590000 ;
      RECT 707.500000 392.410000 708.500000 393.590000 ;
      RECT 666.500000 392.410000 699.500000 393.590000 ;
      RECT 657.500000 392.410000 658.500000 393.590000 ;
      RECT 616.500000 392.410000 649.500000 393.590000 ;
      RECT 607.500000 392.410000 608.500000 393.590000 ;
      RECT 566.500000 392.410000 599.500000 393.590000 ;
      RECT 557.500000 392.410000 558.500000 393.590000 ;
      RECT 516.500000 392.410000 549.500000 393.590000 ;
      RECT 507.500000 392.410000 508.500000 393.590000 ;
      RECT 466.500000 392.410000 499.500000 393.590000 ;
      RECT 457.500000 392.410000 458.500000 393.590000 ;
      RECT 416.500000 392.410000 449.500000 393.590000 ;
      RECT 407.500000 392.410000 408.500000 393.590000 ;
      RECT 366.500000 392.410000 399.500000 393.590000 ;
      RECT 357.500000 392.410000 358.500000 393.590000 ;
      RECT 316.500000 392.410000 349.500000 393.590000 ;
      RECT 307.500000 392.410000 308.500000 393.590000 ;
      RECT 266.500000 392.410000 299.500000 393.590000 ;
      RECT 257.500000 392.410000 258.500000 393.590000 ;
      RECT 216.500000 392.410000 249.500000 393.590000 ;
      RECT 207.500000 392.410000 208.500000 393.590000 ;
      RECT 166.500000 392.410000 199.500000 393.590000 ;
      RECT 157.500000 392.410000 158.500000 393.590000 ;
      RECT 116.500000 392.410000 149.500000 393.590000 ;
      RECT 107.500000 392.410000 108.500000 393.590000 ;
      RECT 66.500000 392.410000 99.500000 393.590000 ;
      RECT 57.500000 392.410000 58.500000 393.590000 ;
      RECT 29.500000 392.410000 49.500000 393.590000 ;
      RECT 15.500000 392.410000 16.500000 393.590000 ;
      RECT 0.000000 392.410000 2.500000 395.590000 ;
      RECT 1169.500000 391.590000 1183.980000 392.410000 ;
      RECT 1116.500000 391.590000 1156.500000 392.410000 ;
      RECT 1066.500000 391.590000 1108.500000 392.410000 ;
      RECT 1016.500000 391.590000 1058.500000 392.410000 ;
      RECT 966.500000 391.590000 1008.500000 392.410000 ;
      RECT 916.500000 391.590000 958.500000 392.410000 ;
      RECT 866.500000 391.590000 908.500000 392.410000 ;
      RECT 816.500000 391.590000 858.500000 392.410000 ;
      RECT 766.500000 391.590000 808.500000 392.410000 ;
      RECT 716.500000 391.590000 758.500000 392.410000 ;
      RECT 666.500000 391.590000 708.500000 392.410000 ;
      RECT 616.500000 391.590000 658.500000 392.410000 ;
      RECT 566.500000 391.590000 608.500000 392.410000 ;
      RECT 516.500000 391.590000 558.500000 392.410000 ;
      RECT 466.500000 391.590000 508.500000 392.410000 ;
      RECT 416.500000 391.590000 458.500000 392.410000 ;
      RECT 366.500000 391.590000 408.500000 392.410000 ;
      RECT 316.500000 391.590000 358.500000 392.410000 ;
      RECT 266.500000 391.590000 308.500000 392.410000 ;
      RECT 216.500000 391.590000 258.500000 392.410000 ;
      RECT 166.500000 391.590000 208.500000 392.410000 ;
      RECT 116.500000 391.590000 158.500000 392.410000 ;
      RECT 66.500000 391.590000 108.500000 392.410000 ;
      RECT 29.500000 391.590000 58.500000 392.410000 ;
      RECT 0.000000 391.590000 16.500000 392.410000 ;
      RECT 1169.500000 390.410000 1170.500000 391.590000 ;
      RECT 1116.500000 390.410000 1149.500000 391.590000 ;
      RECT 1107.500000 390.410000 1108.500000 391.590000 ;
      RECT 1066.500000 390.410000 1099.500000 391.590000 ;
      RECT 1057.500000 390.410000 1058.500000 391.590000 ;
      RECT 1016.500000 390.410000 1049.500000 391.590000 ;
      RECT 1007.500000 390.410000 1008.500000 391.590000 ;
      RECT 966.500000 390.410000 999.500000 391.590000 ;
      RECT 957.500000 390.410000 958.500000 391.590000 ;
      RECT 916.500000 390.410000 949.500000 391.590000 ;
      RECT 907.500000 390.410000 908.500000 391.590000 ;
      RECT 866.500000 390.410000 899.500000 391.590000 ;
      RECT 857.500000 390.410000 858.500000 391.590000 ;
      RECT 816.500000 390.410000 849.500000 391.590000 ;
      RECT 807.500000 390.410000 808.500000 391.590000 ;
      RECT 766.500000 390.410000 799.500000 391.590000 ;
      RECT 757.500000 390.410000 758.500000 391.590000 ;
      RECT 716.500000 390.410000 749.500000 391.590000 ;
      RECT 707.500000 390.410000 708.500000 391.590000 ;
      RECT 666.500000 390.410000 699.500000 391.590000 ;
      RECT 657.500000 390.410000 658.500000 391.590000 ;
      RECT 616.500000 390.410000 649.500000 391.590000 ;
      RECT 607.500000 390.410000 608.500000 391.590000 ;
      RECT 566.500000 390.410000 599.500000 391.590000 ;
      RECT 557.500000 390.410000 558.500000 391.590000 ;
      RECT 516.500000 390.410000 549.500000 391.590000 ;
      RECT 507.500000 390.410000 508.500000 391.590000 ;
      RECT 466.500000 390.410000 499.500000 391.590000 ;
      RECT 457.500000 390.410000 458.500000 391.590000 ;
      RECT 416.500000 390.410000 449.500000 391.590000 ;
      RECT 407.500000 390.410000 408.500000 391.590000 ;
      RECT 366.500000 390.410000 399.500000 391.590000 ;
      RECT 357.500000 390.410000 358.500000 391.590000 ;
      RECT 316.500000 390.410000 349.500000 391.590000 ;
      RECT 307.500000 390.410000 308.500000 391.590000 ;
      RECT 266.500000 390.410000 299.500000 391.590000 ;
      RECT 257.500000 390.410000 258.500000 391.590000 ;
      RECT 216.500000 390.410000 249.500000 391.590000 ;
      RECT 207.500000 390.410000 208.500000 391.590000 ;
      RECT 166.500000 390.410000 199.500000 391.590000 ;
      RECT 157.500000 390.410000 158.500000 391.590000 ;
      RECT 116.500000 390.410000 149.500000 391.590000 ;
      RECT 107.500000 390.410000 108.500000 391.590000 ;
      RECT 66.500000 390.410000 99.500000 391.590000 ;
      RECT 57.500000 390.410000 58.500000 391.590000 ;
      RECT 29.500000 390.410000 49.500000 391.590000 ;
      RECT 15.500000 390.410000 16.500000 391.590000 ;
      RECT 1183.500000 390.385000 1183.980000 391.590000 ;
      RECT 1157.500000 389.590000 1170.500000 390.410000 ;
      RECT 1107.500000 389.590000 1149.500000 390.410000 ;
      RECT 1057.500000 389.590000 1099.500000 390.410000 ;
      RECT 1007.500000 389.590000 1049.500000 390.410000 ;
      RECT 957.500000 389.590000 999.500000 390.410000 ;
      RECT 907.500000 389.590000 949.500000 390.410000 ;
      RECT 857.500000 389.590000 899.500000 390.410000 ;
      RECT 807.500000 389.590000 849.500000 390.410000 ;
      RECT 757.500000 389.590000 799.500000 390.410000 ;
      RECT 707.500000 389.590000 749.500000 390.410000 ;
      RECT 657.500000 389.590000 699.500000 390.410000 ;
      RECT 607.500000 389.590000 649.500000 390.410000 ;
      RECT 557.500000 389.590000 599.500000 390.410000 ;
      RECT 507.500000 389.590000 549.500000 390.410000 ;
      RECT 457.500000 389.590000 499.500000 390.410000 ;
      RECT 407.500000 389.590000 449.500000 390.410000 ;
      RECT 357.500000 389.590000 399.500000 390.410000 ;
      RECT 307.500000 389.590000 349.500000 390.410000 ;
      RECT 257.500000 389.590000 299.500000 390.410000 ;
      RECT 207.500000 389.590000 249.500000 390.410000 ;
      RECT 157.500000 389.590000 199.500000 390.410000 ;
      RECT 107.500000 389.590000 149.500000 390.410000 ;
      RECT 57.500000 389.590000 99.500000 390.410000 ;
      RECT 15.500000 389.590000 49.500000 390.410000 ;
      RECT 1183.500000 389.525000 1186.000000 390.385000 ;
      RECT 0.000000 388.575000 2.500000 391.590000 ;
      RECT 1183.500000 388.410000 1183.980000 389.525000 ;
      RECT 1169.500000 388.410000 1170.500000 389.590000 ;
      RECT 1116.500000 388.410000 1149.500000 389.590000 ;
      RECT 1107.500000 388.410000 1108.500000 389.590000 ;
      RECT 1066.500000 388.410000 1099.500000 389.590000 ;
      RECT 1057.500000 388.410000 1058.500000 389.590000 ;
      RECT 1016.500000 388.410000 1049.500000 389.590000 ;
      RECT 1007.500000 388.410000 1008.500000 389.590000 ;
      RECT 966.500000 388.410000 999.500000 389.590000 ;
      RECT 957.500000 388.410000 958.500000 389.590000 ;
      RECT 916.500000 388.410000 949.500000 389.590000 ;
      RECT 907.500000 388.410000 908.500000 389.590000 ;
      RECT 866.500000 388.410000 899.500000 389.590000 ;
      RECT 857.500000 388.410000 858.500000 389.590000 ;
      RECT 816.500000 388.410000 849.500000 389.590000 ;
      RECT 807.500000 388.410000 808.500000 389.590000 ;
      RECT 766.500000 388.410000 799.500000 389.590000 ;
      RECT 757.500000 388.410000 758.500000 389.590000 ;
      RECT 716.500000 388.410000 749.500000 389.590000 ;
      RECT 707.500000 388.410000 708.500000 389.590000 ;
      RECT 666.500000 388.410000 699.500000 389.590000 ;
      RECT 657.500000 388.410000 658.500000 389.590000 ;
      RECT 616.500000 388.410000 649.500000 389.590000 ;
      RECT 607.500000 388.410000 608.500000 389.590000 ;
      RECT 566.500000 388.410000 599.500000 389.590000 ;
      RECT 557.500000 388.410000 558.500000 389.590000 ;
      RECT 516.500000 388.410000 549.500000 389.590000 ;
      RECT 507.500000 388.410000 508.500000 389.590000 ;
      RECT 466.500000 388.410000 499.500000 389.590000 ;
      RECT 457.500000 388.410000 458.500000 389.590000 ;
      RECT 416.500000 388.410000 449.500000 389.590000 ;
      RECT 407.500000 388.410000 408.500000 389.590000 ;
      RECT 366.500000 388.410000 399.500000 389.590000 ;
      RECT 357.500000 388.410000 358.500000 389.590000 ;
      RECT 316.500000 388.410000 349.500000 389.590000 ;
      RECT 307.500000 388.410000 308.500000 389.590000 ;
      RECT 266.500000 388.410000 299.500000 389.590000 ;
      RECT 257.500000 388.410000 258.500000 389.590000 ;
      RECT 216.500000 388.410000 249.500000 389.590000 ;
      RECT 207.500000 388.410000 208.500000 389.590000 ;
      RECT 166.500000 388.410000 199.500000 389.590000 ;
      RECT 157.500000 388.410000 158.500000 389.590000 ;
      RECT 116.500000 388.410000 149.500000 389.590000 ;
      RECT 107.500000 388.410000 108.500000 389.590000 ;
      RECT 66.500000 388.410000 99.500000 389.590000 ;
      RECT 57.500000 388.410000 58.500000 389.590000 ;
      RECT 29.500000 388.410000 49.500000 389.590000 ;
      RECT 15.500000 388.410000 16.500000 389.590000 ;
      RECT 2.020000 388.410000 2.500000 388.575000 ;
      RECT 1169.500000 387.590000 1183.980000 388.410000 ;
      RECT 1116.500000 387.590000 1156.500000 388.410000 ;
      RECT 1066.500000 387.590000 1108.500000 388.410000 ;
      RECT 1016.500000 387.590000 1058.500000 388.410000 ;
      RECT 966.500000 387.590000 1008.500000 388.410000 ;
      RECT 916.500000 387.590000 958.500000 388.410000 ;
      RECT 866.500000 387.590000 908.500000 388.410000 ;
      RECT 816.500000 387.590000 858.500000 388.410000 ;
      RECT 766.500000 387.590000 808.500000 388.410000 ;
      RECT 716.500000 387.590000 758.500000 388.410000 ;
      RECT 666.500000 387.590000 708.500000 388.410000 ;
      RECT 616.500000 387.590000 658.500000 388.410000 ;
      RECT 566.500000 387.590000 608.500000 388.410000 ;
      RECT 516.500000 387.590000 558.500000 388.410000 ;
      RECT 466.500000 387.590000 508.500000 388.410000 ;
      RECT 416.500000 387.590000 458.500000 388.410000 ;
      RECT 366.500000 387.590000 408.500000 388.410000 ;
      RECT 316.500000 387.590000 358.500000 388.410000 ;
      RECT 266.500000 387.590000 308.500000 388.410000 ;
      RECT 216.500000 387.590000 258.500000 388.410000 ;
      RECT 166.500000 387.590000 208.500000 388.410000 ;
      RECT 116.500000 387.590000 158.500000 388.410000 ;
      RECT 66.500000 387.590000 108.500000 388.410000 ;
      RECT 29.500000 387.590000 58.500000 388.410000 ;
      RECT 2.020000 387.590000 16.500000 388.410000 ;
      RECT 1183.500000 386.425000 1183.980000 387.590000 ;
      RECT 1169.500000 386.410000 1170.500000 387.590000 ;
      RECT 1116.500000 386.410000 1149.500000 387.590000 ;
      RECT 1107.500000 386.410000 1108.500000 387.590000 ;
      RECT 1066.500000 386.410000 1099.500000 387.590000 ;
      RECT 1057.500000 386.410000 1058.500000 387.590000 ;
      RECT 1016.500000 386.410000 1049.500000 387.590000 ;
      RECT 1007.500000 386.410000 1008.500000 387.590000 ;
      RECT 966.500000 386.410000 999.500000 387.590000 ;
      RECT 957.500000 386.410000 958.500000 387.590000 ;
      RECT 916.500000 386.410000 949.500000 387.590000 ;
      RECT 907.500000 386.410000 908.500000 387.590000 ;
      RECT 866.500000 386.410000 899.500000 387.590000 ;
      RECT 857.500000 386.410000 858.500000 387.590000 ;
      RECT 816.500000 386.410000 849.500000 387.590000 ;
      RECT 807.500000 386.410000 808.500000 387.590000 ;
      RECT 766.500000 386.410000 799.500000 387.590000 ;
      RECT 757.500000 386.410000 758.500000 387.590000 ;
      RECT 716.500000 386.410000 749.500000 387.590000 ;
      RECT 707.500000 386.410000 708.500000 387.590000 ;
      RECT 666.500000 386.410000 699.500000 387.590000 ;
      RECT 657.500000 386.410000 658.500000 387.590000 ;
      RECT 616.500000 386.410000 649.500000 387.590000 ;
      RECT 607.500000 386.410000 608.500000 387.590000 ;
      RECT 566.500000 386.410000 599.500000 387.590000 ;
      RECT 557.500000 386.410000 558.500000 387.590000 ;
      RECT 516.500000 386.410000 549.500000 387.590000 ;
      RECT 507.500000 386.410000 508.500000 387.590000 ;
      RECT 466.500000 386.410000 499.500000 387.590000 ;
      RECT 457.500000 386.410000 458.500000 387.590000 ;
      RECT 416.500000 386.410000 449.500000 387.590000 ;
      RECT 407.500000 386.410000 408.500000 387.590000 ;
      RECT 366.500000 386.410000 399.500000 387.590000 ;
      RECT 357.500000 386.410000 358.500000 387.590000 ;
      RECT 316.500000 386.410000 349.500000 387.590000 ;
      RECT 307.500000 386.410000 308.500000 387.590000 ;
      RECT 266.500000 386.410000 299.500000 387.590000 ;
      RECT 257.500000 386.410000 258.500000 387.590000 ;
      RECT 216.500000 386.410000 249.500000 387.590000 ;
      RECT 207.500000 386.410000 208.500000 387.590000 ;
      RECT 166.500000 386.410000 199.500000 387.590000 ;
      RECT 157.500000 386.410000 158.500000 387.590000 ;
      RECT 116.500000 386.410000 149.500000 387.590000 ;
      RECT 107.500000 386.410000 108.500000 387.590000 ;
      RECT 66.500000 386.410000 99.500000 387.590000 ;
      RECT 57.500000 386.410000 58.500000 387.590000 ;
      RECT 29.500000 386.410000 49.500000 387.590000 ;
      RECT 15.500000 386.410000 16.500000 387.590000 ;
      RECT 1157.500000 385.590000 1170.500000 386.410000 ;
      RECT 1107.500000 385.590000 1149.500000 386.410000 ;
      RECT 1057.500000 385.590000 1099.500000 386.410000 ;
      RECT 1007.500000 385.590000 1049.500000 386.410000 ;
      RECT 957.500000 385.590000 999.500000 386.410000 ;
      RECT 907.500000 385.590000 949.500000 386.410000 ;
      RECT 857.500000 385.590000 899.500000 386.410000 ;
      RECT 807.500000 385.590000 849.500000 386.410000 ;
      RECT 757.500000 385.590000 799.500000 386.410000 ;
      RECT 707.500000 385.590000 749.500000 386.410000 ;
      RECT 657.500000 385.590000 699.500000 386.410000 ;
      RECT 607.500000 385.590000 649.500000 386.410000 ;
      RECT 557.500000 385.590000 599.500000 386.410000 ;
      RECT 507.500000 385.590000 549.500000 386.410000 ;
      RECT 457.500000 385.590000 499.500000 386.410000 ;
      RECT 407.500000 385.590000 449.500000 386.410000 ;
      RECT 357.500000 385.590000 399.500000 386.410000 ;
      RECT 307.500000 385.590000 349.500000 386.410000 ;
      RECT 257.500000 385.590000 299.500000 386.410000 ;
      RECT 207.500000 385.590000 249.500000 386.410000 ;
      RECT 157.500000 385.590000 199.500000 386.410000 ;
      RECT 107.500000 385.590000 149.500000 386.410000 ;
      RECT 57.500000 385.590000 99.500000 386.410000 ;
      RECT 15.500000 385.590000 49.500000 386.410000 ;
      RECT 2.020000 385.475000 2.500000 387.590000 ;
      RECT 0.000000 384.615000 2.500000 385.475000 ;
      RECT 1183.500000 384.410000 1186.000000 386.425000 ;
      RECT 1169.500000 384.410000 1170.500000 385.590000 ;
      RECT 1116.500000 384.410000 1149.500000 385.590000 ;
      RECT 1107.500000 384.410000 1108.500000 385.590000 ;
      RECT 1066.500000 384.410000 1099.500000 385.590000 ;
      RECT 1057.500000 384.410000 1058.500000 385.590000 ;
      RECT 1016.500000 384.410000 1049.500000 385.590000 ;
      RECT 1007.500000 384.410000 1008.500000 385.590000 ;
      RECT 966.500000 384.410000 999.500000 385.590000 ;
      RECT 957.500000 384.410000 958.500000 385.590000 ;
      RECT 916.500000 384.410000 949.500000 385.590000 ;
      RECT 907.500000 384.410000 908.500000 385.590000 ;
      RECT 866.500000 384.410000 899.500000 385.590000 ;
      RECT 857.500000 384.410000 858.500000 385.590000 ;
      RECT 816.500000 384.410000 849.500000 385.590000 ;
      RECT 807.500000 384.410000 808.500000 385.590000 ;
      RECT 766.500000 384.410000 799.500000 385.590000 ;
      RECT 757.500000 384.410000 758.500000 385.590000 ;
      RECT 716.500000 384.410000 749.500000 385.590000 ;
      RECT 707.500000 384.410000 708.500000 385.590000 ;
      RECT 666.500000 384.410000 699.500000 385.590000 ;
      RECT 657.500000 384.410000 658.500000 385.590000 ;
      RECT 616.500000 384.410000 649.500000 385.590000 ;
      RECT 607.500000 384.410000 608.500000 385.590000 ;
      RECT 566.500000 384.410000 599.500000 385.590000 ;
      RECT 557.500000 384.410000 558.500000 385.590000 ;
      RECT 516.500000 384.410000 549.500000 385.590000 ;
      RECT 507.500000 384.410000 508.500000 385.590000 ;
      RECT 466.500000 384.410000 499.500000 385.590000 ;
      RECT 457.500000 384.410000 458.500000 385.590000 ;
      RECT 416.500000 384.410000 449.500000 385.590000 ;
      RECT 407.500000 384.410000 408.500000 385.590000 ;
      RECT 366.500000 384.410000 399.500000 385.590000 ;
      RECT 357.500000 384.410000 358.500000 385.590000 ;
      RECT 316.500000 384.410000 349.500000 385.590000 ;
      RECT 307.500000 384.410000 308.500000 385.590000 ;
      RECT 266.500000 384.410000 299.500000 385.590000 ;
      RECT 257.500000 384.410000 258.500000 385.590000 ;
      RECT 216.500000 384.410000 249.500000 385.590000 ;
      RECT 207.500000 384.410000 208.500000 385.590000 ;
      RECT 166.500000 384.410000 199.500000 385.590000 ;
      RECT 157.500000 384.410000 158.500000 385.590000 ;
      RECT 116.500000 384.410000 149.500000 385.590000 ;
      RECT 107.500000 384.410000 108.500000 385.590000 ;
      RECT 66.500000 384.410000 99.500000 385.590000 ;
      RECT 57.500000 384.410000 58.500000 385.590000 ;
      RECT 29.500000 384.410000 49.500000 385.590000 ;
      RECT 15.500000 384.410000 16.500000 385.590000 ;
      RECT 2.020000 384.410000 2.500000 384.615000 ;
      RECT 1169.500000 383.590000 1186.000000 384.410000 ;
      RECT 1116.500000 383.590000 1156.500000 384.410000 ;
      RECT 1066.500000 383.590000 1108.500000 384.410000 ;
      RECT 1016.500000 383.590000 1058.500000 384.410000 ;
      RECT 966.500000 383.590000 1008.500000 384.410000 ;
      RECT 916.500000 383.590000 958.500000 384.410000 ;
      RECT 866.500000 383.590000 908.500000 384.410000 ;
      RECT 816.500000 383.590000 858.500000 384.410000 ;
      RECT 766.500000 383.590000 808.500000 384.410000 ;
      RECT 716.500000 383.590000 758.500000 384.410000 ;
      RECT 666.500000 383.590000 708.500000 384.410000 ;
      RECT 616.500000 383.590000 658.500000 384.410000 ;
      RECT 566.500000 383.590000 608.500000 384.410000 ;
      RECT 516.500000 383.590000 558.500000 384.410000 ;
      RECT 466.500000 383.590000 508.500000 384.410000 ;
      RECT 416.500000 383.590000 458.500000 384.410000 ;
      RECT 366.500000 383.590000 408.500000 384.410000 ;
      RECT 316.500000 383.590000 358.500000 384.410000 ;
      RECT 266.500000 383.590000 308.500000 384.410000 ;
      RECT 216.500000 383.590000 258.500000 384.410000 ;
      RECT 166.500000 383.590000 208.500000 384.410000 ;
      RECT 116.500000 383.590000 158.500000 384.410000 ;
      RECT 66.500000 383.590000 108.500000 384.410000 ;
      RECT 29.500000 383.590000 58.500000 384.410000 ;
      RECT 2.020000 383.590000 16.500000 384.410000 ;
      RECT 1169.500000 382.410000 1170.500000 383.590000 ;
      RECT 1116.500000 382.410000 1149.500000 383.590000 ;
      RECT 1107.500000 382.410000 1108.500000 383.590000 ;
      RECT 1066.500000 382.410000 1099.500000 383.590000 ;
      RECT 1057.500000 382.410000 1058.500000 383.590000 ;
      RECT 1016.500000 382.410000 1049.500000 383.590000 ;
      RECT 1007.500000 382.410000 1008.500000 383.590000 ;
      RECT 966.500000 382.410000 999.500000 383.590000 ;
      RECT 957.500000 382.410000 958.500000 383.590000 ;
      RECT 916.500000 382.410000 949.500000 383.590000 ;
      RECT 907.500000 382.410000 908.500000 383.590000 ;
      RECT 866.500000 382.410000 899.500000 383.590000 ;
      RECT 857.500000 382.410000 858.500000 383.590000 ;
      RECT 816.500000 382.410000 849.500000 383.590000 ;
      RECT 807.500000 382.410000 808.500000 383.590000 ;
      RECT 766.500000 382.410000 799.500000 383.590000 ;
      RECT 757.500000 382.410000 758.500000 383.590000 ;
      RECT 716.500000 382.410000 749.500000 383.590000 ;
      RECT 707.500000 382.410000 708.500000 383.590000 ;
      RECT 666.500000 382.410000 699.500000 383.590000 ;
      RECT 657.500000 382.410000 658.500000 383.590000 ;
      RECT 616.500000 382.410000 649.500000 383.590000 ;
      RECT 607.500000 382.410000 608.500000 383.590000 ;
      RECT 566.500000 382.410000 599.500000 383.590000 ;
      RECT 557.500000 382.410000 558.500000 383.590000 ;
      RECT 516.500000 382.410000 549.500000 383.590000 ;
      RECT 507.500000 382.410000 508.500000 383.590000 ;
      RECT 466.500000 382.410000 499.500000 383.590000 ;
      RECT 457.500000 382.410000 458.500000 383.590000 ;
      RECT 416.500000 382.410000 449.500000 383.590000 ;
      RECT 407.500000 382.410000 408.500000 383.590000 ;
      RECT 366.500000 382.410000 399.500000 383.590000 ;
      RECT 357.500000 382.410000 358.500000 383.590000 ;
      RECT 316.500000 382.410000 349.500000 383.590000 ;
      RECT 307.500000 382.410000 308.500000 383.590000 ;
      RECT 266.500000 382.410000 299.500000 383.590000 ;
      RECT 257.500000 382.410000 258.500000 383.590000 ;
      RECT 216.500000 382.410000 249.500000 383.590000 ;
      RECT 207.500000 382.410000 208.500000 383.590000 ;
      RECT 166.500000 382.410000 199.500000 383.590000 ;
      RECT 157.500000 382.410000 158.500000 383.590000 ;
      RECT 116.500000 382.410000 149.500000 383.590000 ;
      RECT 107.500000 382.410000 108.500000 383.590000 ;
      RECT 66.500000 382.410000 99.500000 383.590000 ;
      RECT 57.500000 382.410000 58.500000 383.590000 ;
      RECT 29.500000 382.410000 49.500000 383.590000 ;
      RECT 15.500000 382.410000 16.500000 383.590000 ;
      RECT 1157.500000 381.590000 1170.500000 382.410000 ;
      RECT 1107.500000 381.590000 1149.500000 382.410000 ;
      RECT 1057.500000 381.590000 1099.500000 382.410000 ;
      RECT 1007.500000 381.590000 1049.500000 382.410000 ;
      RECT 957.500000 381.590000 999.500000 382.410000 ;
      RECT 907.500000 381.590000 949.500000 382.410000 ;
      RECT 857.500000 381.590000 899.500000 382.410000 ;
      RECT 807.500000 381.590000 849.500000 382.410000 ;
      RECT 757.500000 381.590000 799.500000 382.410000 ;
      RECT 707.500000 381.590000 749.500000 382.410000 ;
      RECT 657.500000 381.590000 699.500000 382.410000 ;
      RECT 607.500000 381.590000 649.500000 382.410000 ;
      RECT 557.500000 381.590000 599.500000 382.410000 ;
      RECT 507.500000 381.590000 549.500000 382.410000 ;
      RECT 457.500000 381.590000 499.500000 382.410000 ;
      RECT 407.500000 381.590000 449.500000 382.410000 ;
      RECT 357.500000 381.590000 399.500000 382.410000 ;
      RECT 307.500000 381.590000 349.500000 382.410000 ;
      RECT 257.500000 381.590000 299.500000 382.410000 ;
      RECT 207.500000 381.590000 249.500000 382.410000 ;
      RECT 157.500000 381.590000 199.500000 382.410000 ;
      RECT 107.500000 381.590000 149.500000 382.410000 ;
      RECT 57.500000 381.590000 99.500000 382.410000 ;
      RECT 15.500000 381.590000 49.500000 382.410000 ;
      RECT 2.020000 381.515000 2.500000 383.590000 ;
      RECT 1183.500000 380.410000 1186.000000 383.590000 ;
      RECT 1169.500000 380.410000 1170.500000 381.590000 ;
      RECT 1116.500000 380.410000 1149.500000 381.590000 ;
      RECT 1107.500000 380.410000 1108.500000 381.590000 ;
      RECT 1066.500000 380.410000 1099.500000 381.590000 ;
      RECT 1057.500000 380.410000 1058.500000 381.590000 ;
      RECT 1016.500000 380.410000 1049.500000 381.590000 ;
      RECT 1007.500000 380.410000 1008.500000 381.590000 ;
      RECT 966.500000 380.410000 999.500000 381.590000 ;
      RECT 957.500000 380.410000 958.500000 381.590000 ;
      RECT 916.500000 380.410000 949.500000 381.590000 ;
      RECT 907.500000 380.410000 908.500000 381.590000 ;
      RECT 866.500000 380.410000 899.500000 381.590000 ;
      RECT 857.500000 380.410000 858.500000 381.590000 ;
      RECT 816.500000 380.410000 849.500000 381.590000 ;
      RECT 807.500000 380.410000 808.500000 381.590000 ;
      RECT 766.500000 380.410000 799.500000 381.590000 ;
      RECT 757.500000 380.410000 758.500000 381.590000 ;
      RECT 716.500000 380.410000 749.500000 381.590000 ;
      RECT 707.500000 380.410000 708.500000 381.590000 ;
      RECT 666.500000 380.410000 699.500000 381.590000 ;
      RECT 657.500000 380.410000 658.500000 381.590000 ;
      RECT 616.500000 380.410000 649.500000 381.590000 ;
      RECT 607.500000 380.410000 608.500000 381.590000 ;
      RECT 566.500000 380.410000 599.500000 381.590000 ;
      RECT 557.500000 380.410000 558.500000 381.590000 ;
      RECT 516.500000 380.410000 549.500000 381.590000 ;
      RECT 507.500000 380.410000 508.500000 381.590000 ;
      RECT 466.500000 380.410000 499.500000 381.590000 ;
      RECT 457.500000 380.410000 458.500000 381.590000 ;
      RECT 416.500000 380.410000 449.500000 381.590000 ;
      RECT 407.500000 380.410000 408.500000 381.590000 ;
      RECT 366.500000 380.410000 399.500000 381.590000 ;
      RECT 357.500000 380.410000 358.500000 381.590000 ;
      RECT 316.500000 380.410000 349.500000 381.590000 ;
      RECT 307.500000 380.410000 308.500000 381.590000 ;
      RECT 266.500000 380.410000 299.500000 381.590000 ;
      RECT 257.500000 380.410000 258.500000 381.590000 ;
      RECT 216.500000 380.410000 249.500000 381.590000 ;
      RECT 207.500000 380.410000 208.500000 381.590000 ;
      RECT 166.500000 380.410000 199.500000 381.590000 ;
      RECT 157.500000 380.410000 158.500000 381.590000 ;
      RECT 116.500000 380.410000 149.500000 381.590000 ;
      RECT 107.500000 380.410000 108.500000 381.590000 ;
      RECT 66.500000 380.410000 99.500000 381.590000 ;
      RECT 57.500000 380.410000 58.500000 381.590000 ;
      RECT 29.500000 380.410000 49.500000 381.590000 ;
      RECT 15.500000 380.410000 16.500000 381.590000 ;
      RECT 0.000000 380.410000 2.500000 381.515000 ;
      RECT 1169.500000 379.590000 1186.000000 380.410000 ;
      RECT 1116.500000 379.590000 1156.500000 380.410000 ;
      RECT 1066.500000 379.590000 1108.500000 380.410000 ;
      RECT 1016.500000 379.590000 1058.500000 380.410000 ;
      RECT 966.500000 379.590000 1008.500000 380.410000 ;
      RECT 916.500000 379.590000 958.500000 380.410000 ;
      RECT 866.500000 379.590000 908.500000 380.410000 ;
      RECT 816.500000 379.590000 858.500000 380.410000 ;
      RECT 766.500000 379.590000 808.500000 380.410000 ;
      RECT 716.500000 379.590000 758.500000 380.410000 ;
      RECT 666.500000 379.590000 708.500000 380.410000 ;
      RECT 616.500000 379.590000 658.500000 380.410000 ;
      RECT 566.500000 379.590000 608.500000 380.410000 ;
      RECT 516.500000 379.590000 558.500000 380.410000 ;
      RECT 466.500000 379.590000 508.500000 380.410000 ;
      RECT 416.500000 379.590000 458.500000 380.410000 ;
      RECT 366.500000 379.590000 408.500000 380.410000 ;
      RECT 316.500000 379.590000 358.500000 380.410000 ;
      RECT 266.500000 379.590000 308.500000 380.410000 ;
      RECT 216.500000 379.590000 258.500000 380.410000 ;
      RECT 166.500000 379.590000 208.500000 380.410000 ;
      RECT 116.500000 379.590000 158.500000 380.410000 ;
      RECT 66.500000 379.590000 108.500000 380.410000 ;
      RECT 29.500000 379.590000 58.500000 380.410000 ;
      RECT 0.000000 379.590000 16.500000 380.410000 ;
      RECT 0.000000 378.935000 2.500000 379.590000 ;
      RECT 1183.500000 378.930000 1186.000000 379.590000 ;
      RECT 1169.500000 378.410000 1170.500000 379.590000 ;
      RECT 1116.500000 378.410000 1149.500000 379.590000 ;
      RECT 1107.500000 378.410000 1108.500000 379.590000 ;
      RECT 1066.500000 378.410000 1099.500000 379.590000 ;
      RECT 1057.500000 378.410000 1058.500000 379.590000 ;
      RECT 1016.500000 378.410000 1049.500000 379.590000 ;
      RECT 1007.500000 378.410000 1008.500000 379.590000 ;
      RECT 966.500000 378.410000 999.500000 379.590000 ;
      RECT 957.500000 378.410000 958.500000 379.590000 ;
      RECT 916.500000 378.410000 949.500000 379.590000 ;
      RECT 907.500000 378.410000 908.500000 379.590000 ;
      RECT 866.500000 378.410000 899.500000 379.590000 ;
      RECT 857.500000 378.410000 858.500000 379.590000 ;
      RECT 816.500000 378.410000 849.500000 379.590000 ;
      RECT 807.500000 378.410000 808.500000 379.590000 ;
      RECT 766.500000 378.410000 799.500000 379.590000 ;
      RECT 757.500000 378.410000 758.500000 379.590000 ;
      RECT 716.500000 378.410000 749.500000 379.590000 ;
      RECT 707.500000 378.410000 708.500000 379.590000 ;
      RECT 666.500000 378.410000 699.500000 379.590000 ;
      RECT 657.500000 378.410000 658.500000 379.590000 ;
      RECT 616.500000 378.410000 649.500000 379.590000 ;
      RECT 607.500000 378.410000 608.500000 379.590000 ;
      RECT 566.500000 378.410000 599.500000 379.590000 ;
      RECT 557.500000 378.410000 558.500000 379.590000 ;
      RECT 516.500000 378.410000 549.500000 379.590000 ;
      RECT 507.500000 378.410000 508.500000 379.590000 ;
      RECT 466.500000 378.410000 499.500000 379.590000 ;
      RECT 457.500000 378.410000 458.500000 379.590000 ;
      RECT 416.500000 378.410000 449.500000 379.590000 ;
      RECT 407.500000 378.410000 408.500000 379.590000 ;
      RECT 366.500000 378.410000 399.500000 379.590000 ;
      RECT 357.500000 378.410000 358.500000 379.590000 ;
      RECT 316.500000 378.410000 349.500000 379.590000 ;
      RECT 307.500000 378.410000 308.500000 379.590000 ;
      RECT 266.500000 378.410000 299.500000 379.590000 ;
      RECT 257.500000 378.410000 258.500000 379.590000 ;
      RECT 216.500000 378.410000 249.500000 379.590000 ;
      RECT 207.500000 378.410000 208.500000 379.590000 ;
      RECT 166.500000 378.410000 199.500000 379.590000 ;
      RECT 157.500000 378.410000 158.500000 379.590000 ;
      RECT 116.500000 378.410000 149.500000 379.590000 ;
      RECT 107.500000 378.410000 108.500000 379.590000 ;
      RECT 66.500000 378.410000 99.500000 379.590000 ;
      RECT 57.500000 378.410000 58.500000 379.590000 ;
      RECT 29.500000 378.410000 49.500000 379.590000 ;
      RECT 15.500000 378.410000 16.500000 379.590000 ;
      RECT 1157.500000 377.590000 1170.500000 378.410000 ;
      RECT 1107.500000 377.590000 1149.500000 378.410000 ;
      RECT 1057.500000 377.590000 1099.500000 378.410000 ;
      RECT 1007.500000 377.590000 1049.500000 378.410000 ;
      RECT 957.500000 377.590000 999.500000 378.410000 ;
      RECT 907.500000 377.590000 949.500000 378.410000 ;
      RECT 857.500000 377.590000 899.500000 378.410000 ;
      RECT 807.500000 377.590000 849.500000 378.410000 ;
      RECT 757.500000 377.590000 799.500000 378.410000 ;
      RECT 707.500000 377.590000 749.500000 378.410000 ;
      RECT 657.500000 377.590000 699.500000 378.410000 ;
      RECT 607.500000 377.590000 649.500000 378.410000 ;
      RECT 557.500000 377.590000 599.500000 378.410000 ;
      RECT 507.500000 377.590000 549.500000 378.410000 ;
      RECT 457.500000 377.590000 499.500000 378.410000 ;
      RECT 407.500000 377.590000 449.500000 378.410000 ;
      RECT 357.500000 377.590000 399.500000 378.410000 ;
      RECT 307.500000 377.590000 349.500000 378.410000 ;
      RECT 257.500000 377.590000 299.500000 378.410000 ;
      RECT 207.500000 377.590000 249.500000 378.410000 ;
      RECT 157.500000 377.590000 199.500000 378.410000 ;
      RECT 107.500000 377.590000 149.500000 378.410000 ;
      RECT 57.500000 377.590000 99.500000 378.410000 ;
      RECT 15.500000 377.590000 49.500000 378.410000 ;
      RECT 1183.500000 376.410000 1183.980000 378.930000 ;
      RECT 1169.500000 376.410000 1170.500000 377.590000 ;
      RECT 1116.500000 376.410000 1149.500000 377.590000 ;
      RECT 1107.500000 376.410000 1108.500000 377.590000 ;
      RECT 1066.500000 376.410000 1099.500000 377.590000 ;
      RECT 1057.500000 376.410000 1058.500000 377.590000 ;
      RECT 1016.500000 376.410000 1049.500000 377.590000 ;
      RECT 1007.500000 376.410000 1008.500000 377.590000 ;
      RECT 966.500000 376.410000 999.500000 377.590000 ;
      RECT 957.500000 376.410000 958.500000 377.590000 ;
      RECT 916.500000 376.410000 949.500000 377.590000 ;
      RECT 907.500000 376.410000 908.500000 377.590000 ;
      RECT 866.500000 376.410000 899.500000 377.590000 ;
      RECT 857.500000 376.410000 858.500000 377.590000 ;
      RECT 816.500000 376.410000 849.500000 377.590000 ;
      RECT 807.500000 376.410000 808.500000 377.590000 ;
      RECT 766.500000 376.410000 799.500000 377.590000 ;
      RECT 757.500000 376.410000 758.500000 377.590000 ;
      RECT 716.500000 376.410000 749.500000 377.590000 ;
      RECT 707.500000 376.410000 708.500000 377.590000 ;
      RECT 666.500000 376.410000 699.500000 377.590000 ;
      RECT 657.500000 376.410000 658.500000 377.590000 ;
      RECT 616.500000 376.410000 649.500000 377.590000 ;
      RECT 607.500000 376.410000 608.500000 377.590000 ;
      RECT 566.500000 376.410000 599.500000 377.590000 ;
      RECT 557.500000 376.410000 558.500000 377.590000 ;
      RECT 516.500000 376.410000 549.500000 377.590000 ;
      RECT 507.500000 376.410000 508.500000 377.590000 ;
      RECT 466.500000 376.410000 499.500000 377.590000 ;
      RECT 457.500000 376.410000 458.500000 377.590000 ;
      RECT 416.500000 376.410000 449.500000 377.590000 ;
      RECT 407.500000 376.410000 408.500000 377.590000 ;
      RECT 366.500000 376.410000 399.500000 377.590000 ;
      RECT 357.500000 376.410000 358.500000 377.590000 ;
      RECT 316.500000 376.410000 349.500000 377.590000 ;
      RECT 307.500000 376.410000 308.500000 377.590000 ;
      RECT 266.500000 376.410000 299.500000 377.590000 ;
      RECT 257.500000 376.410000 258.500000 377.590000 ;
      RECT 216.500000 376.410000 249.500000 377.590000 ;
      RECT 207.500000 376.410000 208.500000 377.590000 ;
      RECT 166.500000 376.410000 199.500000 377.590000 ;
      RECT 157.500000 376.410000 158.500000 377.590000 ;
      RECT 116.500000 376.410000 149.500000 377.590000 ;
      RECT 107.500000 376.410000 108.500000 377.590000 ;
      RECT 66.500000 376.410000 99.500000 377.590000 ;
      RECT 57.500000 376.410000 58.500000 377.590000 ;
      RECT 29.500000 376.410000 49.500000 377.590000 ;
      RECT 15.500000 376.410000 16.500000 377.590000 ;
      RECT 2.020000 376.410000 2.500000 378.935000 ;
      RECT 2.020000 375.835000 16.500000 376.410000 ;
      RECT 1169.500000 375.830000 1183.980000 376.410000 ;
      RECT 1169.500000 375.590000 1186.000000 375.830000 ;
      RECT 1116.500000 375.590000 1156.500000 376.410000 ;
      RECT 1066.500000 375.590000 1108.500000 376.410000 ;
      RECT 1016.500000 375.590000 1058.500000 376.410000 ;
      RECT 966.500000 375.590000 1008.500000 376.410000 ;
      RECT 916.500000 375.590000 958.500000 376.410000 ;
      RECT 866.500000 375.590000 908.500000 376.410000 ;
      RECT 816.500000 375.590000 858.500000 376.410000 ;
      RECT 766.500000 375.590000 808.500000 376.410000 ;
      RECT 716.500000 375.590000 758.500000 376.410000 ;
      RECT 666.500000 375.590000 708.500000 376.410000 ;
      RECT 616.500000 375.590000 658.500000 376.410000 ;
      RECT 566.500000 375.590000 608.500000 376.410000 ;
      RECT 516.500000 375.590000 558.500000 376.410000 ;
      RECT 466.500000 375.590000 508.500000 376.410000 ;
      RECT 416.500000 375.590000 458.500000 376.410000 ;
      RECT 366.500000 375.590000 408.500000 376.410000 ;
      RECT 316.500000 375.590000 358.500000 376.410000 ;
      RECT 266.500000 375.590000 308.500000 376.410000 ;
      RECT 216.500000 375.590000 258.500000 376.410000 ;
      RECT 166.500000 375.590000 208.500000 376.410000 ;
      RECT 116.500000 375.590000 158.500000 376.410000 ;
      RECT 66.500000 375.590000 108.500000 376.410000 ;
      RECT 29.500000 375.590000 58.500000 376.410000 ;
      RECT 0.000000 375.590000 16.500000 375.835000 ;
      RECT 1169.500000 374.410000 1170.500000 375.590000 ;
      RECT 1116.500000 374.410000 1149.500000 375.590000 ;
      RECT 1107.500000 374.410000 1108.500000 375.590000 ;
      RECT 1066.500000 374.410000 1099.500000 375.590000 ;
      RECT 1057.500000 374.410000 1058.500000 375.590000 ;
      RECT 1016.500000 374.410000 1049.500000 375.590000 ;
      RECT 1007.500000 374.410000 1008.500000 375.590000 ;
      RECT 966.500000 374.410000 999.500000 375.590000 ;
      RECT 957.500000 374.410000 958.500000 375.590000 ;
      RECT 916.500000 374.410000 949.500000 375.590000 ;
      RECT 907.500000 374.410000 908.500000 375.590000 ;
      RECT 866.500000 374.410000 899.500000 375.590000 ;
      RECT 857.500000 374.410000 858.500000 375.590000 ;
      RECT 816.500000 374.410000 849.500000 375.590000 ;
      RECT 807.500000 374.410000 808.500000 375.590000 ;
      RECT 766.500000 374.410000 799.500000 375.590000 ;
      RECT 757.500000 374.410000 758.500000 375.590000 ;
      RECT 716.500000 374.410000 749.500000 375.590000 ;
      RECT 707.500000 374.410000 708.500000 375.590000 ;
      RECT 666.500000 374.410000 699.500000 375.590000 ;
      RECT 657.500000 374.410000 658.500000 375.590000 ;
      RECT 616.500000 374.410000 649.500000 375.590000 ;
      RECT 607.500000 374.410000 608.500000 375.590000 ;
      RECT 566.500000 374.410000 599.500000 375.590000 ;
      RECT 557.500000 374.410000 558.500000 375.590000 ;
      RECT 516.500000 374.410000 549.500000 375.590000 ;
      RECT 507.500000 374.410000 508.500000 375.590000 ;
      RECT 466.500000 374.410000 499.500000 375.590000 ;
      RECT 457.500000 374.410000 458.500000 375.590000 ;
      RECT 416.500000 374.410000 449.500000 375.590000 ;
      RECT 407.500000 374.410000 408.500000 375.590000 ;
      RECT 366.500000 374.410000 399.500000 375.590000 ;
      RECT 357.500000 374.410000 358.500000 375.590000 ;
      RECT 316.500000 374.410000 349.500000 375.590000 ;
      RECT 307.500000 374.410000 308.500000 375.590000 ;
      RECT 266.500000 374.410000 299.500000 375.590000 ;
      RECT 257.500000 374.410000 258.500000 375.590000 ;
      RECT 216.500000 374.410000 249.500000 375.590000 ;
      RECT 207.500000 374.410000 208.500000 375.590000 ;
      RECT 166.500000 374.410000 199.500000 375.590000 ;
      RECT 157.500000 374.410000 158.500000 375.590000 ;
      RECT 116.500000 374.410000 149.500000 375.590000 ;
      RECT 107.500000 374.410000 108.500000 375.590000 ;
      RECT 66.500000 374.410000 99.500000 375.590000 ;
      RECT 57.500000 374.410000 58.500000 375.590000 ;
      RECT 29.500000 374.410000 49.500000 375.590000 ;
      RECT 15.500000 374.410000 16.500000 375.590000 ;
      RECT 1157.500000 373.590000 1170.500000 374.410000 ;
      RECT 1107.500000 373.590000 1149.500000 374.410000 ;
      RECT 1057.500000 373.590000 1099.500000 374.410000 ;
      RECT 1007.500000 373.590000 1049.500000 374.410000 ;
      RECT 957.500000 373.590000 999.500000 374.410000 ;
      RECT 907.500000 373.590000 949.500000 374.410000 ;
      RECT 857.500000 373.590000 899.500000 374.410000 ;
      RECT 807.500000 373.590000 849.500000 374.410000 ;
      RECT 757.500000 373.590000 799.500000 374.410000 ;
      RECT 707.500000 373.590000 749.500000 374.410000 ;
      RECT 657.500000 373.590000 699.500000 374.410000 ;
      RECT 607.500000 373.590000 649.500000 374.410000 ;
      RECT 557.500000 373.590000 599.500000 374.410000 ;
      RECT 507.500000 373.590000 549.500000 374.410000 ;
      RECT 457.500000 373.590000 499.500000 374.410000 ;
      RECT 407.500000 373.590000 449.500000 374.410000 ;
      RECT 357.500000 373.590000 399.500000 374.410000 ;
      RECT 307.500000 373.590000 349.500000 374.410000 ;
      RECT 257.500000 373.590000 299.500000 374.410000 ;
      RECT 207.500000 373.590000 249.500000 374.410000 ;
      RECT 157.500000 373.590000 199.500000 374.410000 ;
      RECT 107.500000 373.590000 149.500000 374.410000 ;
      RECT 57.500000 373.590000 99.500000 374.410000 ;
      RECT 15.500000 373.590000 49.500000 374.410000 ;
      RECT 1183.500000 372.410000 1186.000000 375.590000 ;
      RECT 1169.500000 372.410000 1170.500000 373.590000 ;
      RECT 1116.500000 372.410000 1149.500000 373.590000 ;
      RECT 1107.500000 372.410000 1108.500000 373.590000 ;
      RECT 1066.500000 372.410000 1099.500000 373.590000 ;
      RECT 1057.500000 372.410000 1058.500000 373.590000 ;
      RECT 1016.500000 372.410000 1049.500000 373.590000 ;
      RECT 1007.500000 372.410000 1008.500000 373.590000 ;
      RECT 966.500000 372.410000 999.500000 373.590000 ;
      RECT 957.500000 372.410000 958.500000 373.590000 ;
      RECT 916.500000 372.410000 949.500000 373.590000 ;
      RECT 907.500000 372.410000 908.500000 373.590000 ;
      RECT 866.500000 372.410000 899.500000 373.590000 ;
      RECT 857.500000 372.410000 858.500000 373.590000 ;
      RECT 816.500000 372.410000 849.500000 373.590000 ;
      RECT 807.500000 372.410000 808.500000 373.590000 ;
      RECT 766.500000 372.410000 799.500000 373.590000 ;
      RECT 757.500000 372.410000 758.500000 373.590000 ;
      RECT 716.500000 372.410000 749.500000 373.590000 ;
      RECT 707.500000 372.410000 708.500000 373.590000 ;
      RECT 666.500000 372.410000 699.500000 373.590000 ;
      RECT 657.500000 372.410000 658.500000 373.590000 ;
      RECT 616.500000 372.410000 649.500000 373.590000 ;
      RECT 607.500000 372.410000 608.500000 373.590000 ;
      RECT 566.500000 372.410000 599.500000 373.590000 ;
      RECT 557.500000 372.410000 558.500000 373.590000 ;
      RECT 516.500000 372.410000 549.500000 373.590000 ;
      RECT 507.500000 372.410000 508.500000 373.590000 ;
      RECT 466.500000 372.410000 499.500000 373.590000 ;
      RECT 457.500000 372.410000 458.500000 373.590000 ;
      RECT 416.500000 372.410000 449.500000 373.590000 ;
      RECT 407.500000 372.410000 408.500000 373.590000 ;
      RECT 366.500000 372.410000 399.500000 373.590000 ;
      RECT 357.500000 372.410000 358.500000 373.590000 ;
      RECT 316.500000 372.410000 349.500000 373.590000 ;
      RECT 307.500000 372.410000 308.500000 373.590000 ;
      RECT 266.500000 372.410000 299.500000 373.590000 ;
      RECT 257.500000 372.410000 258.500000 373.590000 ;
      RECT 216.500000 372.410000 249.500000 373.590000 ;
      RECT 207.500000 372.410000 208.500000 373.590000 ;
      RECT 166.500000 372.410000 199.500000 373.590000 ;
      RECT 157.500000 372.410000 158.500000 373.590000 ;
      RECT 116.500000 372.410000 149.500000 373.590000 ;
      RECT 107.500000 372.410000 108.500000 373.590000 ;
      RECT 66.500000 372.410000 99.500000 373.590000 ;
      RECT 57.500000 372.410000 58.500000 373.590000 ;
      RECT 29.500000 372.410000 49.500000 373.590000 ;
      RECT 15.500000 372.410000 16.500000 373.590000 ;
      RECT 0.000000 372.410000 2.500000 375.590000 ;
      RECT 1169.500000 371.590000 1186.000000 372.410000 ;
      RECT 1116.500000 371.590000 1156.500000 372.410000 ;
      RECT 1066.500000 371.590000 1108.500000 372.410000 ;
      RECT 1016.500000 371.590000 1058.500000 372.410000 ;
      RECT 966.500000 371.590000 1008.500000 372.410000 ;
      RECT 916.500000 371.590000 958.500000 372.410000 ;
      RECT 866.500000 371.590000 908.500000 372.410000 ;
      RECT 816.500000 371.590000 858.500000 372.410000 ;
      RECT 766.500000 371.590000 808.500000 372.410000 ;
      RECT 716.500000 371.590000 758.500000 372.410000 ;
      RECT 666.500000 371.590000 708.500000 372.410000 ;
      RECT 616.500000 371.590000 658.500000 372.410000 ;
      RECT 566.500000 371.590000 608.500000 372.410000 ;
      RECT 516.500000 371.590000 558.500000 372.410000 ;
      RECT 466.500000 371.590000 508.500000 372.410000 ;
      RECT 416.500000 371.590000 458.500000 372.410000 ;
      RECT 366.500000 371.590000 408.500000 372.410000 ;
      RECT 316.500000 371.590000 358.500000 372.410000 ;
      RECT 266.500000 371.590000 308.500000 372.410000 ;
      RECT 216.500000 371.590000 258.500000 372.410000 ;
      RECT 166.500000 371.590000 208.500000 372.410000 ;
      RECT 116.500000 371.590000 158.500000 372.410000 ;
      RECT 66.500000 371.590000 108.500000 372.410000 ;
      RECT 29.500000 371.590000 58.500000 372.410000 ;
      RECT 0.000000 371.590000 16.500000 372.410000 ;
      RECT 1169.500000 370.410000 1170.500000 371.590000 ;
      RECT 1116.500000 370.410000 1149.500000 371.590000 ;
      RECT 1107.500000 370.410000 1108.500000 371.590000 ;
      RECT 1066.500000 370.410000 1099.500000 371.590000 ;
      RECT 1057.500000 370.410000 1058.500000 371.590000 ;
      RECT 1016.500000 370.410000 1049.500000 371.590000 ;
      RECT 1007.500000 370.410000 1008.500000 371.590000 ;
      RECT 966.500000 370.410000 999.500000 371.590000 ;
      RECT 957.500000 370.410000 958.500000 371.590000 ;
      RECT 916.500000 370.410000 949.500000 371.590000 ;
      RECT 907.500000 370.410000 908.500000 371.590000 ;
      RECT 866.500000 370.410000 899.500000 371.590000 ;
      RECT 857.500000 370.410000 858.500000 371.590000 ;
      RECT 816.500000 370.410000 849.500000 371.590000 ;
      RECT 807.500000 370.410000 808.500000 371.590000 ;
      RECT 766.500000 370.410000 799.500000 371.590000 ;
      RECT 757.500000 370.410000 758.500000 371.590000 ;
      RECT 716.500000 370.410000 749.500000 371.590000 ;
      RECT 707.500000 370.410000 708.500000 371.590000 ;
      RECT 666.500000 370.410000 699.500000 371.590000 ;
      RECT 657.500000 370.410000 658.500000 371.590000 ;
      RECT 616.500000 370.410000 649.500000 371.590000 ;
      RECT 607.500000 370.410000 608.500000 371.590000 ;
      RECT 566.500000 370.410000 599.500000 371.590000 ;
      RECT 557.500000 370.410000 558.500000 371.590000 ;
      RECT 516.500000 370.410000 549.500000 371.590000 ;
      RECT 507.500000 370.410000 508.500000 371.590000 ;
      RECT 466.500000 370.410000 499.500000 371.590000 ;
      RECT 457.500000 370.410000 458.500000 371.590000 ;
      RECT 416.500000 370.410000 449.500000 371.590000 ;
      RECT 407.500000 370.410000 408.500000 371.590000 ;
      RECT 366.500000 370.410000 399.500000 371.590000 ;
      RECT 357.500000 370.410000 358.500000 371.590000 ;
      RECT 316.500000 370.410000 349.500000 371.590000 ;
      RECT 307.500000 370.410000 308.500000 371.590000 ;
      RECT 266.500000 370.410000 299.500000 371.590000 ;
      RECT 257.500000 370.410000 258.500000 371.590000 ;
      RECT 216.500000 370.410000 249.500000 371.590000 ;
      RECT 207.500000 370.410000 208.500000 371.590000 ;
      RECT 166.500000 370.410000 199.500000 371.590000 ;
      RECT 157.500000 370.410000 158.500000 371.590000 ;
      RECT 116.500000 370.410000 149.500000 371.590000 ;
      RECT 107.500000 370.410000 108.500000 371.590000 ;
      RECT 66.500000 370.410000 99.500000 371.590000 ;
      RECT 57.500000 370.410000 58.500000 371.590000 ;
      RECT 29.500000 370.410000 49.500000 371.590000 ;
      RECT 15.500000 370.410000 16.500000 371.590000 ;
      RECT 1157.500000 369.590000 1170.500000 370.410000 ;
      RECT 1107.500000 369.590000 1149.500000 370.410000 ;
      RECT 1057.500000 369.590000 1099.500000 370.410000 ;
      RECT 1007.500000 369.590000 1049.500000 370.410000 ;
      RECT 957.500000 369.590000 999.500000 370.410000 ;
      RECT 907.500000 369.590000 949.500000 370.410000 ;
      RECT 857.500000 369.590000 899.500000 370.410000 ;
      RECT 807.500000 369.590000 849.500000 370.410000 ;
      RECT 757.500000 369.590000 799.500000 370.410000 ;
      RECT 707.500000 369.590000 749.500000 370.410000 ;
      RECT 657.500000 369.590000 699.500000 370.410000 ;
      RECT 607.500000 369.590000 649.500000 370.410000 ;
      RECT 557.500000 369.590000 599.500000 370.410000 ;
      RECT 507.500000 369.590000 549.500000 370.410000 ;
      RECT 407.500000 369.590000 449.500000 370.410000 ;
      RECT 357.500000 369.590000 399.500000 370.410000 ;
      RECT 307.500000 369.590000 349.500000 370.410000 ;
      RECT 257.500000 369.590000 299.500000 370.410000 ;
      RECT 207.500000 369.590000 249.500000 370.410000 ;
      RECT 157.500000 369.590000 199.500000 370.410000 ;
      RECT 107.500000 369.590000 149.500000 370.410000 ;
      RECT 57.500000 369.590000 99.500000 370.410000 ;
      RECT 15.500000 369.590000 49.500000 370.410000 ;
      RECT 1183.500000 368.410000 1186.000000 371.590000 ;
      RECT 1169.500000 368.410000 1170.500000 369.590000 ;
      RECT 1116.500000 368.410000 1149.500000 369.590000 ;
      RECT 1107.500000 368.410000 1108.500000 369.590000 ;
      RECT 1066.500000 368.410000 1099.500000 369.590000 ;
      RECT 1057.500000 368.410000 1058.500000 369.590000 ;
      RECT 1016.500000 368.410000 1049.500000 369.590000 ;
      RECT 1007.500000 368.410000 1008.500000 369.590000 ;
      RECT 966.500000 368.410000 999.500000 369.590000 ;
      RECT 957.500000 368.410000 958.500000 369.590000 ;
      RECT 916.500000 368.410000 949.500000 369.590000 ;
      RECT 907.500000 368.410000 908.500000 369.590000 ;
      RECT 866.500000 368.410000 899.500000 369.590000 ;
      RECT 857.500000 368.410000 858.500000 369.590000 ;
      RECT 816.500000 368.410000 849.500000 369.590000 ;
      RECT 807.500000 368.410000 808.500000 369.590000 ;
      RECT 766.500000 368.410000 799.500000 369.590000 ;
      RECT 757.500000 368.410000 758.500000 369.590000 ;
      RECT 716.500000 368.410000 749.500000 369.590000 ;
      RECT 707.500000 368.410000 708.500000 369.590000 ;
      RECT 666.500000 368.410000 699.500000 369.590000 ;
      RECT 657.500000 368.410000 658.500000 369.590000 ;
      RECT 616.500000 368.410000 649.500000 369.590000 ;
      RECT 607.500000 368.410000 608.500000 369.590000 ;
      RECT 566.500000 368.410000 599.500000 369.590000 ;
      RECT 557.500000 368.410000 558.500000 369.590000 ;
      RECT 516.500000 368.410000 549.500000 369.590000 ;
      RECT 507.500000 368.410000 508.500000 369.590000 ;
      RECT 457.500000 368.410000 499.500000 370.410000 ;
      RECT 416.500000 368.410000 449.500000 369.590000 ;
      RECT 407.500000 368.410000 408.500000 369.590000 ;
      RECT 366.500000 368.410000 399.500000 369.590000 ;
      RECT 357.500000 368.410000 358.500000 369.590000 ;
      RECT 316.500000 368.410000 349.500000 369.590000 ;
      RECT 307.500000 368.410000 308.500000 369.590000 ;
      RECT 266.500000 368.410000 299.500000 369.590000 ;
      RECT 257.500000 368.410000 258.500000 369.590000 ;
      RECT 216.500000 368.410000 249.500000 369.590000 ;
      RECT 207.500000 368.410000 208.500000 369.590000 ;
      RECT 166.500000 368.410000 199.500000 369.590000 ;
      RECT 157.500000 368.410000 158.500000 369.590000 ;
      RECT 116.500000 368.410000 149.500000 369.590000 ;
      RECT 107.500000 368.410000 108.500000 369.590000 ;
      RECT 66.500000 368.410000 99.500000 369.590000 ;
      RECT 57.500000 368.410000 58.500000 369.590000 ;
      RECT 29.500000 368.410000 49.500000 369.590000 ;
      RECT 15.500000 368.410000 16.500000 369.590000 ;
      RECT 0.000000 368.410000 2.500000 371.590000 ;
      RECT 1169.500000 367.590000 1186.000000 368.410000 ;
      RECT 1116.500000 367.590000 1156.500000 368.410000 ;
      RECT 1066.500000 367.590000 1108.500000 368.410000 ;
      RECT 1016.500000 367.590000 1058.500000 368.410000 ;
      RECT 966.500000 367.590000 1008.500000 368.410000 ;
      RECT 916.500000 367.590000 958.500000 368.410000 ;
      RECT 866.500000 367.590000 908.500000 368.410000 ;
      RECT 816.500000 367.590000 858.500000 368.410000 ;
      RECT 766.500000 367.590000 808.500000 368.410000 ;
      RECT 716.500000 367.590000 758.500000 368.410000 ;
      RECT 666.500000 367.590000 708.500000 368.410000 ;
      RECT 616.500000 367.590000 658.500000 368.410000 ;
      RECT 566.500000 367.590000 608.500000 368.410000 ;
      RECT 516.500000 367.590000 558.500000 368.410000 ;
      RECT 416.500000 367.590000 508.500000 368.410000 ;
      RECT 366.500000 367.590000 408.500000 368.410000 ;
      RECT 316.500000 367.590000 358.500000 368.410000 ;
      RECT 266.500000 367.590000 308.500000 368.410000 ;
      RECT 216.500000 367.590000 258.500000 368.410000 ;
      RECT 166.500000 367.590000 208.500000 368.410000 ;
      RECT 116.500000 367.590000 158.500000 368.410000 ;
      RECT 66.500000 367.590000 108.500000 368.410000 ;
      RECT 29.500000 367.590000 58.500000 368.410000 ;
      RECT 0.000000 367.590000 16.500000 368.410000 ;
      RECT 1169.500000 366.410000 1170.500000 367.590000 ;
      RECT 1116.500000 366.410000 1149.500000 367.590000 ;
      RECT 1107.500000 366.410000 1108.500000 367.590000 ;
      RECT 1066.500000 366.410000 1099.500000 367.590000 ;
      RECT 1057.500000 366.410000 1058.500000 367.590000 ;
      RECT 1016.500000 366.410000 1049.500000 367.590000 ;
      RECT 1007.500000 366.410000 1008.500000 367.590000 ;
      RECT 966.500000 366.410000 999.500000 367.590000 ;
      RECT 957.500000 366.410000 958.500000 367.590000 ;
      RECT 916.500000 366.410000 949.500000 367.590000 ;
      RECT 907.500000 366.410000 908.500000 367.590000 ;
      RECT 866.500000 366.410000 899.500000 367.590000 ;
      RECT 857.500000 366.410000 858.500000 367.590000 ;
      RECT 816.500000 366.410000 849.500000 367.590000 ;
      RECT 807.500000 366.410000 808.500000 367.590000 ;
      RECT 766.500000 366.410000 799.500000 367.590000 ;
      RECT 757.500000 366.410000 758.500000 367.590000 ;
      RECT 716.500000 366.410000 749.500000 367.590000 ;
      RECT 707.500000 366.410000 708.500000 367.590000 ;
      RECT 666.500000 366.410000 699.500000 367.590000 ;
      RECT 657.500000 366.410000 658.500000 367.590000 ;
      RECT 616.500000 366.410000 649.500000 367.590000 ;
      RECT 607.500000 366.410000 608.500000 367.590000 ;
      RECT 566.500000 366.410000 599.500000 367.590000 ;
      RECT 557.500000 366.410000 558.500000 367.590000 ;
      RECT 516.500000 366.410000 549.500000 367.590000 ;
      RECT 507.500000 366.410000 508.500000 367.590000 ;
      RECT 416.500000 366.410000 499.500000 367.590000 ;
      RECT 407.500000 366.410000 408.500000 367.590000 ;
      RECT 366.500000 366.410000 399.500000 367.590000 ;
      RECT 357.500000 366.410000 358.500000 367.590000 ;
      RECT 316.500000 366.410000 349.500000 367.590000 ;
      RECT 307.500000 366.410000 308.500000 367.590000 ;
      RECT 266.500000 366.410000 299.500000 367.590000 ;
      RECT 257.500000 366.410000 258.500000 367.590000 ;
      RECT 216.500000 366.410000 249.500000 367.590000 ;
      RECT 207.500000 366.410000 208.500000 367.590000 ;
      RECT 166.500000 366.410000 199.500000 367.590000 ;
      RECT 157.500000 366.410000 158.500000 367.590000 ;
      RECT 116.500000 366.410000 149.500000 367.590000 ;
      RECT 107.500000 366.410000 108.500000 367.590000 ;
      RECT 66.500000 366.410000 99.500000 367.590000 ;
      RECT 57.500000 366.410000 58.500000 367.590000 ;
      RECT 29.500000 366.410000 49.500000 367.590000 ;
      RECT 15.500000 366.410000 16.500000 367.590000 ;
      RECT 1157.500000 365.590000 1170.500000 366.410000 ;
      RECT 1107.500000 365.590000 1149.500000 366.410000 ;
      RECT 1057.500000 365.590000 1099.500000 366.410000 ;
      RECT 1007.500000 365.590000 1049.500000 366.410000 ;
      RECT 957.500000 365.590000 999.500000 366.410000 ;
      RECT 907.500000 365.590000 949.500000 366.410000 ;
      RECT 857.500000 365.590000 899.500000 366.410000 ;
      RECT 807.500000 365.590000 849.500000 366.410000 ;
      RECT 757.500000 365.590000 799.500000 366.410000 ;
      RECT 707.500000 365.590000 749.500000 366.410000 ;
      RECT 657.500000 365.590000 699.500000 366.410000 ;
      RECT 607.500000 365.590000 649.500000 366.410000 ;
      RECT 557.500000 365.590000 599.500000 366.410000 ;
      RECT 507.500000 365.590000 549.500000 366.410000 ;
      RECT 407.500000 365.590000 499.500000 366.410000 ;
      RECT 357.500000 365.590000 399.500000 366.410000 ;
      RECT 307.500000 365.590000 349.500000 366.410000 ;
      RECT 257.500000 365.590000 299.500000 366.410000 ;
      RECT 207.500000 365.590000 249.500000 366.410000 ;
      RECT 157.500000 365.590000 199.500000 366.410000 ;
      RECT 107.500000 365.590000 149.500000 366.410000 ;
      RECT 57.500000 365.590000 99.500000 366.410000 ;
      RECT 15.500000 365.590000 49.500000 366.410000 ;
      RECT 1183.500000 364.410000 1186.000000 367.590000 ;
      RECT 1169.500000 364.410000 1170.500000 365.590000 ;
      RECT 1116.500000 364.410000 1149.500000 365.590000 ;
      RECT 1107.500000 364.410000 1108.500000 365.590000 ;
      RECT 1066.500000 364.410000 1099.500000 365.590000 ;
      RECT 1057.500000 364.410000 1058.500000 365.590000 ;
      RECT 1016.500000 364.410000 1049.500000 365.590000 ;
      RECT 1007.500000 364.410000 1008.500000 365.590000 ;
      RECT 966.500000 364.410000 999.500000 365.590000 ;
      RECT 957.500000 364.410000 958.500000 365.590000 ;
      RECT 916.500000 364.410000 949.500000 365.590000 ;
      RECT 907.500000 364.410000 908.500000 365.590000 ;
      RECT 866.500000 364.410000 899.500000 365.590000 ;
      RECT 857.500000 364.410000 858.500000 365.590000 ;
      RECT 816.500000 364.410000 849.500000 365.590000 ;
      RECT 807.500000 364.410000 808.500000 365.590000 ;
      RECT 766.500000 364.410000 799.500000 365.590000 ;
      RECT 757.500000 364.410000 758.500000 365.590000 ;
      RECT 716.500000 364.410000 749.500000 365.590000 ;
      RECT 707.500000 364.410000 708.500000 365.590000 ;
      RECT 666.500000 364.410000 699.500000 365.590000 ;
      RECT 657.500000 364.410000 658.500000 365.590000 ;
      RECT 616.500000 364.410000 649.500000 365.590000 ;
      RECT 607.500000 364.410000 608.500000 365.590000 ;
      RECT 566.500000 364.410000 599.500000 365.590000 ;
      RECT 557.500000 364.410000 558.500000 365.590000 ;
      RECT 516.500000 364.410000 549.500000 365.590000 ;
      RECT 507.500000 364.410000 508.500000 365.590000 ;
      RECT 416.500000 364.410000 499.500000 365.590000 ;
      RECT 407.500000 364.410000 408.500000 365.590000 ;
      RECT 366.500000 364.410000 399.500000 365.590000 ;
      RECT 357.500000 364.410000 358.500000 365.590000 ;
      RECT 316.500000 364.410000 349.500000 365.590000 ;
      RECT 307.500000 364.410000 308.500000 365.590000 ;
      RECT 266.500000 364.410000 299.500000 365.590000 ;
      RECT 257.500000 364.410000 258.500000 365.590000 ;
      RECT 216.500000 364.410000 249.500000 365.590000 ;
      RECT 207.500000 364.410000 208.500000 365.590000 ;
      RECT 166.500000 364.410000 199.500000 365.590000 ;
      RECT 157.500000 364.410000 158.500000 365.590000 ;
      RECT 116.500000 364.410000 149.500000 365.590000 ;
      RECT 107.500000 364.410000 108.500000 365.590000 ;
      RECT 66.500000 364.410000 99.500000 365.590000 ;
      RECT 57.500000 364.410000 58.500000 365.590000 ;
      RECT 29.500000 364.410000 49.500000 365.590000 ;
      RECT 15.500000 364.410000 16.500000 365.590000 ;
      RECT 0.000000 364.410000 2.500000 367.590000 ;
      RECT 1169.500000 363.590000 1186.000000 364.410000 ;
      RECT 1116.500000 363.590000 1156.500000 364.410000 ;
      RECT 1066.500000 363.590000 1108.500000 364.410000 ;
      RECT 1016.500000 363.590000 1058.500000 364.410000 ;
      RECT 966.500000 363.590000 1008.500000 364.410000 ;
      RECT 916.500000 363.590000 958.500000 364.410000 ;
      RECT 866.500000 363.590000 908.500000 364.410000 ;
      RECT 816.500000 363.590000 858.500000 364.410000 ;
      RECT 766.500000 363.590000 808.500000 364.410000 ;
      RECT 716.500000 363.590000 758.500000 364.410000 ;
      RECT 666.500000 363.590000 708.500000 364.410000 ;
      RECT 616.500000 363.590000 658.500000 364.410000 ;
      RECT 566.500000 363.590000 608.500000 364.410000 ;
      RECT 516.500000 363.590000 558.500000 364.410000 ;
      RECT 416.500000 363.590000 508.500000 364.410000 ;
      RECT 366.500000 363.590000 408.500000 364.410000 ;
      RECT 316.500000 363.590000 358.500000 364.410000 ;
      RECT 266.500000 363.590000 308.500000 364.410000 ;
      RECT 216.500000 363.590000 258.500000 364.410000 ;
      RECT 166.500000 363.590000 208.500000 364.410000 ;
      RECT 116.500000 363.590000 158.500000 364.410000 ;
      RECT 66.500000 363.590000 108.500000 364.410000 ;
      RECT 29.500000 363.590000 58.500000 364.410000 ;
      RECT 0.000000 363.590000 16.500000 364.410000 ;
      RECT 1169.500000 362.410000 1170.500000 363.590000 ;
      RECT 1116.500000 362.410000 1149.500000 363.590000 ;
      RECT 1107.500000 362.410000 1108.500000 363.590000 ;
      RECT 1066.500000 362.410000 1099.500000 363.590000 ;
      RECT 1057.500000 362.410000 1058.500000 363.590000 ;
      RECT 1016.500000 362.410000 1049.500000 363.590000 ;
      RECT 1007.500000 362.410000 1008.500000 363.590000 ;
      RECT 966.500000 362.410000 999.500000 363.590000 ;
      RECT 957.500000 362.410000 958.500000 363.590000 ;
      RECT 916.500000 362.410000 949.500000 363.590000 ;
      RECT 907.500000 362.410000 908.500000 363.590000 ;
      RECT 866.500000 362.410000 899.500000 363.590000 ;
      RECT 857.500000 362.410000 858.500000 363.590000 ;
      RECT 816.500000 362.410000 849.500000 363.590000 ;
      RECT 807.500000 362.410000 808.500000 363.590000 ;
      RECT 766.500000 362.410000 799.500000 363.590000 ;
      RECT 757.500000 362.410000 758.500000 363.590000 ;
      RECT 716.500000 362.410000 749.500000 363.590000 ;
      RECT 707.500000 362.410000 708.500000 363.590000 ;
      RECT 666.500000 362.410000 699.500000 363.590000 ;
      RECT 657.500000 362.410000 658.500000 363.590000 ;
      RECT 616.500000 362.410000 649.500000 363.590000 ;
      RECT 607.500000 362.410000 608.500000 363.590000 ;
      RECT 566.500000 362.410000 599.500000 363.590000 ;
      RECT 557.500000 362.410000 558.500000 363.590000 ;
      RECT 516.500000 362.410000 549.500000 363.590000 ;
      RECT 507.500000 362.410000 508.500000 363.590000 ;
      RECT 416.500000 362.410000 499.500000 363.590000 ;
      RECT 407.500000 362.410000 408.500000 363.590000 ;
      RECT 366.500000 362.410000 399.500000 363.590000 ;
      RECT 357.500000 362.410000 358.500000 363.590000 ;
      RECT 316.500000 362.410000 349.500000 363.590000 ;
      RECT 307.500000 362.410000 308.500000 363.590000 ;
      RECT 266.500000 362.410000 299.500000 363.590000 ;
      RECT 257.500000 362.410000 258.500000 363.590000 ;
      RECT 216.500000 362.410000 249.500000 363.590000 ;
      RECT 207.500000 362.410000 208.500000 363.590000 ;
      RECT 166.500000 362.410000 199.500000 363.590000 ;
      RECT 157.500000 362.410000 158.500000 363.590000 ;
      RECT 116.500000 362.410000 149.500000 363.590000 ;
      RECT 107.500000 362.410000 108.500000 363.590000 ;
      RECT 66.500000 362.410000 99.500000 363.590000 ;
      RECT 57.500000 362.410000 58.500000 363.590000 ;
      RECT 29.500000 362.410000 49.500000 363.590000 ;
      RECT 15.500000 362.410000 16.500000 363.590000 ;
      RECT 1157.500000 361.590000 1170.500000 362.410000 ;
      RECT 1107.500000 361.590000 1149.500000 362.410000 ;
      RECT 1057.500000 361.590000 1099.500000 362.410000 ;
      RECT 1007.500000 361.590000 1049.500000 362.410000 ;
      RECT 957.500000 361.590000 999.500000 362.410000 ;
      RECT 907.500000 361.590000 949.500000 362.410000 ;
      RECT 857.500000 361.590000 899.500000 362.410000 ;
      RECT 807.500000 361.590000 849.500000 362.410000 ;
      RECT 757.500000 361.590000 799.500000 362.410000 ;
      RECT 707.500000 361.590000 749.500000 362.410000 ;
      RECT 657.500000 361.590000 699.500000 362.410000 ;
      RECT 607.500000 361.590000 649.500000 362.410000 ;
      RECT 557.500000 361.590000 599.500000 362.410000 ;
      RECT 507.500000 361.590000 549.500000 362.410000 ;
      RECT 407.500000 361.590000 499.500000 362.410000 ;
      RECT 357.500000 361.590000 399.500000 362.410000 ;
      RECT 307.500000 361.590000 349.500000 362.410000 ;
      RECT 257.500000 361.590000 299.500000 362.410000 ;
      RECT 207.500000 361.590000 249.500000 362.410000 ;
      RECT 157.500000 361.590000 199.500000 362.410000 ;
      RECT 107.500000 361.590000 149.500000 362.410000 ;
      RECT 15.500000 361.590000 49.500000 362.410000 ;
      RECT 1183.500000 360.410000 1186.000000 363.590000 ;
      RECT 1169.500000 360.410000 1170.500000 361.590000 ;
      RECT 1116.500000 360.410000 1149.500000 361.590000 ;
      RECT 1107.500000 360.410000 1108.500000 361.590000 ;
      RECT 1066.500000 360.410000 1099.500000 361.590000 ;
      RECT 1057.500000 360.410000 1058.500000 361.590000 ;
      RECT 1016.500000 360.410000 1049.500000 361.590000 ;
      RECT 1007.500000 360.410000 1008.500000 361.590000 ;
      RECT 966.500000 360.410000 999.500000 361.590000 ;
      RECT 957.500000 360.410000 958.500000 361.590000 ;
      RECT 916.500000 360.410000 949.500000 361.590000 ;
      RECT 907.500000 360.410000 908.500000 361.590000 ;
      RECT 866.500000 360.410000 899.500000 361.590000 ;
      RECT 857.500000 360.410000 858.500000 361.590000 ;
      RECT 816.500000 360.410000 849.500000 361.590000 ;
      RECT 807.500000 360.410000 808.500000 361.590000 ;
      RECT 766.500000 360.410000 799.500000 361.590000 ;
      RECT 757.500000 360.410000 758.500000 361.590000 ;
      RECT 716.500000 360.410000 749.500000 361.590000 ;
      RECT 707.500000 360.410000 708.500000 361.590000 ;
      RECT 666.500000 360.410000 699.500000 361.590000 ;
      RECT 657.500000 360.410000 658.500000 361.590000 ;
      RECT 616.500000 360.410000 649.500000 361.590000 ;
      RECT 607.500000 360.410000 608.500000 361.590000 ;
      RECT 566.500000 360.410000 599.500000 361.590000 ;
      RECT 557.500000 360.410000 558.500000 361.590000 ;
      RECT 516.500000 360.410000 549.500000 361.590000 ;
      RECT 507.500000 360.410000 508.500000 361.590000 ;
      RECT 416.500000 360.410000 499.500000 361.590000 ;
      RECT 407.500000 360.410000 408.500000 361.590000 ;
      RECT 366.500000 360.410000 399.500000 361.590000 ;
      RECT 357.500000 360.410000 358.500000 361.590000 ;
      RECT 316.500000 360.410000 349.500000 361.590000 ;
      RECT 307.500000 360.410000 308.500000 361.590000 ;
      RECT 266.500000 360.410000 299.500000 361.590000 ;
      RECT 257.500000 360.410000 258.500000 361.590000 ;
      RECT 216.500000 360.410000 249.500000 361.590000 ;
      RECT 207.500000 360.410000 208.500000 361.590000 ;
      RECT 166.500000 360.410000 199.500000 361.590000 ;
      RECT 157.500000 360.410000 158.500000 361.590000 ;
      RECT 116.500000 360.410000 149.500000 361.590000 ;
      RECT 107.500000 360.410000 108.500000 361.590000 ;
      RECT 57.500000 360.410000 99.500000 362.410000 ;
      RECT 29.500000 360.410000 49.500000 361.590000 ;
      RECT 15.500000 360.410000 16.500000 361.590000 ;
      RECT 0.000000 360.410000 2.500000 363.590000 ;
      RECT 1169.500000 359.590000 1186.000000 360.410000 ;
      RECT 1116.500000 359.590000 1156.500000 360.410000 ;
      RECT 1066.500000 359.590000 1108.500000 360.410000 ;
      RECT 1016.500000 359.590000 1058.500000 360.410000 ;
      RECT 966.500000 359.590000 1008.500000 360.410000 ;
      RECT 916.500000 359.590000 958.500000 360.410000 ;
      RECT 866.500000 359.590000 908.500000 360.410000 ;
      RECT 816.500000 359.590000 858.500000 360.410000 ;
      RECT 766.500000 359.590000 808.500000 360.410000 ;
      RECT 716.500000 359.590000 758.500000 360.410000 ;
      RECT 666.500000 359.590000 708.500000 360.410000 ;
      RECT 616.500000 359.590000 658.500000 360.410000 ;
      RECT 566.500000 359.590000 608.500000 360.410000 ;
      RECT 516.500000 359.590000 558.500000 360.410000 ;
      RECT 416.500000 359.590000 508.500000 360.410000 ;
      RECT 366.500000 359.590000 408.500000 360.410000 ;
      RECT 316.500000 359.590000 358.500000 360.410000 ;
      RECT 266.500000 359.590000 308.500000 360.410000 ;
      RECT 216.500000 359.590000 258.500000 360.410000 ;
      RECT 166.500000 359.590000 208.500000 360.410000 ;
      RECT 116.500000 359.590000 158.500000 360.410000 ;
      RECT 29.500000 359.590000 108.500000 360.410000 ;
      RECT 0.000000 359.590000 16.500000 360.410000 ;
      RECT 1169.500000 358.410000 1170.500000 359.590000 ;
      RECT 1116.500000 358.410000 1149.500000 359.590000 ;
      RECT 1107.500000 358.410000 1108.500000 359.590000 ;
      RECT 1066.500000 358.410000 1099.500000 359.590000 ;
      RECT 1057.500000 358.410000 1058.500000 359.590000 ;
      RECT 1016.500000 358.410000 1049.500000 359.590000 ;
      RECT 1007.500000 358.410000 1008.500000 359.590000 ;
      RECT 966.500000 358.410000 999.500000 359.590000 ;
      RECT 957.500000 358.410000 958.500000 359.590000 ;
      RECT 916.500000 358.410000 949.500000 359.590000 ;
      RECT 907.500000 358.410000 908.500000 359.590000 ;
      RECT 866.500000 358.410000 899.500000 359.590000 ;
      RECT 857.500000 358.410000 858.500000 359.590000 ;
      RECT 816.500000 358.410000 849.500000 359.590000 ;
      RECT 807.500000 358.410000 808.500000 359.590000 ;
      RECT 766.500000 358.410000 799.500000 359.590000 ;
      RECT 757.500000 358.410000 758.500000 359.590000 ;
      RECT 716.500000 358.410000 749.500000 359.590000 ;
      RECT 707.500000 358.410000 708.500000 359.590000 ;
      RECT 666.500000 358.410000 699.500000 359.590000 ;
      RECT 657.500000 358.410000 658.500000 359.590000 ;
      RECT 616.500000 358.410000 649.500000 359.590000 ;
      RECT 607.500000 358.410000 608.500000 359.590000 ;
      RECT 566.500000 358.410000 599.500000 359.590000 ;
      RECT 557.500000 358.410000 558.500000 359.590000 ;
      RECT 516.500000 358.410000 549.500000 359.590000 ;
      RECT 507.500000 358.410000 508.500000 359.590000 ;
      RECT 416.500000 358.410000 499.500000 359.590000 ;
      RECT 407.500000 358.410000 408.500000 359.590000 ;
      RECT 366.500000 358.410000 399.500000 359.590000 ;
      RECT 357.500000 358.410000 358.500000 359.590000 ;
      RECT 316.500000 358.410000 349.500000 359.590000 ;
      RECT 307.500000 358.410000 308.500000 359.590000 ;
      RECT 266.500000 358.410000 299.500000 359.590000 ;
      RECT 257.500000 358.410000 258.500000 359.590000 ;
      RECT 216.500000 358.410000 249.500000 359.590000 ;
      RECT 207.500000 358.410000 208.500000 359.590000 ;
      RECT 166.500000 358.410000 199.500000 359.590000 ;
      RECT 157.500000 358.410000 158.500000 359.590000 ;
      RECT 116.500000 358.410000 149.500000 359.590000 ;
      RECT 107.500000 358.410000 108.500000 359.590000 ;
      RECT 29.500000 358.410000 99.500000 359.590000 ;
      RECT 15.500000 358.410000 16.500000 359.590000 ;
      RECT 1157.500000 357.590000 1170.500000 358.410000 ;
      RECT 1107.500000 357.590000 1149.500000 358.410000 ;
      RECT 1057.500000 357.590000 1099.500000 358.410000 ;
      RECT 1007.500000 357.590000 1049.500000 358.410000 ;
      RECT 957.500000 357.590000 999.500000 358.410000 ;
      RECT 907.500000 357.590000 949.500000 358.410000 ;
      RECT 857.500000 357.590000 899.500000 358.410000 ;
      RECT 807.500000 357.590000 849.500000 358.410000 ;
      RECT 757.500000 357.590000 799.500000 358.410000 ;
      RECT 707.500000 357.590000 749.500000 358.410000 ;
      RECT 657.500000 357.590000 699.500000 358.410000 ;
      RECT 607.500000 357.590000 649.500000 358.410000 ;
      RECT 557.500000 357.590000 599.500000 358.410000 ;
      RECT 507.500000 357.590000 549.500000 358.410000 ;
      RECT 407.500000 357.590000 499.500000 358.410000 ;
      RECT 357.500000 357.590000 399.500000 358.410000 ;
      RECT 307.500000 357.590000 349.500000 358.410000 ;
      RECT 257.500000 357.590000 299.500000 358.410000 ;
      RECT 207.500000 357.590000 249.500000 358.410000 ;
      RECT 157.500000 357.590000 199.500000 358.410000 ;
      RECT 107.500000 357.590000 149.500000 358.410000 ;
      RECT 15.500000 357.590000 99.500000 358.410000 ;
      RECT 1183.500000 356.410000 1186.000000 359.590000 ;
      RECT 1169.500000 356.410000 1170.500000 357.590000 ;
      RECT 1116.500000 356.410000 1149.500000 357.590000 ;
      RECT 1107.500000 356.410000 1108.500000 357.590000 ;
      RECT 1066.500000 356.410000 1099.500000 357.590000 ;
      RECT 1057.500000 356.410000 1058.500000 357.590000 ;
      RECT 1016.500000 356.410000 1049.500000 357.590000 ;
      RECT 1007.500000 356.410000 1008.500000 357.590000 ;
      RECT 966.500000 356.410000 999.500000 357.590000 ;
      RECT 957.500000 356.410000 958.500000 357.590000 ;
      RECT 916.500000 356.410000 949.500000 357.590000 ;
      RECT 907.500000 356.410000 908.500000 357.590000 ;
      RECT 866.500000 356.410000 899.500000 357.590000 ;
      RECT 857.500000 356.410000 858.500000 357.590000 ;
      RECT 816.500000 356.410000 849.500000 357.590000 ;
      RECT 807.500000 356.410000 808.500000 357.590000 ;
      RECT 766.500000 356.410000 799.500000 357.590000 ;
      RECT 757.500000 356.410000 758.500000 357.590000 ;
      RECT 716.500000 356.410000 749.500000 357.590000 ;
      RECT 707.500000 356.410000 708.500000 357.590000 ;
      RECT 666.500000 356.410000 699.500000 357.590000 ;
      RECT 657.500000 356.410000 658.500000 357.590000 ;
      RECT 616.500000 356.410000 649.500000 357.590000 ;
      RECT 607.500000 356.410000 608.500000 357.590000 ;
      RECT 566.500000 356.410000 599.500000 357.590000 ;
      RECT 557.500000 356.410000 558.500000 357.590000 ;
      RECT 516.500000 356.410000 549.500000 357.590000 ;
      RECT 507.500000 356.410000 508.500000 357.590000 ;
      RECT 416.500000 356.410000 499.500000 357.590000 ;
      RECT 407.500000 356.410000 408.500000 357.590000 ;
      RECT 366.500000 356.410000 399.500000 357.590000 ;
      RECT 357.500000 356.410000 358.500000 357.590000 ;
      RECT 316.500000 356.410000 349.500000 357.590000 ;
      RECT 307.500000 356.410000 308.500000 357.590000 ;
      RECT 266.500000 356.410000 299.500000 357.590000 ;
      RECT 257.500000 356.410000 258.500000 357.590000 ;
      RECT 216.500000 356.410000 249.500000 357.590000 ;
      RECT 207.500000 356.410000 208.500000 357.590000 ;
      RECT 166.500000 356.410000 199.500000 357.590000 ;
      RECT 157.500000 356.410000 158.500000 357.590000 ;
      RECT 116.500000 356.410000 149.500000 357.590000 ;
      RECT 107.500000 356.410000 108.500000 357.590000 ;
      RECT 29.500000 356.410000 99.500000 357.590000 ;
      RECT 15.500000 356.410000 16.500000 357.590000 ;
      RECT 0.000000 356.410000 2.500000 359.590000 ;
      RECT 1169.500000 355.590000 1186.000000 356.410000 ;
      RECT 1116.500000 355.590000 1156.500000 356.410000 ;
      RECT 1066.500000 355.590000 1108.500000 356.410000 ;
      RECT 1016.500000 355.590000 1058.500000 356.410000 ;
      RECT 966.500000 355.590000 1008.500000 356.410000 ;
      RECT 916.500000 355.590000 958.500000 356.410000 ;
      RECT 866.500000 355.590000 908.500000 356.410000 ;
      RECT 816.500000 355.590000 858.500000 356.410000 ;
      RECT 766.500000 355.590000 808.500000 356.410000 ;
      RECT 716.500000 355.590000 758.500000 356.410000 ;
      RECT 666.500000 355.590000 708.500000 356.410000 ;
      RECT 616.500000 355.590000 658.500000 356.410000 ;
      RECT 566.500000 355.590000 608.500000 356.410000 ;
      RECT 516.500000 355.590000 558.500000 356.410000 ;
      RECT 416.500000 355.590000 508.500000 356.410000 ;
      RECT 366.500000 355.590000 408.500000 356.410000 ;
      RECT 316.500000 355.590000 358.500000 356.410000 ;
      RECT 266.500000 355.590000 308.500000 356.410000 ;
      RECT 216.500000 355.590000 258.500000 356.410000 ;
      RECT 166.500000 355.590000 208.500000 356.410000 ;
      RECT 116.500000 355.590000 158.500000 356.410000 ;
      RECT 29.500000 355.590000 108.500000 356.410000 ;
      RECT 0.000000 355.590000 16.500000 356.410000 ;
      RECT 1169.500000 354.410000 1170.500000 355.590000 ;
      RECT 1116.500000 354.410000 1149.500000 355.590000 ;
      RECT 1107.500000 354.410000 1108.500000 355.590000 ;
      RECT 1066.500000 354.410000 1099.500000 355.590000 ;
      RECT 1057.500000 354.410000 1058.500000 355.590000 ;
      RECT 1016.500000 354.410000 1049.500000 355.590000 ;
      RECT 1007.500000 354.410000 1008.500000 355.590000 ;
      RECT 966.500000 354.410000 999.500000 355.590000 ;
      RECT 957.500000 354.410000 958.500000 355.590000 ;
      RECT 916.500000 354.410000 949.500000 355.590000 ;
      RECT 907.500000 354.410000 908.500000 355.590000 ;
      RECT 866.500000 354.410000 899.500000 355.590000 ;
      RECT 857.500000 354.410000 858.500000 355.590000 ;
      RECT 816.500000 354.410000 849.500000 355.590000 ;
      RECT 807.500000 354.410000 808.500000 355.590000 ;
      RECT 766.500000 354.410000 799.500000 355.590000 ;
      RECT 757.500000 354.410000 758.500000 355.590000 ;
      RECT 716.500000 354.410000 749.500000 355.590000 ;
      RECT 707.500000 354.410000 708.500000 355.590000 ;
      RECT 666.500000 354.410000 699.500000 355.590000 ;
      RECT 657.500000 354.410000 658.500000 355.590000 ;
      RECT 616.500000 354.410000 649.500000 355.590000 ;
      RECT 607.500000 354.410000 608.500000 355.590000 ;
      RECT 566.500000 354.410000 599.500000 355.590000 ;
      RECT 557.500000 354.410000 558.500000 355.590000 ;
      RECT 516.500000 354.410000 549.500000 355.590000 ;
      RECT 507.500000 354.410000 508.500000 355.590000 ;
      RECT 416.500000 354.410000 499.500000 355.590000 ;
      RECT 407.500000 354.410000 408.500000 355.590000 ;
      RECT 366.500000 354.410000 399.500000 355.590000 ;
      RECT 357.500000 354.410000 358.500000 355.590000 ;
      RECT 316.500000 354.410000 349.500000 355.590000 ;
      RECT 307.500000 354.410000 308.500000 355.590000 ;
      RECT 266.500000 354.410000 299.500000 355.590000 ;
      RECT 257.500000 354.410000 258.500000 355.590000 ;
      RECT 216.500000 354.410000 249.500000 355.590000 ;
      RECT 207.500000 354.410000 208.500000 355.590000 ;
      RECT 166.500000 354.410000 199.500000 355.590000 ;
      RECT 157.500000 354.410000 158.500000 355.590000 ;
      RECT 116.500000 354.410000 149.500000 355.590000 ;
      RECT 107.500000 354.410000 108.500000 355.590000 ;
      RECT 29.500000 354.410000 99.500000 355.590000 ;
      RECT 15.500000 354.410000 16.500000 355.590000 ;
      RECT 1157.500000 353.590000 1170.500000 354.410000 ;
      RECT 1107.500000 353.590000 1149.500000 354.410000 ;
      RECT 1057.500000 353.590000 1099.500000 354.410000 ;
      RECT 1007.500000 353.590000 1049.500000 354.410000 ;
      RECT 957.500000 353.590000 999.500000 354.410000 ;
      RECT 907.500000 353.590000 949.500000 354.410000 ;
      RECT 857.500000 353.590000 899.500000 354.410000 ;
      RECT 807.500000 353.590000 849.500000 354.410000 ;
      RECT 757.500000 353.590000 799.500000 354.410000 ;
      RECT 707.500000 353.590000 749.500000 354.410000 ;
      RECT 657.500000 353.590000 699.500000 354.410000 ;
      RECT 607.500000 353.590000 649.500000 354.410000 ;
      RECT 557.500000 353.590000 599.500000 354.410000 ;
      RECT 507.500000 353.590000 549.500000 354.410000 ;
      RECT 407.500000 353.590000 499.500000 354.410000 ;
      RECT 357.500000 353.590000 399.500000 354.410000 ;
      RECT 307.500000 353.590000 349.500000 354.410000 ;
      RECT 257.500000 353.590000 299.500000 354.410000 ;
      RECT 207.500000 353.590000 249.500000 354.410000 ;
      RECT 157.500000 353.590000 199.500000 354.410000 ;
      RECT 107.500000 353.590000 149.500000 354.410000 ;
      RECT 15.500000 353.590000 99.500000 354.410000 ;
      RECT 1183.500000 352.410000 1186.000000 355.590000 ;
      RECT 1169.500000 352.410000 1170.500000 353.590000 ;
      RECT 1116.500000 352.410000 1149.500000 353.590000 ;
      RECT 1107.500000 352.410000 1108.500000 353.590000 ;
      RECT 1066.500000 352.410000 1099.500000 353.590000 ;
      RECT 1057.500000 352.410000 1058.500000 353.590000 ;
      RECT 1016.500000 352.410000 1049.500000 353.590000 ;
      RECT 1007.500000 352.410000 1008.500000 353.590000 ;
      RECT 966.500000 352.410000 999.500000 353.590000 ;
      RECT 957.500000 352.410000 958.500000 353.590000 ;
      RECT 916.500000 352.410000 949.500000 353.590000 ;
      RECT 907.500000 352.410000 908.500000 353.590000 ;
      RECT 866.500000 352.410000 899.500000 353.590000 ;
      RECT 857.500000 352.410000 858.500000 353.590000 ;
      RECT 816.500000 352.410000 849.500000 353.590000 ;
      RECT 807.500000 352.410000 808.500000 353.590000 ;
      RECT 766.500000 352.410000 799.500000 353.590000 ;
      RECT 757.500000 352.410000 758.500000 353.590000 ;
      RECT 716.500000 352.410000 749.500000 353.590000 ;
      RECT 707.500000 352.410000 708.500000 353.590000 ;
      RECT 666.500000 352.410000 699.500000 353.590000 ;
      RECT 657.500000 352.410000 658.500000 353.590000 ;
      RECT 616.500000 352.410000 649.500000 353.590000 ;
      RECT 607.500000 352.410000 608.500000 353.590000 ;
      RECT 566.500000 352.410000 599.500000 353.590000 ;
      RECT 557.500000 352.410000 558.500000 353.590000 ;
      RECT 516.500000 352.410000 549.500000 353.590000 ;
      RECT 507.500000 352.410000 508.500000 353.590000 ;
      RECT 416.500000 352.410000 499.500000 353.590000 ;
      RECT 407.500000 352.410000 408.500000 353.590000 ;
      RECT 366.500000 352.410000 399.500000 353.590000 ;
      RECT 357.500000 352.410000 358.500000 353.590000 ;
      RECT 316.500000 352.410000 349.500000 353.590000 ;
      RECT 307.500000 352.410000 308.500000 353.590000 ;
      RECT 266.500000 352.410000 299.500000 353.590000 ;
      RECT 257.500000 352.410000 258.500000 353.590000 ;
      RECT 216.500000 352.410000 249.500000 353.590000 ;
      RECT 207.500000 352.410000 208.500000 353.590000 ;
      RECT 166.500000 352.410000 199.500000 353.590000 ;
      RECT 157.500000 352.410000 158.500000 353.590000 ;
      RECT 116.500000 352.410000 149.500000 353.590000 ;
      RECT 107.500000 352.410000 108.500000 353.590000 ;
      RECT 29.500000 352.410000 99.500000 353.590000 ;
      RECT 15.500000 352.410000 16.500000 353.590000 ;
      RECT 0.000000 352.410000 2.500000 355.590000 ;
      RECT 1169.500000 351.590000 1186.000000 352.410000 ;
      RECT 1116.500000 351.590000 1156.500000 352.410000 ;
      RECT 1066.500000 351.590000 1108.500000 352.410000 ;
      RECT 1016.500000 351.590000 1058.500000 352.410000 ;
      RECT 966.500000 351.590000 1008.500000 352.410000 ;
      RECT 916.500000 351.590000 958.500000 352.410000 ;
      RECT 866.500000 351.590000 908.500000 352.410000 ;
      RECT 816.500000 351.590000 858.500000 352.410000 ;
      RECT 766.500000 351.590000 808.500000 352.410000 ;
      RECT 716.500000 351.590000 758.500000 352.410000 ;
      RECT 666.500000 351.590000 708.500000 352.410000 ;
      RECT 616.500000 351.590000 658.500000 352.410000 ;
      RECT 566.500000 351.590000 608.500000 352.410000 ;
      RECT 516.500000 351.590000 558.500000 352.410000 ;
      RECT 416.500000 351.590000 508.500000 352.410000 ;
      RECT 366.500000 351.590000 408.500000 352.410000 ;
      RECT 316.500000 351.590000 358.500000 352.410000 ;
      RECT 266.500000 351.590000 308.500000 352.410000 ;
      RECT 216.500000 351.590000 258.500000 352.410000 ;
      RECT 166.500000 351.590000 208.500000 352.410000 ;
      RECT 116.500000 351.590000 158.500000 352.410000 ;
      RECT 29.500000 351.590000 108.500000 352.410000 ;
      RECT 0.000000 351.590000 16.500000 352.410000 ;
      RECT 1169.500000 350.410000 1170.500000 351.590000 ;
      RECT 1116.500000 350.410000 1149.500000 351.590000 ;
      RECT 1107.500000 350.410000 1108.500000 351.590000 ;
      RECT 1066.500000 350.410000 1099.500000 351.590000 ;
      RECT 1057.500000 350.410000 1058.500000 351.590000 ;
      RECT 1016.500000 350.410000 1049.500000 351.590000 ;
      RECT 1007.500000 350.410000 1008.500000 351.590000 ;
      RECT 966.500000 350.410000 999.500000 351.590000 ;
      RECT 957.500000 350.410000 958.500000 351.590000 ;
      RECT 916.500000 350.410000 949.500000 351.590000 ;
      RECT 907.500000 350.410000 908.500000 351.590000 ;
      RECT 866.500000 350.410000 899.500000 351.590000 ;
      RECT 857.500000 350.410000 858.500000 351.590000 ;
      RECT 816.500000 350.410000 849.500000 351.590000 ;
      RECT 807.500000 350.410000 808.500000 351.590000 ;
      RECT 766.500000 350.410000 799.500000 351.590000 ;
      RECT 757.500000 350.410000 758.500000 351.590000 ;
      RECT 716.500000 350.410000 749.500000 351.590000 ;
      RECT 707.500000 350.410000 708.500000 351.590000 ;
      RECT 666.500000 350.410000 699.500000 351.590000 ;
      RECT 657.500000 350.410000 658.500000 351.590000 ;
      RECT 616.500000 350.410000 649.500000 351.590000 ;
      RECT 607.500000 350.410000 608.500000 351.590000 ;
      RECT 566.500000 350.410000 599.500000 351.590000 ;
      RECT 557.500000 350.410000 558.500000 351.590000 ;
      RECT 516.500000 350.410000 549.500000 351.590000 ;
      RECT 507.500000 350.410000 508.500000 351.590000 ;
      RECT 416.500000 350.410000 499.500000 351.590000 ;
      RECT 407.500000 350.410000 408.500000 351.590000 ;
      RECT 366.500000 350.410000 399.500000 351.590000 ;
      RECT 357.500000 350.410000 358.500000 351.590000 ;
      RECT 316.500000 350.410000 349.500000 351.590000 ;
      RECT 307.500000 350.410000 308.500000 351.590000 ;
      RECT 266.500000 350.410000 299.500000 351.590000 ;
      RECT 257.500000 350.410000 258.500000 351.590000 ;
      RECT 216.500000 350.410000 249.500000 351.590000 ;
      RECT 207.500000 350.410000 208.500000 351.590000 ;
      RECT 166.500000 350.410000 199.500000 351.590000 ;
      RECT 157.500000 350.410000 158.500000 351.590000 ;
      RECT 116.500000 350.410000 149.500000 351.590000 ;
      RECT 107.500000 350.410000 108.500000 351.590000 ;
      RECT 29.500000 350.410000 99.500000 351.590000 ;
      RECT 15.500000 350.410000 16.500000 351.590000 ;
      RECT 1157.500000 349.590000 1170.500000 350.410000 ;
      RECT 1107.500000 349.590000 1149.500000 350.410000 ;
      RECT 1057.500000 349.590000 1099.500000 350.410000 ;
      RECT 1007.500000 349.590000 1049.500000 350.410000 ;
      RECT 957.500000 349.590000 999.500000 350.410000 ;
      RECT 907.500000 349.590000 949.500000 350.410000 ;
      RECT 857.500000 349.590000 899.500000 350.410000 ;
      RECT 807.500000 349.590000 849.500000 350.410000 ;
      RECT 757.500000 349.590000 799.500000 350.410000 ;
      RECT 707.500000 349.590000 749.500000 350.410000 ;
      RECT 657.500000 349.590000 699.500000 350.410000 ;
      RECT 607.500000 349.590000 649.500000 350.410000 ;
      RECT 557.500000 349.590000 599.500000 350.410000 ;
      RECT 507.500000 349.590000 549.500000 350.410000 ;
      RECT 407.500000 349.590000 499.500000 350.410000 ;
      RECT 357.500000 349.590000 399.500000 350.410000 ;
      RECT 307.500000 349.590000 349.500000 350.410000 ;
      RECT 257.500000 349.590000 299.500000 350.410000 ;
      RECT 207.500000 349.590000 249.500000 350.410000 ;
      RECT 157.500000 349.590000 199.500000 350.410000 ;
      RECT 107.500000 349.590000 149.500000 350.410000 ;
      RECT 15.500000 349.590000 99.500000 350.410000 ;
      RECT 1183.500000 348.410000 1186.000000 351.590000 ;
      RECT 1169.500000 348.410000 1170.500000 349.590000 ;
      RECT 1116.500000 348.410000 1149.500000 349.590000 ;
      RECT 1107.500000 348.410000 1108.500000 349.590000 ;
      RECT 1066.500000 348.410000 1099.500000 349.590000 ;
      RECT 1057.500000 348.410000 1058.500000 349.590000 ;
      RECT 1016.500000 348.410000 1049.500000 349.590000 ;
      RECT 1007.500000 348.410000 1008.500000 349.590000 ;
      RECT 966.500000 348.410000 999.500000 349.590000 ;
      RECT 957.500000 348.410000 958.500000 349.590000 ;
      RECT 916.500000 348.410000 949.500000 349.590000 ;
      RECT 907.500000 348.410000 908.500000 349.590000 ;
      RECT 866.500000 348.410000 899.500000 349.590000 ;
      RECT 857.500000 348.410000 858.500000 349.590000 ;
      RECT 816.500000 348.410000 849.500000 349.590000 ;
      RECT 807.500000 348.410000 808.500000 349.590000 ;
      RECT 766.500000 348.410000 799.500000 349.590000 ;
      RECT 757.500000 348.410000 758.500000 349.590000 ;
      RECT 716.500000 348.410000 749.500000 349.590000 ;
      RECT 707.500000 348.410000 708.500000 349.590000 ;
      RECT 666.500000 348.410000 699.500000 349.590000 ;
      RECT 657.500000 348.410000 658.500000 349.590000 ;
      RECT 616.500000 348.410000 649.500000 349.590000 ;
      RECT 607.500000 348.410000 608.500000 349.590000 ;
      RECT 566.500000 348.410000 599.500000 349.590000 ;
      RECT 557.500000 348.410000 558.500000 349.590000 ;
      RECT 516.500000 348.410000 549.500000 349.590000 ;
      RECT 507.500000 348.410000 508.500000 349.590000 ;
      RECT 466.500000 348.410000 499.500000 349.590000 ;
      RECT 407.500000 348.410000 408.500000 349.590000 ;
      RECT 366.500000 348.410000 399.500000 349.590000 ;
      RECT 357.500000 348.410000 358.500000 349.590000 ;
      RECT 316.500000 348.410000 349.500000 349.590000 ;
      RECT 307.500000 348.410000 308.500000 349.590000 ;
      RECT 266.500000 348.410000 299.500000 349.590000 ;
      RECT 257.500000 348.410000 258.500000 349.590000 ;
      RECT 216.500000 348.410000 249.500000 349.590000 ;
      RECT 207.500000 348.410000 208.500000 349.590000 ;
      RECT 166.500000 348.410000 199.500000 349.590000 ;
      RECT 157.500000 348.410000 158.500000 349.590000 ;
      RECT 116.500000 348.410000 149.500000 349.590000 ;
      RECT 107.500000 348.410000 108.500000 349.590000 ;
      RECT 66.500000 348.410000 99.500000 349.590000 ;
      RECT 15.500000 348.410000 16.500000 349.590000 ;
      RECT 0.000000 348.410000 2.500000 351.590000 ;
      RECT 1169.500000 347.590000 1186.000000 348.410000 ;
      RECT 1116.500000 347.590000 1156.500000 348.410000 ;
      RECT 1066.500000 347.590000 1108.500000 348.410000 ;
      RECT 1016.500000 347.590000 1058.500000 348.410000 ;
      RECT 966.500000 347.590000 1008.500000 348.410000 ;
      RECT 916.500000 347.590000 958.500000 348.410000 ;
      RECT 866.500000 347.590000 908.500000 348.410000 ;
      RECT 816.500000 347.590000 858.500000 348.410000 ;
      RECT 766.500000 347.590000 808.500000 348.410000 ;
      RECT 716.500000 347.590000 758.500000 348.410000 ;
      RECT 666.500000 347.590000 708.500000 348.410000 ;
      RECT 616.500000 347.590000 658.500000 348.410000 ;
      RECT 566.500000 347.590000 608.500000 348.410000 ;
      RECT 516.500000 347.590000 558.500000 348.410000 ;
      RECT 466.500000 347.590000 508.500000 348.410000 ;
      RECT 416.500000 347.590000 458.500000 349.590000 ;
      RECT 366.500000 347.590000 408.500000 348.410000 ;
      RECT 316.500000 347.590000 358.500000 348.410000 ;
      RECT 266.500000 347.590000 308.500000 348.410000 ;
      RECT 216.500000 347.590000 258.500000 348.410000 ;
      RECT 166.500000 347.590000 208.500000 348.410000 ;
      RECT 116.500000 347.590000 158.500000 348.410000 ;
      RECT 66.500000 347.590000 108.500000 348.410000 ;
      RECT 29.500000 347.590000 58.500000 349.590000 ;
      RECT 0.000000 347.590000 16.500000 348.410000 ;
      RECT 1169.500000 346.410000 1170.500000 347.590000 ;
      RECT 1116.500000 346.410000 1149.500000 347.590000 ;
      RECT 1107.500000 346.410000 1108.500000 347.590000 ;
      RECT 1066.500000 346.410000 1099.500000 347.590000 ;
      RECT 1057.500000 346.410000 1058.500000 347.590000 ;
      RECT 1016.500000 346.410000 1049.500000 347.590000 ;
      RECT 1007.500000 346.410000 1008.500000 347.590000 ;
      RECT 966.500000 346.410000 999.500000 347.590000 ;
      RECT 957.500000 346.410000 958.500000 347.590000 ;
      RECT 916.500000 346.410000 949.500000 347.590000 ;
      RECT 907.500000 346.410000 908.500000 347.590000 ;
      RECT 866.500000 346.410000 899.500000 347.590000 ;
      RECT 857.500000 346.410000 858.500000 347.590000 ;
      RECT 816.500000 346.410000 849.500000 347.590000 ;
      RECT 807.500000 346.410000 808.500000 347.590000 ;
      RECT 766.500000 346.410000 799.500000 347.590000 ;
      RECT 757.500000 346.410000 758.500000 347.590000 ;
      RECT 716.500000 346.410000 749.500000 347.590000 ;
      RECT 707.500000 346.410000 708.500000 347.590000 ;
      RECT 666.500000 346.410000 699.500000 347.590000 ;
      RECT 657.500000 346.410000 658.500000 347.590000 ;
      RECT 616.500000 346.410000 649.500000 347.590000 ;
      RECT 607.500000 346.410000 608.500000 347.590000 ;
      RECT 566.500000 346.410000 599.500000 347.590000 ;
      RECT 557.500000 346.410000 558.500000 347.590000 ;
      RECT 516.500000 346.410000 549.500000 347.590000 ;
      RECT 507.500000 346.410000 508.500000 347.590000 ;
      RECT 466.500000 346.410000 499.500000 347.590000 ;
      RECT 457.500000 346.410000 458.500000 347.590000 ;
      RECT 416.500000 346.410000 449.500000 347.590000 ;
      RECT 407.500000 346.410000 408.500000 347.590000 ;
      RECT 366.500000 346.410000 399.500000 347.590000 ;
      RECT 357.500000 346.410000 358.500000 347.590000 ;
      RECT 316.500000 346.410000 349.500000 347.590000 ;
      RECT 307.500000 346.410000 308.500000 347.590000 ;
      RECT 266.500000 346.410000 299.500000 347.590000 ;
      RECT 257.500000 346.410000 258.500000 347.590000 ;
      RECT 216.500000 346.410000 249.500000 347.590000 ;
      RECT 207.500000 346.410000 208.500000 347.590000 ;
      RECT 166.500000 346.410000 199.500000 347.590000 ;
      RECT 157.500000 346.410000 158.500000 347.590000 ;
      RECT 116.500000 346.410000 149.500000 347.590000 ;
      RECT 107.500000 346.410000 108.500000 347.590000 ;
      RECT 66.500000 346.410000 99.500000 347.590000 ;
      RECT 57.500000 346.410000 58.500000 347.590000 ;
      RECT 29.500000 346.410000 49.500000 347.590000 ;
      RECT 15.500000 346.410000 16.500000 347.590000 ;
      RECT 1157.500000 345.590000 1170.500000 346.410000 ;
      RECT 1107.500000 345.590000 1149.500000 346.410000 ;
      RECT 1057.500000 345.590000 1099.500000 346.410000 ;
      RECT 1007.500000 345.590000 1049.500000 346.410000 ;
      RECT 957.500000 345.590000 999.500000 346.410000 ;
      RECT 907.500000 345.590000 949.500000 346.410000 ;
      RECT 857.500000 345.590000 899.500000 346.410000 ;
      RECT 807.500000 345.590000 849.500000 346.410000 ;
      RECT 757.500000 345.590000 799.500000 346.410000 ;
      RECT 707.500000 345.590000 749.500000 346.410000 ;
      RECT 657.500000 345.590000 699.500000 346.410000 ;
      RECT 607.500000 345.590000 649.500000 346.410000 ;
      RECT 557.500000 345.590000 599.500000 346.410000 ;
      RECT 507.500000 345.590000 549.500000 346.410000 ;
      RECT 457.500000 345.590000 499.500000 346.410000 ;
      RECT 407.500000 345.590000 449.500000 346.410000 ;
      RECT 357.500000 345.590000 399.500000 346.410000 ;
      RECT 307.500000 345.590000 349.500000 346.410000 ;
      RECT 257.500000 345.590000 299.500000 346.410000 ;
      RECT 207.500000 345.590000 249.500000 346.410000 ;
      RECT 157.500000 345.590000 199.500000 346.410000 ;
      RECT 107.500000 345.590000 149.500000 346.410000 ;
      RECT 57.500000 345.590000 99.500000 346.410000 ;
      RECT 15.500000 345.590000 49.500000 346.410000 ;
      RECT 1183.500000 344.410000 1186.000000 347.590000 ;
      RECT 1169.500000 344.410000 1170.500000 345.590000 ;
      RECT 1116.500000 344.410000 1149.500000 345.590000 ;
      RECT 1107.500000 344.410000 1108.500000 345.590000 ;
      RECT 1066.500000 344.410000 1099.500000 345.590000 ;
      RECT 1057.500000 344.410000 1058.500000 345.590000 ;
      RECT 1016.500000 344.410000 1049.500000 345.590000 ;
      RECT 1007.500000 344.410000 1008.500000 345.590000 ;
      RECT 966.500000 344.410000 999.500000 345.590000 ;
      RECT 957.500000 344.410000 958.500000 345.590000 ;
      RECT 916.500000 344.410000 949.500000 345.590000 ;
      RECT 907.500000 344.410000 908.500000 345.590000 ;
      RECT 866.500000 344.410000 899.500000 345.590000 ;
      RECT 857.500000 344.410000 858.500000 345.590000 ;
      RECT 816.500000 344.410000 849.500000 345.590000 ;
      RECT 807.500000 344.410000 808.500000 345.590000 ;
      RECT 766.500000 344.410000 799.500000 345.590000 ;
      RECT 757.500000 344.410000 758.500000 345.590000 ;
      RECT 716.500000 344.410000 749.500000 345.590000 ;
      RECT 707.500000 344.410000 708.500000 345.590000 ;
      RECT 666.500000 344.410000 699.500000 345.590000 ;
      RECT 657.500000 344.410000 658.500000 345.590000 ;
      RECT 616.500000 344.410000 649.500000 345.590000 ;
      RECT 607.500000 344.410000 608.500000 345.590000 ;
      RECT 566.500000 344.410000 599.500000 345.590000 ;
      RECT 557.500000 344.410000 558.500000 345.590000 ;
      RECT 516.500000 344.410000 549.500000 345.590000 ;
      RECT 507.500000 344.410000 508.500000 345.590000 ;
      RECT 466.500000 344.410000 499.500000 345.590000 ;
      RECT 457.500000 344.410000 458.500000 345.590000 ;
      RECT 416.500000 344.410000 449.500000 345.590000 ;
      RECT 407.500000 344.410000 408.500000 345.590000 ;
      RECT 366.500000 344.410000 399.500000 345.590000 ;
      RECT 357.500000 344.410000 358.500000 345.590000 ;
      RECT 316.500000 344.410000 349.500000 345.590000 ;
      RECT 307.500000 344.410000 308.500000 345.590000 ;
      RECT 266.500000 344.410000 299.500000 345.590000 ;
      RECT 257.500000 344.410000 258.500000 345.590000 ;
      RECT 216.500000 344.410000 249.500000 345.590000 ;
      RECT 207.500000 344.410000 208.500000 345.590000 ;
      RECT 166.500000 344.410000 199.500000 345.590000 ;
      RECT 157.500000 344.410000 158.500000 345.590000 ;
      RECT 116.500000 344.410000 149.500000 345.590000 ;
      RECT 107.500000 344.410000 108.500000 345.590000 ;
      RECT 66.500000 344.410000 99.500000 345.590000 ;
      RECT 57.500000 344.410000 58.500000 345.590000 ;
      RECT 29.500000 344.410000 49.500000 345.590000 ;
      RECT 15.500000 344.410000 16.500000 345.590000 ;
      RECT 0.000000 344.410000 2.500000 347.590000 ;
      RECT 1169.500000 343.590000 1186.000000 344.410000 ;
      RECT 1116.500000 343.590000 1156.500000 344.410000 ;
      RECT 1066.500000 343.590000 1108.500000 344.410000 ;
      RECT 1016.500000 343.590000 1058.500000 344.410000 ;
      RECT 966.500000 343.590000 1008.500000 344.410000 ;
      RECT 916.500000 343.590000 958.500000 344.410000 ;
      RECT 866.500000 343.590000 908.500000 344.410000 ;
      RECT 816.500000 343.590000 858.500000 344.410000 ;
      RECT 766.500000 343.590000 808.500000 344.410000 ;
      RECT 716.500000 343.590000 758.500000 344.410000 ;
      RECT 666.500000 343.590000 708.500000 344.410000 ;
      RECT 616.500000 343.590000 658.500000 344.410000 ;
      RECT 566.500000 343.590000 608.500000 344.410000 ;
      RECT 516.500000 343.590000 558.500000 344.410000 ;
      RECT 466.500000 343.590000 508.500000 344.410000 ;
      RECT 416.500000 343.590000 458.500000 344.410000 ;
      RECT 366.500000 343.590000 408.500000 344.410000 ;
      RECT 316.500000 343.590000 358.500000 344.410000 ;
      RECT 266.500000 343.590000 308.500000 344.410000 ;
      RECT 216.500000 343.590000 258.500000 344.410000 ;
      RECT 166.500000 343.590000 208.500000 344.410000 ;
      RECT 116.500000 343.590000 158.500000 344.410000 ;
      RECT 66.500000 343.590000 108.500000 344.410000 ;
      RECT 29.500000 343.590000 58.500000 344.410000 ;
      RECT 0.000000 343.590000 16.500000 344.410000 ;
      RECT 1169.500000 342.410000 1170.500000 343.590000 ;
      RECT 1116.500000 342.410000 1149.500000 343.590000 ;
      RECT 1107.500000 342.410000 1108.500000 343.590000 ;
      RECT 1066.500000 342.410000 1099.500000 343.590000 ;
      RECT 1057.500000 342.410000 1058.500000 343.590000 ;
      RECT 1016.500000 342.410000 1049.500000 343.590000 ;
      RECT 1007.500000 342.410000 1008.500000 343.590000 ;
      RECT 966.500000 342.410000 999.500000 343.590000 ;
      RECT 957.500000 342.410000 958.500000 343.590000 ;
      RECT 916.500000 342.410000 949.500000 343.590000 ;
      RECT 907.500000 342.410000 908.500000 343.590000 ;
      RECT 866.500000 342.410000 899.500000 343.590000 ;
      RECT 857.500000 342.410000 858.500000 343.590000 ;
      RECT 816.500000 342.410000 849.500000 343.590000 ;
      RECT 807.500000 342.410000 808.500000 343.590000 ;
      RECT 766.500000 342.410000 799.500000 343.590000 ;
      RECT 757.500000 342.410000 758.500000 343.590000 ;
      RECT 716.500000 342.410000 749.500000 343.590000 ;
      RECT 707.500000 342.410000 708.500000 343.590000 ;
      RECT 666.500000 342.410000 699.500000 343.590000 ;
      RECT 657.500000 342.410000 658.500000 343.590000 ;
      RECT 616.500000 342.410000 649.500000 343.590000 ;
      RECT 607.500000 342.410000 608.500000 343.590000 ;
      RECT 566.500000 342.410000 599.500000 343.590000 ;
      RECT 557.500000 342.410000 558.500000 343.590000 ;
      RECT 516.500000 342.410000 549.500000 343.590000 ;
      RECT 507.500000 342.410000 508.500000 343.590000 ;
      RECT 466.500000 342.410000 499.500000 343.590000 ;
      RECT 457.500000 342.410000 458.500000 343.590000 ;
      RECT 416.500000 342.410000 449.500000 343.590000 ;
      RECT 407.500000 342.410000 408.500000 343.590000 ;
      RECT 366.500000 342.410000 399.500000 343.590000 ;
      RECT 357.500000 342.410000 358.500000 343.590000 ;
      RECT 316.500000 342.410000 349.500000 343.590000 ;
      RECT 307.500000 342.410000 308.500000 343.590000 ;
      RECT 266.500000 342.410000 299.500000 343.590000 ;
      RECT 257.500000 342.410000 258.500000 343.590000 ;
      RECT 216.500000 342.410000 249.500000 343.590000 ;
      RECT 207.500000 342.410000 208.500000 343.590000 ;
      RECT 166.500000 342.410000 199.500000 343.590000 ;
      RECT 157.500000 342.410000 158.500000 343.590000 ;
      RECT 116.500000 342.410000 149.500000 343.590000 ;
      RECT 107.500000 342.410000 108.500000 343.590000 ;
      RECT 66.500000 342.410000 99.500000 343.590000 ;
      RECT 57.500000 342.410000 58.500000 343.590000 ;
      RECT 29.500000 342.410000 49.500000 343.590000 ;
      RECT 15.500000 342.410000 16.500000 343.590000 ;
      RECT 1157.500000 341.590000 1170.500000 342.410000 ;
      RECT 1107.500000 341.590000 1149.500000 342.410000 ;
      RECT 1057.500000 341.590000 1099.500000 342.410000 ;
      RECT 1007.500000 341.590000 1049.500000 342.410000 ;
      RECT 957.500000 341.590000 999.500000 342.410000 ;
      RECT 907.500000 341.590000 949.500000 342.410000 ;
      RECT 857.500000 341.590000 899.500000 342.410000 ;
      RECT 807.500000 341.590000 849.500000 342.410000 ;
      RECT 757.500000 341.590000 799.500000 342.410000 ;
      RECT 707.500000 341.590000 749.500000 342.410000 ;
      RECT 657.500000 341.590000 699.500000 342.410000 ;
      RECT 607.500000 341.590000 649.500000 342.410000 ;
      RECT 557.500000 341.590000 599.500000 342.410000 ;
      RECT 507.500000 341.590000 549.500000 342.410000 ;
      RECT 457.500000 341.590000 499.500000 342.410000 ;
      RECT 407.500000 341.590000 449.500000 342.410000 ;
      RECT 357.500000 341.590000 399.500000 342.410000 ;
      RECT 307.500000 341.590000 349.500000 342.410000 ;
      RECT 257.500000 341.590000 299.500000 342.410000 ;
      RECT 207.500000 341.590000 249.500000 342.410000 ;
      RECT 157.500000 341.590000 199.500000 342.410000 ;
      RECT 107.500000 341.590000 149.500000 342.410000 ;
      RECT 57.500000 341.590000 99.500000 342.410000 ;
      RECT 15.500000 341.590000 49.500000 342.410000 ;
      RECT 1183.500000 340.410000 1186.000000 343.590000 ;
      RECT 1169.500000 340.410000 1170.500000 341.590000 ;
      RECT 1116.500000 340.410000 1149.500000 341.590000 ;
      RECT 1107.500000 340.410000 1108.500000 341.590000 ;
      RECT 1066.500000 340.410000 1099.500000 341.590000 ;
      RECT 1057.500000 340.410000 1058.500000 341.590000 ;
      RECT 1016.500000 340.410000 1049.500000 341.590000 ;
      RECT 1007.500000 340.410000 1008.500000 341.590000 ;
      RECT 966.500000 340.410000 999.500000 341.590000 ;
      RECT 957.500000 340.410000 958.500000 341.590000 ;
      RECT 916.500000 340.410000 949.500000 341.590000 ;
      RECT 907.500000 340.410000 908.500000 341.590000 ;
      RECT 866.500000 340.410000 899.500000 341.590000 ;
      RECT 857.500000 340.410000 858.500000 341.590000 ;
      RECT 816.500000 340.410000 849.500000 341.590000 ;
      RECT 807.500000 340.410000 808.500000 341.590000 ;
      RECT 766.500000 340.410000 799.500000 341.590000 ;
      RECT 757.500000 340.410000 758.500000 341.590000 ;
      RECT 716.500000 340.410000 749.500000 341.590000 ;
      RECT 707.500000 340.410000 708.500000 341.590000 ;
      RECT 666.500000 340.410000 699.500000 341.590000 ;
      RECT 657.500000 340.410000 658.500000 341.590000 ;
      RECT 616.500000 340.410000 649.500000 341.590000 ;
      RECT 607.500000 340.410000 608.500000 341.590000 ;
      RECT 566.500000 340.410000 599.500000 341.590000 ;
      RECT 557.500000 340.410000 558.500000 341.590000 ;
      RECT 516.500000 340.410000 549.500000 341.590000 ;
      RECT 507.500000 340.410000 508.500000 341.590000 ;
      RECT 466.500000 340.410000 499.500000 341.590000 ;
      RECT 457.500000 340.410000 458.500000 341.590000 ;
      RECT 416.500000 340.410000 449.500000 341.590000 ;
      RECT 407.500000 340.410000 408.500000 341.590000 ;
      RECT 366.500000 340.410000 399.500000 341.590000 ;
      RECT 357.500000 340.410000 358.500000 341.590000 ;
      RECT 316.500000 340.410000 349.500000 341.590000 ;
      RECT 307.500000 340.410000 308.500000 341.590000 ;
      RECT 266.500000 340.410000 299.500000 341.590000 ;
      RECT 257.500000 340.410000 258.500000 341.590000 ;
      RECT 216.500000 340.410000 249.500000 341.590000 ;
      RECT 207.500000 340.410000 208.500000 341.590000 ;
      RECT 166.500000 340.410000 199.500000 341.590000 ;
      RECT 157.500000 340.410000 158.500000 341.590000 ;
      RECT 116.500000 340.410000 149.500000 341.590000 ;
      RECT 107.500000 340.410000 108.500000 341.590000 ;
      RECT 66.500000 340.410000 99.500000 341.590000 ;
      RECT 57.500000 340.410000 58.500000 341.590000 ;
      RECT 29.500000 340.410000 49.500000 341.590000 ;
      RECT 15.500000 340.410000 16.500000 341.590000 ;
      RECT 0.000000 340.410000 2.500000 343.590000 ;
      RECT 1169.500000 339.590000 1186.000000 340.410000 ;
      RECT 1116.500000 339.590000 1156.500000 340.410000 ;
      RECT 1066.500000 339.590000 1108.500000 340.410000 ;
      RECT 1016.500000 339.590000 1058.500000 340.410000 ;
      RECT 966.500000 339.590000 1008.500000 340.410000 ;
      RECT 916.500000 339.590000 958.500000 340.410000 ;
      RECT 866.500000 339.590000 908.500000 340.410000 ;
      RECT 816.500000 339.590000 858.500000 340.410000 ;
      RECT 766.500000 339.590000 808.500000 340.410000 ;
      RECT 716.500000 339.590000 758.500000 340.410000 ;
      RECT 666.500000 339.590000 708.500000 340.410000 ;
      RECT 616.500000 339.590000 658.500000 340.410000 ;
      RECT 566.500000 339.590000 608.500000 340.410000 ;
      RECT 516.500000 339.590000 558.500000 340.410000 ;
      RECT 466.500000 339.590000 508.500000 340.410000 ;
      RECT 416.500000 339.590000 458.500000 340.410000 ;
      RECT 366.500000 339.590000 408.500000 340.410000 ;
      RECT 316.500000 339.590000 358.500000 340.410000 ;
      RECT 266.500000 339.590000 308.500000 340.410000 ;
      RECT 216.500000 339.590000 258.500000 340.410000 ;
      RECT 166.500000 339.590000 208.500000 340.410000 ;
      RECT 116.500000 339.590000 158.500000 340.410000 ;
      RECT 66.500000 339.590000 108.500000 340.410000 ;
      RECT 29.500000 339.590000 58.500000 340.410000 ;
      RECT 0.000000 339.590000 16.500000 340.410000 ;
      RECT 1169.500000 338.410000 1170.500000 339.590000 ;
      RECT 1116.500000 338.410000 1149.500000 339.590000 ;
      RECT 1107.500000 338.410000 1108.500000 339.590000 ;
      RECT 1066.500000 338.410000 1099.500000 339.590000 ;
      RECT 1057.500000 338.410000 1058.500000 339.590000 ;
      RECT 1016.500000 338.410000 1049.500000 339.590000 ;
      RECT 1007.500000 338.410000 1008.500000 339.590000 ;
      RECT 966.500000 338.410000 999.500000 339.590000 ;
      RECT 957.500000 338.410000 958.500000 339.590000 ;
      RECT 916.500000 338.410000 949.500000 339.590000 ;
      RECT 907.500000 338.410000 908.500000 339.590000 ;
      RECT 866.500000 338.410000 899.500000 339.590000 ;
      RECT 857.500000 338.410000 858.500000 339.590000 ;
      RECT 816.500000 338.410000 849.500000 339.590000 ;
      RECT 807.500000 338.410000 808.500000 339.590000 ;
      RECT 766.500000 338.410000 799.500000 339.590000 ;
      RECT 757.500000 338.410000 758.500000 339.590000 ;
      RECT 716.500000 338.410000 749.500000 339.590000 ;
      RECT 707.500000 338.410000 708.500000 339.590000 ;
      RECT 666.500000 338.410000 699.500000 339.590000 ;
      RECT 657.500000 338.410000 658.500000 339.590000 ;
      RECT 616.500000 338.410000 649.500000 339.590000 ;
      RECT 607.500000 338.410000 608.500000 339.590000 ;
      RECT 566.500000 338.410000 599.500000 339.590000 ;
      RECT 557.500000 338.410000 558.500000 339.590000 ;
      RECT 516.500000 338.410000 549.500000 339.590000 ;
      RECT 507.500000 338.410000 508.500000 339.590000 ;
      RECT 466.500000 338.410000 499.500000 339.590000 ;
      RECT 457.500000 338.410000 458.500000 339.590000 ;
      RECT 416.500000 338.410000 449.500000 339.590000 ;
      RECT 407.500000 338.410000 408.500000 339.590000 ;
      RECT 366.500000 338.410000 399.500000 339.590000 ;
      RECT 357.500000 338.410000 358.500000 339.590000 ;
      RECT 316.500000 338.410000 349.500000 339.590000 ;
      RECT 307.500000 338.410000 308.500000 339.590000 ;
      RECT 266.500000 338.410000 299.500000 339.590000 ;
      RECT 257.500000 338.410000 258.500000 339.590000 ;
      RECT 216.500000 338.410000 249.500000 339.590000 ;
      RECT 207.500000 338.410000 208.500000 339.590000 ;
      RECT 166.500000 338.410000 199.500000 339.590000 ;
      RECT 157.500000 338.410000 158.500000 339.590000 ;
      RECT 116.500000 338.410000 149.500000 339.590000 ;
      RECT 107.500000 338.410000 108.500000 339.590000 ;
      RECT 66.500000 338.410000 99.500000 339.590000 ;
      RECT 57.500000 338.410000 58.500000 339.590000 ;
      RECT 29.500000 338.410000 49.500000 339.590000 ;
      RECT 15.500000 338.410000 16.500000 339.590000 ;
      RECT 1157.500000 337.590000 1170.500000 338.410000 ;
      RECT 1107.500000 337.590000 1149.500000 338.410000 ;
      RECT 1057.500000 337.590000 1099.500000 338.410000 ;
      RECT 1007.500000 337.590000 1049.500000 338.410000 ;
      RECT 957.500000 337.590000 999.500000 338.410000 ;
      RECT 907.500000 337.590000 949.500000 338.410000 ;
      RECT 857.500000 337.590000 899.500000 338.410000 ;
      RECT 807.500000 337.590000 849.500000 338.410000 ;
      RECT 757.500000 337.590000 799.500000 338.410000 ;
      RECT 707.500000 337.590000 749.500000 338.410000 ;
      RECT 657.500000 337.590000 699.500000 338.410000 ;
      RECT 607.500000 337.590000 649.500000 338.410000 ;
      RECT 557.500000 337.590000 599.500000 338.410000 ;
      RECT 507.500000 337.590000 549.500000 338.410000 ;
      RECT 457.500000 337.590000 499.500000 338.410000 ;
      RECT 407.500000 337.590000 449.500000 338.410000 ;
      RECT 357.500000 337.590000 399.500000 338.410000 ;
      RECT 307.500000 337.590000 349.500000 338.410000 ;
      RECT 257.500000 337.590000 299.500000 338.410000 ;
      RECT 207.500000 337.590000 249.500000 338.410000 ;
      RECT 157.500000 337.590000 199.500000 338.410000 ;
      RECT 107.500000 337.590000 149.500000 338.410000 ;
      RECT 57.500000 337.590000 99.500000 338.410000 ;
      RECT 15.500000 337.590000 49.500000 338.410000 ;
      RECT 1183.500000 336.410000 1186.000000 339.590000 ;
      RECT 1169.500000 336.410000 1170.500000 337.590000 ;
      RECT 1116.500000 336.410000 1149.500000 337.590000 ;
      RECT 1107.500000 336.410000 1108.500000 337.590000 ;
      RECT 1066.500000 336.410000 1099.500000 337.590000 ;
      RECT 1057.500000 336.410000 1058.500000 337.590000 ;
      RECT 1016.500000 336.410000 1049.500000 337.590000 ;
      RECT 1007.500000 336.410000 1008.500000 337.590000 ;
      RECT 966.500000 336.410000 999.500000 337.590000 ;
      RECT 957.500000 336.410000 958.500000 337.590000 ;
      RECT 916.500000 336.410000 949.500000 337.590000 ;
      RECT 907.500000 336.410000 908.500000 337.590000 ;
      RECT 866.500000 336.410000 899.500000 337.590000 ;
      RECT 857.500000 336.410000 858.500000 337.590000 ;
      RECT 816.500000 336.410000 849.500000 337.590000 ;
      RECT 807.500000 336.410000 808.500000 337.590000 ;
      RECT 766.500000 336.410000 799.500000 337.590000 ;
      RECT 757.500000 336.410000 758.500000 337.590000 ;
      RECT 716.500000 336.410000 749.500000 337.590000 ;
      RECT 707.500000 336.410000 708.500000 337.590000 ;
      RECT 666.500000 336.410000 699.500000 337.590000 ;
      RECT 657.500000 336.410000 658.500000 337.590000 ;
      RECT 616.500000 336.410000 649.500000 337.590000 ;
      RECT 607.500000 336.410000 608.500000 337.590000 ;
      RECT 566.500000 336.410000 599.500000 337.590000 ;
      RECT 557.500000 336.410000 558.500000 337.590000 ;
      RECT 516.500000 336.410000 549.500000 337.590000 ;
      RECT 507.500000 336.410000 508.500000 337.590000 ;
      RECT 466.500000 336.410000 499.500000 337.590000 ;
      RECT 457.500000 336.410000 458.500000 337.590000 ;
      RECT 416.500000 336.410000 449.500000 337.590000 ;
      RECT 407.500000 336.410000 408.500000 337.590000 ;
      RECT 366.500000 336.410000 399.500000 337.590000 ;
      RECT 357.500000 336.410000 358.500000 337.590000 ;
      RECT 316.500000 336.410000 349.500000 337.590000 ;
      RECT 307.500000 336.410000 308.500000 337.590000 ;
      RECT 266.500000 336.410000 299.500000 337.590000 ;
      RECT 257.500000 336.410000 258.500000 337.590000 ;
      RECT 216.500000 336.410000 249.500000 337.590000 ;
      RECT 207.500000 336.410000 208.500000 337.590000 ;
      RECT 166.500000 336.410000 199.500000 337.590000 ;
      RECT 157.500000 336.410000 158.500000 337.590000 ;
      RECT 116.500000 336.410000 149.500000 337.590000 ;
      RECT 107.500000 336.410000 108.500000 337.590000 ;
      RECT 66.500000 336.410000 99.500000 337.590000 ;
      RECT 57.500000 336.410000 58.500000 337.590000 ;
      RECT 29.500000 336.410000 49.500000 337.590000 ;
      RECT 15.500000 336.410000 16.500000 337.590000 ;
      RECT 0.000000 336.410000 2.500000 339.590000 ;
      RECT 1169.500000 335.590000 1186.000000 336.410000 ;
      RECT 1116.500000 335.590000 1156.500000 336.410000 ;
      RECT 1066.500000 335.590000 1108.500000 336.410000 ;
      RECT 1016.500000 335.590000 1058.500000 336.410000 ;
      RECT 966.500000 335.590000 1008.500000 336.410000 ;
      RECT 916.500000 335.590000 958.500000 336.410000 ;
      RECT 866.500000 335.590000 908.500000 336.410000 ;
      RECT 816.500000 335.590000 858.500000 336.410000 ;
      RECT 766.500000 335.590000 808.500000 336.410000 ;
      RECT 716.500000 335.590000 758.500000 336.410000 ;
      RECT 666.500000 335.590000 708.500000 336.410000 ;
      RECT 616.500000 335.590000 658.500000 336.410000 ;
      RECT 566.500000 335.590000 608.500000 336.410000 ;
      RECT 516.500000 335.590000 558.500000 336.410000 ;
      RECT 466.500000 335.590000 508.500000 336.410000 ;
      RECT 416.500000 335.590000 458.500000 336.410000 ;
      RECT 366.500000 335.590000 408.500000 336.410000 ;
      RECT 316.500000 335.590000 358.500000 336.410000 ;
      RECT 266.500000 335.590000 308.500000 336.410000 ;
      RECT 216.500000 335.590000 258.500000 336.410000 ;
      RECT 166.500000 335.590000 208.500000 336.410000 ;
      RECT 116.500000 335.590000 158.500000 336.410000 ;
      RECT 66.500000 335.590000 108.500000 336.410000 ;
      RECT 29.500000 335.590000 58.500000 336.410000 ;
      RECT 0.000000 335.590000 16.500000 336.410000 ;
      RECT 1169.500000 334.410000 1170.500000 335.590000 ;
      RECT 1116.500000 334.410000 1149.500000 335.590000 ;
      RECT 1107.500000 334.410000 1108.500000 335.590000 ;
      RECT 1066.500000 334.410000 1099.500000 335.590000 ;
      RECT 1057.500000 334.410000 1058.500000 335.590000 ;
      RECT 1016.500000 334.410000 1049.500000 335.590000 ;
      RECT 1007.500000 334.410000 1008.500000 335.590000 ;
      RECT 966.500000 334.410000 999.500000 335.590000 ;
      RECT 957.500000 334.410000 958.500000 335.590000 ;
      RECT 916.500000 334.410000 949.500000 335.590000 ;
      RECT 907.500000 334.410000 908.500000 335.590000 ;
      RECT 866.500000 334.410000 899.500000 335.590000 ;
      RECT 857.500000 334.410000 858.500000 335.590000 ;
      RECT 816.500000 334.410000 849.500000 335.590000 ;
      RECT 807.500000 334.410000 808.500000 335.590000 ;
      RECT 766.500000 334.410000 799.500000 335.590000 ;
      RECT 757.500000 334.410000 758.500000 335.590000 ;
      RECT 716.500000 334.410000 749.500000 335.590000 ;
      RECT 707.500000 334.410000 708.500000 335.590000 ;
      RECT 666.500000 334.410000 699.500000 335.590000 ;
      RECT 657.500000 334.410000 658.500000 335.590000 ;
      RECT 616.500000 334.410000 649.500000 335.590000 ;
      RECT 607.500000 334.410000 608.500000 335.590000 ;
      RECT 566.500000 334.410000 599.500000 335.590000 ;
      RECT 557.500000 334.410000 558.500000 335.590000 ;
      RECT 516.500000 334.410000 549.500000 335.590000 ;
      RECT 507.500000 334.410000 508.500000 335.590000 ;
      RECT 466.500000 334.410000 499.500000 335.590000 ;
      RECT 457.500000 334.410000 458.500000 335.590000 ;
      RECT 416.500000 334.410000 449.500000 335.590000 ;
      RECT 407.500000 334.410000 408.500000 335.590000 ;
      RECT 366.500000 334.410000 399.500000 335.590000 ;
      RECT 357.500000 334.410000 358.500000 335.590000 ;
      RECT 316.500000 334.410000 349.500000 335.590000 ;
      RECT 307.500000 334.410000 308.500000 335.590000 ;
      RECT 266.500000 334.410000 299.500000 335.590000 ;
      RECT 257.500000 334.410000 258.500000 335.590000 ;
      RECT 216.500000 334.410000 249.500000 335.590000 ;
      RECT 207.500000 334.410000 208.500000 335.590000 ;
      RECT 166.500000 334.410000 199.500000 335.590000 ;
      RECT 157.500000 334.410000 158.500000 335.590000 ;
      RECT 116.500000 334.410000 149.500000 335.590000 ;
      RECT 107.500000 334.410000 108.500000 335.590000 ;
      RECT 66.500000 334.410000 99.500000 335.590000 ;
      RECT 57.500000 334.410000 58.500000 335.590000 ;
      RECT 29.500000 334.410000 49.500000 335.590000 ;
      RECT 15.500000 334.410000 16.500000 335.590000 ;
      RECT 1157.500000 333.590000 1170.500000 334.410000 ;
      RECT 1107.500000 333.590000 1149.500000 334.410000 ;
      RECT 1057.500000 333.590000 1099.500000 334.410000 ;
      RECT 1007.500000 333.590000 1049.500000 334.410000 ;
      RECT 957.500000 333.590000 999.500000 334.410000 ;
      RECT 907.500000 333.590000 949.500000 334.410000 ;
      RECT 857.500000 333.590000 899.500000 334.410000 ;
      RECT 807.500000 333.590000 849.500000 334.410000 ;
      RECT 757.500000 333.590000 799.500000 334.410000 ;
      RECT 707.500000 333.590000 749.500000 334.410000 ;
      RECT 657.500000 333.590000 699.500000 334.410000 ;
      RECT 607.500000 333.590000 649.500000 334.410000 ;
      RECT 557.500000 333.590000 599.500000 334.410000 ;
      RECT 507.500000 333.590000 549.500000 334.410000 ;
      RECT 457.500000 333.590000 499.500000 334.410000 ;
      RECT 407.500000 333.590000 449.500000 334.410000 ;
      RECT 357.500000 333.590000 399.500000 334.410000 ;
      RECT 307.500000 333.590000 349.500000 334.410000 ;
      RECT 257.500000 333.590000 299.500000 334.410000 ;
      RECT 207.500000 333.590000 249.500000 334.410000 ;
      RECT 157.500000 333.590000 199.500000 334.410000 ;
      RECT 107.500000 333.590000 149.500000 334.410000 ;
      RECT 57.500000 333.590000 99.500000 334.410000 ;
      RECT 15.500000 333.590000 49.500000 334.410000 ;
      RECT 1183.500000 332.410000 1186.000000 335.590000 ;
      RECT 1169.500000 332.410000 1170.500000 333.590000 ;
      RECT 1116.500000 332.410000 1149.500000 333.590000 ;
      RECT 1107.500000 332.410000 1108.500000 333.590000 ;
      RECT 1066.500000 332.410000 1099.500000 333.590000 ;
      RECT 1057.500000 332.410000 1058.500000 333.590000 ;
      RECT 1016.500000 332.410000 1049.500000 333.590000 ;
      RECT 1007.500000 332.410000 1008.500000 333.590000 ;
      RECT 966.500000 332.410000 999.500000 333.590000 ;
      RECT 957.500000 332.410000 958.500000 333.590000 ;
      RECT 916.500000 332.410000 949.500000 333.590000 ;
      RECT 907.500000 332.410000 908.500000 333.590000 ;
      RECT 866.500000 332.410000 899.500000 333.590000 ;
      RECT 857.500000 332.410000 858.500000 333.590000 ;
      RECT 816.500000 332.410000 849.500000 333.590000 ;
      RECT 807.500000 332.410000 808.500000 333.590000 ;
      RECT 766.500000 332.410000 799.500000 333.590000 ;
      RECT 757.500000 332.410000 758.500000 333.590000 ;
      RECT 716.500000 332.410000 749.500000 333.590000 ;
      RECT 707.500000 332.410000 708.500000 333.590000 ;
      RECT 666.500000 332.410000 699.500000 333.590000 ;
      RECT 657.500000 332.410000 658.500000 333.590000 ;
      RECT 616.500000 332.410000 649.500000 333.590000 ;
      RECT 607.500000 332.410000 608.500000 333.590000 ;
      RECT 566.500000 332.410000 599.500000 333.590000 ;
      RECT 557.500000 332.410000 558.500000 333.590000 ;
      RECT 516.500000 332.410000 549.500000 333.590000 ;
      RECT 507.500000 332.410000 508.500000 333.590000 ;
      RECT 466.500000 332.410000 499.500000 333.590000 ;
      RECT 457.500000 332.410000 458.500000 333.590000 ;
      RECT 416.500000 332.410000 449.500000 333.590000 ;
      RECT 407.500000 332.410000 408.500000 333.590000 ;
      RECT 366.500000 332.410000 399.500000 333.590000 ;
      RECT 357.500000 332.410000 358.500000 333.590000 ;
      RECT 316.500000 332.410000 349.500000 333.590000 ;
      RECT 307.500000 332.410000 308.500000 333.590000 ;
      RECT 266.500000 332.410000 299.500000 333.590000 ;
      RECT 257.500000 332.410000 258.500000 333.590000 ;
      RECT 216.500000 332.410000 249.500000 333.590000 ;
      RECT 207.500000 332.410000 208.500000 333.590000 ;
      RECT 166.500000 332.410000 199.500000 333.590000 ;
      RECT 157.500000 332.410000 158.500000 333.590000 ;
      RECT 116.500000 332.410000 149.500000 333.590000 ;
      RECT 107.500000 332.410000 108.500000 333.590000 ;
      RECT 66.500000 332.410000 99.500000 333.590000 ;
      RECT 57.500000 332.410000 58.500000 333.590000 ;
      RECT 29.500000 332.410000 49.500000 333.590000 ;
      RECT 15.500000 332.410000 16.500000 333.590000 ;
      RECT 0.000000 332.410000 2.500000 335.590000 ;
      RECT 1169.500000 331.590000 1186.000000 332.410000 ;
      RECT 1116.500000 331.590000 1156.500000 332.410000 ;
      RECT 1066.500000 331.590000 1108.500000 332.410000 ;
      RECT 1016.500000 331.590000 1058.500000 332.410000 ;
      RECT 966.500000 331.590000 1008.500000 332.410000 ;
      RECT 916.500000 331.590000 958.500000 332.410000 ;
      RECT 866.500000 331.590000 908.500000 332.410000 ;
      RECT 816.500000 331.590000 858.500000 332.410000 ;
      RECT 766.500000 331.590000 808.500000 332.410000 ;
      RECT 716.500000 331.590000 758.500000 332.410000 ;
      RECT 666.500000 331.590000 708.500000 332.410000 ;
      RECT 616.500000 331.590000 658.500000 332.410000 ;
      RECT 566.500000 331.590000 608.500000 332.410000 ;
      RECT 516.500000 331.590000 558.500000 332.410000 ;
      RECT 466.500000 331.590000 508.500000 332.410000 ;
      RECT 416.500000 331.590000 458.500000 332.410000 ;
      RECT 366.500000 331.590000 408.500000 332.410000 ;
      RECT 316.500000 331.590000 358.500000 332.410000 ;
      RECT 266.500000 331.590000 308.500000 332.410000 ;
      RECT 216.500000 331.590000 258.500000 332.410000 ;
      RECT 166.500000 331.590000 208.500000 332.410000 ;
      RECT 116.500000 331.590000 158.500000 332.410000 ;
      RECT 66.500000 331.590000 108.500000 332.410000 ;
      RECT 29.500000 331.590000 58.500000 332.410000 ;
      RECT 0.000000 331.590000 16.500000 332.410000 ;
      RECT 1169.500000 330.410000 1170.500000 331.590000 ;
      RECT 1116.500000 330.410000 1149.500000 331.590000 ;
      RECT 1107.500000 330.410000 1108.500000 331.590000 ;
      RECT 1066.500000 330.410000 1099.500000 331.590000 ;
      RECT 1057.500000 330.410000 1058.500000 331.590000 ;
      RECT 1016.500000 330.410000 1049.500000 331.590000 ;
      RECT 1007.500000 330.410000 1008.500000 331.590000 ;
      RECT 966.500000 330.410000 999.500000 331.590000 ;
      RECT 957.500000 330.410000 958.500000 331.590000 ;
      RECT 916.500000 330.410000 949.500000 331.590000 ;
      RECT 907.500000 330.410000 908.500000 331.590000 ;
      RECT 866.500000 330.410000 899.500000 331.590000 ;
      RECT 857.500000 330.410000 858.500000 331.590000 ;
      RECT 816.500000 330.410000 849.500000 331.590000 ;
      RECT 807.500000 330.410000 808.500000 331.590000 ;
      RECT 766.500000 330.410000 799.500000 331.590000 ;
      RECT 757.500000 330.410000 758.500000 331.590000 ;
      RECT 716.500000 330.410000 749.500000 331.590000 ;
      RECT 707.500000 330.410000 708.500000 331.590000 ;
      RECT 666.500000 330.410000 699.500000 331.590000 ;
      RECT 657.500000 330.410000 658.500000 331.590000 ;
      RECT 616.500000 330.410000 649.500000 331.590000 ;
      RECT 607.500000 330.410000 608.500000 331.590000 ;
      RECT 566.500000 330.410000 599.500000 331.590000 ;
      RECT 557.500000 330.410000 558.500000 331.590000 ;
      RECT 516.500000 330.410000 549.500000 331.590000 ;
      RECT 507.500000 330.410000 508.500000 331.590000 ;
      RECT 466.500000 330.410000 499.500000 331.590000 ;
      RECT 457.500000 330.410000 458.500000 331.590000 ;
      RECT 416.500000 330.410000 449.500000 331.590000 ;
      RECT 407.500000 330.410000 408.500000 331.590000 ;
      RECT 366.500000 330.410000 399.500000 331.590000 ;
      RECT 357.500000 330.410000 358.500000 331.590000 ;
      RECT 316.500000 330.410000 349.500000 331.590000 ;
      RECT 307.500000 330.410000 308.500000 331.590000 ;
      RECT 266.500000 330.410000 299.500000 331.590000 ;
      RECT 257.500000 330.410000 258.500000 331.590000 ;
      RECT 216.500000 330.410000 249.500000 331.590000 ;
      RECT 207.500000 330.410000 208.500000 331.590000 ;
      RECT 166.500000 330.410000 199.500000 331.590000 ;
      RECT 157.500000 330.410000 158.500000 331.590000 ;
      RECT 116.500000 330.410000 149.500000 331.590000 ;
      RECT 107.500000 330.410000 108.500000 331.590000 ;
      RECT 66.500000 330.410000 99.500000 331.590000 ;
      RECT 57.500000 330.410000 58.500000 331.590000 ;
      RECT 29.500000 330.410000 49.500000 331.590000 ;
      RECT 15.500000 330.410000 16.500000 331.590000 ;
      RECT 1157.500000 329.590000 1170.500000 330.410000 ;
      RECT 1107.500000 329.590000 1149.500000 330.410000 ;
      RECT 1057.500000 329.590000 1099.500000 330.410000 ;
      RECT 1007.500000 329.590000 1049.500000 330.410000 ;
      RECT 957.500000 329.590000 999.500000 330.410000 ;
      RECT 907.500000 329.590000 949.500000 330.410000 ;
      RECT 857.500000 329.590000 899.500000 330.410000 ;
      RECT 807.500000 329.590000 849.500000 330.410000 ;
      RECT 757.500000 329.590000 799.500000 330.410000 ;
      RECT 707.500000 329.590000 749.500000 330.410000 ;
      RECT 657.500000 329.590000 699.500000 330.410000 ;
      RECT 607.500000 329.590000 649.500000 330.410000 ;
      RECT 557.500000 329.590000 599.500000 330.410000 ;
      RECT 507.500000 329.590000 549.500000 330.410000 ;
      RECT 457.500000 329.590000 499.500000 330.410000 ;
      RECT 407.500000 329.590000 449.500000 330.410000 ;
      RECT 357.500000 329.590000 399.500000 330.410000 ;
      RECT 307.500000 329.590000 349.500000 330.410000 ;
      RECT 257.500000 329.590000 299.500000 330.410000 ;
      RECT 207.500000 329.590000 249.500000 330.410000 ;
      RECT 157.500000 329.590000 199.500000 330.410000 ;
      RECT 107.500000 329.590000 149.500000 330.410000 ;
      RECT 57.500000 329.590000 99.500000 330.410000 ;
      RECT 15.500000 329.590000 49.500000 330.410000 ;
      RECT 1183.500000 328.410000 1186.000000 331.590000 ;
      RECT 1169.500000 328.410000 1170.500000 329.590000 ;
      RECT 1116.500000 328.410000 1149.500000 329.590000 ;
      RECT 1107.500000 328.410000 1108.500000 329.590000 ;
      RECT 1066.500000 328.410000 1099.500000 329.590000 ;
      RECT 1057.500000 328.410000 1058.500000 329.590000 ;
      RECT 1016.500000 328.410000 1049.500000 329.590000 ;
      RECT 1007.500000 328.410000 1008.500000 329.590000 ;
      RECT 966.500000 328.410000 999.500000 329.590000 ;
      RECT 957.500000 328.410000 958.500000 329.590000 ;
      RECT 916.500000 328.410000 949.500000 329.590000 ;
      RECT 907.500000 328.410000 908.500000 329.590000 ;
      RECT 866.500000 328.410000 899.500000 329.590000 ;
      RECT 857.500000 328.410000 858.500000 329.590000 ;
      RECT 816.500000 328.410000 849.500000 329.590000 ;
      RECT 807.500000 328.410000 808.500000 329.590000 ;
      RECT 766.500000 328.410000 799.500000 329.590000 ;
      RECT 757.500000 328.410000 758.500000 329.590000 ;
      RECT 716.500000 328.410000 749.500000 329.590000 ;
      RECT 707.500000 328.410000 708.500000 329.590000 ;
      RECT 666.500000 328.410000 699.500000 329.590000 ;
      RECT 657.500000 328.410000 658.500000 329.590000 ;
      RECT 616.500000 328.410000 649.500000 329.590000 ;
      RECT 607.500000 328.410000 608.500000 329.590000 ;
      RECT 566.500000 328.410000 599.500000 329.590000 ;
      RECT 557.500000 328.410000 558.500000 329.590000 ;
      RECT 516.500000 328.410000 549.500000 329.590000 ;
      RECT 507.500000 328.410000 508.500000 329.590000 ;
      RECT 466.500000 328.410000 499.500000 329.590000 ;
      RECT 457.500000 328.410000 458.500000 329.590000 ;
      RECT 416.500000 328.410000 449.500000 329.590000 ;
      RECT 407.500000 328.410000 408.500000 329.590000 ;
      RECT 366.500000 328.410000 399.500000 329.590000 ;
      RECT 357.500000 328.410000 358.500000 329.590000 ;
      RECT 316.500000 328.410000 349.500000 329.590000 ;
      RECT 307.500000 328.410000 308.500000 329.590000 ;
      RECT 266.500000 328.410000 299.500000 329.590000 ;
      RECT 257.500000 328.410000 258.500000 329.590000 ;
      RECT 216.500000 328.410000 249.500000 329.590000 ;
      RECT 207.500000 328.410000 208.500000 329.590000 ;
      RECT 166.500000 328.410000 199.500000 329.590000 ;
      RECT 157.500000 328.410000 158.500000 329.590000 ;
      RECT 116.500000 328.410000 149.500000 329.590000 ;
      RECT 107.500000 328.410000 108.500000 329.590000 ;
      RECT 66.500000 328.410000 99.500000 329.590000 ;
      RECT 57.500000 328.410000 58.500000 329.590000 ;
      RECT 29.500000 328.410000 49.500000 329.590000 ;
      RECT 15.500000 328.410000 16.500000 329.590000 ;
      RECT 0.000000 328.410000 2.500000 331.590000 ;
      RECT 1169.500000 327.590000 1186.000000 328.410000 ;
      RECT 1116.500000 327.590000 1156.500000 328.410000 ;
      RECT 1066.500000 327.590000 1108.500000 328.410000 ;
      RECT 1016.500000 327.590000 1058.500000 328.410000 ;
      RECT 966.500000 327.590000 1008.500000 328.410000 ;
      RECT 916.500000 327.590000 958.500000 328.410000 ;
      RECT 866.500000 327.590000 908.500000 328.410000 ;
      RECT 816.500000 327.590000 858.500000 328.410000 ;
      RECT 766.500000 327.590000 808.500000 328.410000 ;
      RECT 716.500000 327.590000 758.500000 328.410000 ;
      RECT 666.500000 327.590000 708.500000 328.410000 ;
      RECT 616.500000 327.590000 658.500000 328.410000 ;
      RECT 566.500000 327.590000 608.500000 328.410000 ;
      RECT 516.500000 327.590000 558.500000 328.410000 ;
      RECT 466.500000 327.590000 508.500000 328.410000 ;
      RECT 416.500000 327.590000 458.500000 328.410000 ;
      RECT 366.500000 327.590000 408.500000 328.410000 ;
      RECT 316.500000 327.590000 358.500000 328.410000 ;
      RECT 266.500000 327.590000 308.500000 328.410000 ;
      RECT 216.500000 327.590000 258.500000 328.410000 ;
      RECT 166.500000 327.590000 208.500000 328.410000 ;
      RECT 116.500000 327.590000 158.500000 328.410000 ;
      RECT 66.500000 327.590000 108.500000 328.410000 ;
      RECT 29.500000 327.590000 58.500000 328.410000 ;
      RECT 0.000000 327.590000 16.500000 328.410000 ;
      RECT 1169.500000 326.410000 1170.500000 327.590000 ;
      RECT 1116.500000 326.410000 1149.500000 327.590000 ;
      RECT 1107.500000 326.410000 1108.500000 327.590000 ;
      RECT 1066.500000 326.410000 1099.500000 327.590000 ;
      RECT 1057.500000 326.410000 1058.500000 327.590000 ;
      RECT 1016.500000 326.410000 1049.500000 327.590000 ;
      RECT 1007.500000 326.410000 1008.500000 327.590000 ;
      RECT 966.500000 326.410000 999.500000 327.590000 ;
      RECT 957.500000 326.410000 958.500000 327.590000 ;
      RECT 916.500000 326.410000 949.500000 327.590000 ;
      RECT 907.500000 326.410000 908.500000 327.590000 ;
      RECT 866.500000 326.410000 899.500000 327.590000 ;
      RECT 857.500000 326.410000 858.500000 327.590000 ;
      RECT 816.500000 326.410000 849.500000 327.590000 ;
      RECT 807.500000 326.410000 808.500000 327.590000 ;
      RECT 766.500000 326.410000 799.500000 327.590000 ;
      RECT 757.500000 326.410000 758.500000 327.590000 ;
      RECT 716.500000 326.410000 749.500000 327.590000 ;
      RECT 707.500000 326.410000 708.500000 327.590000 ;
      RECT 666.500000 326.410000 699.500000 327.590000 ;
      RECT 657.500000 326.410000 658.500000 327.590000 ;
      RECT 616.500000 326.410000 649.500000 327.590000 ;
      RECT 607.500000 326.410000 608.500000 327.590000 ;
      RECT 566.500000 326.410000 599.500000 327.590000 ;
      RECT 557.500000 326.410000 558.500000 327.590000 ;
      RECT 516.500000 326.410000 549.500000 327.590000 ;
      RECT 507.500000 326.410000 508.500000 327.590000 ;
      RECT 466.500000 326.410000 499.500000 327.590000 ;
      RECT 457.500000 326.410000 458.500000 327.590000 ;
      RECT 416.500000 326.410000 449.500000 327.590000 ;
      RECT 407.500000 326.410000 408.500000 327.590000 ;
      RECT 366.500000 326.410000 399.500000 327.590000 ;
      RECT 357.500000 326.410000 358.500000 327.590000 ;
      RECT 316.500000 326.410000 349.500000 327.590000 ;
      RECT 307.500000 326.410000 308.500000 327.590000 ;
      RECT 266.500000 326.410000 299.500000 327.590000 ;
      RECT 257.500000 326.410000 258.500000 327.590000 ;
      RECT 216.500000 326.410000 249.500000 327.590000 ;
      RECT 207.500000 326.410000 208.500000 327.590000 ;
      RECT 166.500000 326.410000 199.500000 327.590000 ;
      RECT 157.500000 326.410000 158.500000 327.590000 ;
      RECT 116.500000 326.410000 149.500000 327.590000 ;
      RECT 107.500000 326.410000 108.500000 327.590000 ;
      RECT 66.500000 326.410000 99.500000 327.590000 ;
      RECT 57.500000 326.410000 58.500000 327.590000 ;
      RECT 29.500000 326.410000 49.500000 327.590000 ;
      RECT 15.500000 326.410000 16.500000 327.590000 ;
      RECT 1157.500000 325.590000 1170.500000 326.410000 ;
      RECT 1107.500000 325.590000 1149.500000 326.410000 ;
      RECT 1057.500000 325.590000 1099.500000 326.410000 ;
      RECT 1007.500000 325.590000 1049.500000 326.410000 ;
      RECT 957.500000 325.590000 999.500000 326.410000 ;
      RECT 907.500000 325.590000 949.500000 326.410000 ;
      RECT 857.500000 325.590000 899.500000 326.410000 ;
      RECT 807.500000 325.590000 849.500000 326.410000 ;
      RECT 757.500000 325.590000 799.500000 326.410000 ;
      RECT 707.500000 325.590000 749.500000 326.410000 ;
      RECT 657.500000 325.590000 699.500000 326.410000 ;
      RECT 607.500000 325.590000 649.500000 326.410000 ;
      RECT 557.500000 325.590000 599.500000 326.410000 ;
      RECT 507.500000 325.590000 549.500000 326.410000 ;
      RECT 457.500000 325.590000 499.500000 326.410000 ;
      RECT 407.500000 325.590000 449.500000 326.410000 ;
      RECT 357.500000 325.590000 399.500000 326.410000 ;
      RECT 307.500000 325.590000 349.500000 326.410000 ;
      RECT 257.500000 325.590000 299.500000 326.410000 ;
      RECT 207.500000 325.590000 249.500000 326.410000 ;
      RECT 157.500000 325.590000 199.500000 326.410000 ;
      RECT 107.500000 325.590000 149.500000 326.410000 ;
      RECT 57.500000 325.590000 99.500000 326.410000 ;
      RECT 15.500000 325.590000 49.500000 326.410000 ;
      RECT 1183.500000 324.410000 1186.000000 327.590000 ;
      RECT 1169.500000 324.410000 1170.500000 325.590000 ;
      RECT 1116.500000 324.410000 1149.500000 325.590000 ;
      RECT 1107.500000 324.410000 1108.500000 325.590000 ;
      RECT 1066.500000 324.410000 1099.500000 325.590000 ;
      RECT 1057.500000 324.410000 1058.500000 325.590000 ;
      RECT 1016.500000 324.410000 1049.500000 325.590000 ;
      RECT 1007.500000 324.410000 1008.500000 325.590000 ;
      RECT 966.500000 324.410000 999.500000 325.590000 ;
      RECT 957.500000 324.410000 958.500000 325.590000 ;
      RECT 916.500000 324.410000 949.500000 325.590000 ;
      RECT 907.500000 324.410000 908.500000 325.590000 ;
      RECT 866.500000 324.410000 899.500000 325.590000 ;
      RECT 857.500000 324.410000 858.500000 325.590000 ;
      RECT 816.500000 324.410000 849.500000 325.590000 ;
      RECT 807.500000 324.410000 808.500000 325.590000 ;
      RECT 766.500000 324.410000 799.500000 325.590000 ;
      RECT 757.500000 324.410000 758.500000 325.590000 ;
      RECT 716.500000 324.410000 749.500000 325.590000 ;
      RECT 707.500000 324.410000 708.500000 325.590000 ;
      RECT 666.500000 324.410000 699.500000 325.590000 ;
      RECT 657.500000 324.410000 658.500000 325.590000 ;
      RECT 616.500000 324.410000 649.500000 325.590000 ;
      RECT 607.500000 324.410000 608.500000 325.590000 ;
      RECT 566.500000 324.410000 599.500000 325.590000 ;
      RECT 557.500000 324.410000 558.500000 325.590000 ;
      RECT 516.500000 324.410000 549.500000 325.590000 ;
      RECT 507.500000 324.410000 508.500000 325.590000 ;
      RECT 466.500000 324.410000 499.500000 325.590000 ;
      RECT 457.500000 324.410000 458.500000 325.590000 ;
      RECT 416.500000 324.410000 449.500000 325.590000 ;
      RECT 407.500000 324.410000 408.500000 325.590000 ;
      RECT 366.500000 324.410000 399.500000 325.590000 ;
      RECT 357.500000 324.410000 358.500000 325.590000 ;
      RECT 316.500000 324.410000 349.500000 325.590000 ;
      RECT 307.500000 324.410000 308.500000 325.590000 ;
      RECT 266.500000 324.410000 299.500000 325.590000 ;
      RECT 257.500000 324.410000 258.500000 325.590000 ;
      RECT 216.500000 324.410000 249.500000 325.590000 ;
      RECT 207.500000 324.410000 208.500000 325.590000 ;
      RECT 166.500000 324.410000 199.500000 325.590000 ;
      RECT 157.500000 324.410000 158.500000 325.590000 ;
      RECT 116.500000 324.410000 149.500000 325.590000 ;
      RECT 107.500000 324.410000 108.500000 325.590000 ;
      RECT 66.500000 324.410000 99.500000 325.590000 ;
      RECT 57.500000 324.410000 58.500000 325.590000 ;
      RECT 29.500000 324.410000 49.500000 325.590000 ;
      RECT 15.500000 324.410000 16.500000 325.590000 ;
      RECT 0.000000 324.410000 2.500000 327.590000 ;
      RECT 1169.500000 323.590000 1186.000000 324.410000 ;
      RECT 1116.500000 323.590000 1156.500000 324.410000 ;
      RECT 1066.500000 323.590000 1108.500000 324.410000 ;
      RECT 1016.500000 323.590000 1058.500000 324.410000 ;
      RECT 966.500000 323.590000 1008.500000 324.410000 ;
      RECT 916.500000 323.590000 958.500000 324.410000 ;
      RECT 866.500000 323.590000 908.500000 324.410000 ;
      RECT 816.500000 323.590000 858.500000 324.410000 ;
      RECT 766.500000 323.590000 808.500000 324.410000 ;
      RECT 716.500000 323.590000 758.500000 324.410000 ;
      RECT 666.500000 323.590000 708.500000 324.410000 ;
      RECT 616.500000 323.590000 658.500000 324.410000 ;
      RECT 566.500000 323.590000 608.500000 324.410000 ;
      RECT 516.500000 323.590000 558.500000 324.410000 ;
      RECT 466.500000 323.590000 508.500000 324.410000 ;
      RECT 416.500000 323.590000 458.500000 324.410000 ;
      RECT 366.500000 323.590000 408.500000 324.410000 ;
      RECT 316.500000 323.590000 358.500000 324.410000 ;
      RECT 266.500000 323.590000 308.500000 324.410000 ;
      RECT 216.500000 323.590000 258.500000 324.410000 ;
      RECT 166.500000 323.590000 208.500000 324.410000 ;
      RECT 116.500000 323.590000 158.500000 324.410000 ;
      RECT 66.500000 323.590000 108.500000 324.410000 ;
      RECT 29.500000 323.590000 58.500000 324.410000 ;
      RECT 0.000000 323.590000 16.500000 324.410000 ;
      RECT 1169.500000 322.410000 1170.500000 323.590000 ;
      RECT 1116.500000 322.410000 1149.500000 323.590000 ;
      RECT 1107.500000 322.410000 1108.500000 323.590000 ;
      RECT 1066.500000 322.410000 1099.500000 323.590000 ;
      RECT 1057.500000 322.410000 1058.500000 323.590000 ;
      RECT 1016.500000 322.410000 1049.500000 323.590000 ;
      RECT 1007.500000 322.410000 1008.500000 323.590000 ;
      RECT 966.500000 322.410000 999.500000 323.590000 ;
      RECT 957.500000 322.410000 958.500000 323.590000 ;
      RECT 916.500000 322.410000 949.500000 323.590000 ;
      RECT 907.500000 322.410000 908.500000 323.590000 ;
      RECT 866.500000 322.410000 899.500000 323.590000 ;
      RECT 857.500000 322.410000 858.500000 323.590000 ;
      RECT 816.500000 322.410000 849.500000 323.590000 ;
      RECT 807.500000 322.410000 808.500000 323.590000 ;
      RECT 766.500000 322.410000 799.500000 323.590000 ;
      RECT 757.500000 322.410000 758.500000 323.590000 ;
      RECT 716.500000 322.410000 749.500000 323.590000 ;
      RECT 707.500000 322.410000 708.500000 323.590000 ;
      RECT 666.500000 322.410000 699.500000 323.590000 ;
      RECT 657.500000 322.410000 658.500000 323.590000 ;
      RECT 616.500000 322.410000 649.500000 323.590000 ;
      RECT 607.500000 322.410000 608.500000 323.590000 ;
      RECT 566.500000 322.410000 599.500000 323.590000 ;
      RECT 557.500000 322.410000 558.500000 323.590000 ;
      RECT 516.500000 322.410000 549.500000 323.590000 ;
      RECT 507.500000 322.410000 508.500000 323.590000 ;
      RECT 466.500000 322.410000 499.500000 323.590000 ;
      RECT 457.500000 322.410000 458.500000 323.590000 ;
      RECT 416.500000 322.410000 449.500000 323.590000 ;
      RECT 407.500000 322.410000 408.500000 323.590000 ;
      RECT 366.500000 322.410000 399.500000 323.590000 ;
      RECT 357.500000 322.410000 358.500000 323.590000 ;
      RECT 316.500000 322.410000 349.500000 323.590000 ;
      RECT 307.500000 322.410000 308.500000 323.590000 ;
      RECT 266.500000 322.410000 299.500000 323.590000 ;
      RECT 257.500000 322.410000 258.500000 323.590000 ;
      RECT 216.500000 322.410000 249.500000 323.590000 ;
      RECT 207.500000 322.410000 208.500000 323.590000 ;
      RECT 166.500000 322.410000 199.500000 323.590000 ;
      RECT 157.500000 322.410000 158.500000 323.590000 ;
      RECT 116.500000 322.410000 149.500000 323.590000 ;
      RECT 107.500000 322.410000 108.500000 323.590000 ;
      RECT 66.500000 322.410000 99.500000 323.590000 ;
      RECT 57.500000 322.410000 58.500000 323.590000 ;
      RECT 29.500000 322.410000 49.500000 323.590000 ;
      RECT 15.500000 322.410000 16.500000 323.590000 ;
      RECT 1157.500000 321.590000 1170.500000 322.410000 ;
      RECT 1107.500000 321.590000 1149.500000 322.410000 ;
      RECT 1057.500000 321.590000 1099.500000 322.410000 ;
      RECT 1007.500000 321.590000 1049.500000 322.410000 ;
      RECT 957.500000 321.590000 999.500000 322.410000 ;
      RECT 907.500000 321.590000 949.500000 322.410000 ;
      RECT 857.500000 321.590000 899.500000 322.410000 ;
      RECT 807.500000 321.590000 849.500000 322.410000 ;
      RECT 757.500000 321.590000 799.500000 322.410000 ;
      RECT 707.500000 321.590000 749.500000 322.410000 ;
      RECT 657.500000 321.590000 699.500000 322.410000 ;
      RECT 607.500000 321.590000 649.500000 322.410000 ;
      RECT 557.500000 321.590000 599.500000 322.410000 ;
      RECT 507.500000 321.590000 549.500000 322.410000 ;
      RECT 457.500000 321.590000 499.500000 322.410000 ;
      RECT 407.500000 321.590000 449.500000 322.410000 ;
      RECT 357.500000 321.590000 399.500000 322.410000 ;
      RECT 307.500000 321.590000 349.500000 322.410000 ;
      RECT 257.500000 321.590000 299.500000 322.410000 ;
      RECT 207.500000 321.590000 249.500000 322.410000 ;
      RECT 157.500000 321.590000 199.500000 322.410000 ;
      RECT 107.500000 321.590000 149.500000 322.410000 ;
      RECT 57.500000 321.590000 99.500000 322.410000 ;
      RECT 15.500000 321.590000 49.500000 322.410000 ;
      RECT 1183.500000 320.410000 1186.000000 323.590000 ;
      RECT 1169.500000 320.410000 1170.500000 321.590000 ;
      RECT 1116.500000 320.410000 1149.500000 321.590000 ;
      RECT 1107.500000 320.410000 1108.500000 321.590000 ;
      RECT 1066.500000 320.410000 1099.500000 321.590000 ;
      RECT 1057.500000 320.410000 1058.500000 321.590000 ;
      RECT 1016.500000 320.410000 1049.500000 321.590000 ;
      RECT 1007.500000 320.410000 1008.500000 321.590000 ;
      RECT 966.500000 320.410000 999.500000 321.590000 ;
      RECT 957.500000 320.410000 958.500000 321.590000 ;
      RECT 916.500000 320.410000 949.500000 321.590000 ;
      RECT 907.500000 320.410000 908.500000 321.590000 ;
      RECT 866.500000 320.410000 899.500000 321.590000 ;
      RECT 857.500000 320.410000 858.500000 321.590000 ;
      RECT 816.500000 320.410000 849.500000 321.590000 ;
      RECT 807.500000 320.410000 808.500000 321.590000 ;
      RECT 766.500000 320.410000 799.500000 321.590000 ;
      RECT 757.500000 320.410000 758.500000 321.590000 ;
      RECT 716.500000 320.410000 749.500000 321.590000 ;
      RECT 707.500000 320.410000 708.500000 321.590000 ;
      RECT 666.500000 320.410000 699.500000 321.590000 ;
      RECT 657.500000 320.410000 658.500000 321.590000 ;
      RECT 616.500000 320.410000 649.500000 321.590000 ;
      RECT 607.500000 320.410000 608.500000 321.590000 ;
      RECT 566.500000 320.410000 599.500000 321.590000 ;
      RECT 557.500000 320.410000 558.500000 321.590000 ;
      RECT 516.500000 320.410000 549.500000 321.590000 ;
      RECT 507.500000 320.410000 508.500000 321.590000 ;
      RECT 466.500000 320.410000 499.500000 321.590000 ;
      RECT 457.500000 320.410000 458.500000 321.590000 ;
      RECT 416.500000 320.410000 449.500000 321.590000 ;
      RECT 407.500000 320.410000 408.500000 321.590000 ;
      RECT 366.500000 320.410000 399.500000 321.590000 ;
      RECT 357.500000 320.410000 358.500000 321.590000 ;
      RECT 316.500000 320.410000 349.500000 321.590000 ;
      RECT 307.500000 320.410000 308.500000 321.590000 ;
      RECT 266.500000 320.410000 299.500000 321.590000 ;
      RECT 257.500000 320.410000 258.500000 321.590000 ;
      RECT 216.500000 320.410000 249.500000 321.590000 ;
      RECT 207.500000 320.410000 208.500000 321.590000 ;
      RECT 166.500000 320.410000 199.500000 321.590000 ;
      RECT 157.500000 320.410000 158.500000 321.590000 ;
      RECT 116.500000 320.410000 149.500000 321.590000 ;
      RECT 107.500000 320.410000 108.500000 321.590000 ;
      RECT 66.500000 320.410000 99.500000 321.590000 ;
      RECT 57.500000 320.410000 58.500000 321.590000 ;
      RECT 29.500000 320.410000 49.500000 321.590000 ;
      RECT 15.500000 320.410000 16.500000 321.590000 ;
      RECT 0.000000 320.410000 2.500000 323.590000 ;
      RECT 1169.500000 319.590000 1186.000000 320.410000 ;
      RECT 1116.500000 319.590000 1156.500000 320.410000 ;
      RECT 1066.500000 319.590000 1108.500000 320.410000 ;
      RECT 1016.500000 319.590000 1058.500000 320.410000 ;
      RECT 966.500000 319.590000 1008.500000 320.410000 ;
      RECT 916.500000 319.590000 958.500000 320.410000 ;
      RECT 866.500000 319.590000 908.500000 320.410000 ;
      RECT 816.500000 319.590000 858.500000 320.410000 ;
      RECT 766.500000 319.590000 808.500000 320.410000 ;
      RECT 716.500000 319.590000 758.500000 320.410000 ;
      RECT 666.500000 319.590000 708.500000 320.410000 ;
      RECT 616.500000 319.590000 658.500000 320.410000 ;
      RECT 566.500000 319.590000 608.500000 320.410000 ;
      RECT 516.500000 319.590000 558.500000 320.410000 ;
      RECT 466.500000 319.590000 508.500000 320.410000 ;
      RECT 366.500000 319.590000 408.500000 320.410000 ;
      RECT 316.500000 319.590000 358.500000 320.410000 ;
      RECT 266.500000 319.590000 308.500000 320.410000 ;
      RECT 216.500000 319.590000 258.500000 320.410000 ;
      RECT 166.500000 319.590000 208.500000 320.410000 ;
      RECT 116.500000 319.590000 158.500000 320.410000 ;
      RECT 66.500000 319.590000 108.500000 320.410000 ;
      RECT 29.500000 319.590000 58.500000 320.410000 ;
      RECT 0.000000 319.590000 16.500000 320.410000 ;
      RECT 1169.500000 318.410000 1170.500000 319.590000 ;
      RECT 1116.500000 318.410000 1149.500000 319.590000 ;
      RECT 1107.500000 318.410000 1108.500000 319.590000 ;
      RECT 1066.500000 318.410000 1099.500000 319.590000 ;
      RECT 1057.500000 318.410000 1058.500000 319.590000 ;
      RECT 1016.500000 318.410000 1049.500000 319.590000 ;
      RECT 1007.500000 318.410000 1008.500000 319.590000 ;
      RECT 966.500000 318.410000 999.500000 319.590000 ;
      RECT 957.500000 318.410000 958.500000 319.590000 ;
      RECT 916.500000 318.410000 949.500000 319.590000 ;
      RECT 907.500000 318.410000 908.500000 319.590000 ;
      RECT 866.500000 318.410000 899.500000 319.590000 ;
      RECT 857.500000 318.410000 858.500000 319.590000 ;
      RECT 816.500000 318.410000 849.500000 319.590000 ;
      RECT 807.500000 318.410000 808.500000 319.590000 ;
      RECT 766.500000 318.410000 799.500000 319.590000 ;
      RECT 757.500000 318.410000 758.500000 319.590000 ;
      RECT 716.500000 318.410000 749.500000 319.590000 ;
      RECT 707.500000 318.410000 708.500000 319.590000 ;
      RECT 666.500000 318.410000 699.500000 319.590000 ;
      RECT 657.500000 318.410000 658.500000 319.590000 ;
      RECT 616.500000 318.410000 649.500000 319.590000 ;
      RECT 607.500000 318.410000 608.500000 319.590000 ;
      RECT 566.500000 318.410000 599.500000 319.590000 ;
      RECT 557.500000 318.410000 558.500000 319.590000 ;
      RECT 516.500000 318.410000 549.500000 319.590000 ;
      RECT 507.500000 318.410000 508.500000 319.590000 ;
      RECT 466.500000 318.410000 499.500000 319.590000 ;
      RECT 416.500000 318.410000 458.500000 320.410000 ;
      RECT 407.500000 318.410000 408.500000 319.590000 ;
      RECT 366.500000 318.410000 399.500000 319.590000 ;
      RECT 357.500000 318.410000 358.500000 319.590000 ;
      RECT 316.500000 318.410000 349.500000 319.590000 ;
      RECT 307.500000 318.410000 308.500000 319.590000 ;
      RECT 266.500000 318.410000 299.500000 319.590000 ;
      RECT 257.500000 318.410000 258.500000 319.590000 ;
      RECT 216.500000 318.410000 249.500000 319.590000 ;
      RECT 207.500000 318.410000 208.500000 319.590000 ;
      RECT 166.500000 318.410000 199.500000 319.590000 ;
      RECT 157.500000 318.410000 158.500000 319.590000 ;
      RECT 116.500000 318.410000 149.500000 319.590000 ;
      RECT 107.500000 318.410000 108.500000 319.590000 ;
      RECT 66.500000 318.410000 99.500000 319.590000 ;
      RECT 57.500000 318.410000 58.500000 319.590000 ;
      RECT 29.500000 318.410000 49.500000 319.590000 ;
      RECT 15.500000 318.410000 16.500000 319.590000 ;
      RECT 1157.500000 317.590000 1170.500000 318.410000 ;
      RECT 1107.500000 317.590000 1149.500000 318.410000 ;
      RECT 1057.500000 317.590000 1099.500000 318.410000 ;
      RECT 1007.500000 317.590000 1049.500000 318.410000 ;
      RECT 957.500000 317.590000 999.500000 318.410000 ;
      RECT 907.500000 317.590000 949.500000 318.410000 ;
      RECT 857.500000 317.590000 899.500000 318.410000 ;
      RECT 807.500000 317.590000 849.500000 318.410000 ;
      RECT 757.500000 317.590000 799.500000 318.410000 ;
      RECT 707.500000 317.590000 749.500000 318.410000 ;
      RECT 657.500000 317.590000 699.500000 318.410000 ;
      RECT 607.500000 317.590000 649.500000 318.410000 ;
      RECT 557.500000 317.590000 599.500000 318.410000 ;
      RECT 507.500000 317.590000 549.500000 318.410000 ;
      RECT 407.500000 317.590000 499.500000 318.410000 ;
      RECT 357.500000 317.590000 399.500000 318.410000 ;
      RECT 307.500000 317.590000 349.500000 318.410000 ;
      RECT 257.500000 317.590000 299.500000 318.410000 ;
      RECT 207.500000 317.590000 249.500000 318.410000 ;
      RECT 157.500000 317.590000 199.500000 318.410000 ;
      RECT 107.500000 317.590000 149.500000 318.410000 ;
      RECT 57.500000 317.590000 99.500000 318.410000 ;
      RECT 15.500000 317.590000 49.500000 318.410000 ;
      RECT 1183.500000 316.410000 1186.000000 319.590000 ;
      RECT 1169.500000 316.410000 1170.500000 317.590000 ;
      RECT 1116.500000 316.410000 1149.500000 317.590000 ;
      RECT 1107.500000 316.410000 1108.500000 317.590000 ;
      RECT 1066.500000 316.410000 1099.500000 317.590000 ;
      RECT 1057.500000 316.410000 1058.500000 317.590000 ;
      RECT 1016.500000 316.410000 1049.500000 317.590000 ;
      RECT 1007.500000 316.410000 1008.500000 317.590000 ;
      RECT 966.500000 316.410000 999.500000 317.590000 ;
      RECT 957.500000 316.410000 958.500000 317.590000 ;
      RECT 916.500000 316.410000 949.500000 317.590000 ;
      RECT 907.500000 316.410000 908.500000 317.590000 ;
      RECT 866.500000 316.410000 899.500000 317.590000 ;
      RECT 857.500000 316.410000 858.500000 317.590000 ;
      RECT 816.500000 316.410000 849.500000 317.590000 ;
      RECT 807.500000 316.410000 808.500000 317.590000 ;
      RECT 766.500000 316.410000 799.500000 317.590000 ;
      RECT 757.500000 316.410000 758.500000 317.590000 ;
      RECT 716.500000 316.410000 749.500000 317.590000 ;
      RECT 707.500000 316.410000 708.500000 317.590000 ;
      RECT 666.500000 316.410000 699.500000 317.590000 ;
      RECT 657.500000 316.410000 658.500000 317.590000 ;
      RECT 616.500000 316.410000 649.500000 317.590000 ;
      RECT 607.500000 316.410000 608.500000 317.590000 ;
      RECT 566.500000 316.410000 599.500000 317.590000 ;
      RECT 557.500000 316.410000 558.500000 317.590000 ;
      RECT 516.500000 316.410000 549.500000 317.590000 ;
      RECT 507.500000 316.410000 508.500000 317.590000 ;
      RECT 416.500000 316.410000 499.500000 317.590000 ;
      RECT 407.500000 316.410000 408.500000 317.590000 ;
      RECT 366.500000 316.410000 399.500000 317.590000 ;
      RECT 357.500000 316.410000 358.500000 317.590000 ;
      RECT 316.500000 316.410000 349.500000 317.590000 ;
      RECT 307.500000 316.410000 308.500000 317.590000 ;
      RECT 266.500000 316.410000 299.500000 317.590000 ;
      RECT 257.500000 316.410000 258.500000 317.590000 ;
      RECT 216.500000 316.410000 249.500000 317.590000 ;
      RECT 207.500000 316.410000 208.500000 317.590000 ;
      RECT 166.500000 316.410000 199.500000 317.590000 ;
      RECT 157.500000 316.410000 158.500000 317.590000 ;
      RECT 116.500000 316.410000 149.500000 317.590000 ;
      RECT 107.500000 316.410000 108.500000 317.590000 ;
      RECT 66.500000 316.410000 99.500000 317.590000 ;
      RECT 57.500000 316.410000 58.500000 317.590000 ;
      RECT 29.500000 316.410000 49.500000 317.590000 ;
      RECT 15.500000 316.410000 16.500000 317.590000 ;
      RECT 0.000000 316.410000 2.500000 319.590000 ;
      RECT 1169.500000 315.590000 1186.000000 316.410000 ;
      RECT 1116.500000 315.590000 1156.500000 316.410000 ;
      RECT 1066.500000 315.590000 1108.500000 316.410000 ;
      RECT 1016.500000 315.590000 1058.500000 316.410000 ;
      RECT 966.500000 315.590000 1008.500000 316.410000 ;
      RECT 916.500000 315.590000 958.500000 316.410000 ;
      RECT 866.500000 315.590000 908.500000 316.410000 ;
      RECT 816.500000 315.590000 858.500000 316.410000 ;
      RECT 766.500000 315.590000 808.500000 316.410000 ;
      RECT 716.500000 315.590000 758.500000 316.410000 ;
      RECT 666.500000 315.590000 708.500000 316.410000 ;
      RECT 616.500000 315.590000 658.500000 316.410000 ;
      RECT 566.500000 315.590000 608.500000 316.410000 ;
      RECT 516.500000 315.590000 558.500000 316.410000 ;
      RECT 416.500000 315.590000 508.500000 316.410000 ;
      RECT 366.500000 315.590000 408.500000 316.410000 ;
      RECT 316.500000 315.590000 358.500000 316.410000 ;
      RECT 266.500000 315.590000 308.500000 316.410000 ;
      RECT 216.500000 315.590000 258.500000 316.410000 ;
      RECT 166.500000 315.590000 208.500000 316.410000 ;
      RECT 116.500000 315.590000 158.500000 316.410000 ;
      RECT 66.500000 315.590000 108.500000 316.410000 ;
      RECT 29.500000 315.590000 58.500000 316.410000 ;
      RECT 0.000000 315.590000 16.500000 316.410000 ;
      RECT 1169.500000 314.410000 1170.500000 315.590000 ;
      RECT 1116.500000 314.410000 1149.500000 315.590000 ;
      RECT 1107.500000 314.410000 1108.500000 315.590000 ;
      RECT 1066.500000 314.410000 1099.500000 315.590000 ;
      RECT 1057.500000 314.410000 1058.500000 315.590000 ;
      RECT 1016.500000 314.410000 1049.500000 315.590000 ;
      RECT 1007.500000 314.410000 1008.500000 315.590000 ;
      RECT 966.500000 314.410000 999.500000 315.590000 ;
      RECT 957.500000 314.410000 958.500000 315.590000 ;
      RECT 916.500000 314.410000 949.500000 315.590000 ;
      RECT 907.500000 314.410000 908.500000 315.590000 ;
      RECT 866.500000 314.410000 899.500000 315.590000 ;
      RECT 857.500000 314.410000 858.500000 315.590000 ;
      RECT 816.500000 314.410000 849.500000 315.590000 ;
      RECT 807.500000 314.410000 808.500000 315.590000 ;
      RECT 766.500000 314.410000 799.500000 315.590000 ;
      RECT 757.500000 314.410000 758.500000 315.590000 ;
      RECT 716.500000 314.410000 749.500000 315.590000 ;
      RECT 707.500000 314.410000 708.500000 315.590000 ;
      RECT 666.500000 314.410000 699.500000 315.590000 ;
      RECT 657.500000 314.410000 658.500000 315.590000 ;
      RECT 616.500000 314.410000 649.500000 315.590000 ;
      RECT 607.500000 314.410000 608.500000 315.590000 ;
      RECT 566.500000 314.410000 599.500000 315.590000 ;
      RECT 557.500000 314.410000 558.500000 315.590000 ;
      RECT 516.500000 314.410000 549.500000 315.590000 ;
      RECT 507.500000 314.410000 508.500000 315.590000 ;
      RECT 416.500000 314.410000 499.500000 315.590000 ;
      RECT 407.500000 314.410000 408.500000 315.590000 ;
      RECT 366.500000 314.410000 399.500000 315.590000 ;
      RECT 357.500000 314.410000 358.500000 315.590000 ;
      RECT 316.500000 314.410000 349.500000 315.590000 ;
      RECT 307.500000 314.410000 308.500000 315.590000 ;
      RECT 266.500000 314.410000 299.500000 315.590000 ;
      RECT 257.500000 314.410000 258.500000 315.590000 ;
      RECT 216.500000 314.410000 249.500000 315.590000 ;
      RECT 207.500000 314.410000 208.500000 315.590000 ;
      RECT 166.500000 314.410000 199.500000 315.590000 ;
      RECT 157.500000 314.410000 158.500000 315.590000 ;
      RECT 116.500000 314.410000 149.500000 315.590000 ;
      RECT 107.500000 314.410000 108.500000 315.590000 ;
      RECT 66.500000 314.410000 99.500000 315.590000 ;
      RECT 57.500000 314.410000 58.500000 315.590000 ;
      RECT 29.500000 314.410000 49.500000 315.590000 ;
      RECT 15.500000 314.410000 16.500000 315.590000 ;
      RECT 1157.500000 313.590000 1170.500000 314.410000 ;
      RECT 1107.500000 313.590000 1149.500000 314.410000 ;
      RECT 1057.500000 313.590000 1099.500000 314.410000 ;
      RECT 1007.500000 313.590000 1049.500000 314.410000 ;
      RECT 957.500000 313.590000 999.500000 314.410000 ;
      RECT 907.500000 313.590000 949.500000 314.410000 ;
      RECT 857.500000 313.590000 899.500000 314.410000 ;
      RECT 807.500000 313.590000 849.500000 314.410000 ;
      RECT 757.500000 313.590000 799.500000 314.410000 ;
      RECT 707.500000 313.590000 749.500000 314.410000 ;
      RECT 657.500000 313.590000 699.500000 314.410000 ;
      RECT 607.500000 313.590000 649.500000 314.410000 ;
      RECT 557.500000 313.590000 599.500000 314.410000 ;
      RECT 507.500000 313.590000 549.500000 314.410000 ;
      RECT 407.500000 313.590000 499.500000 314.410000 ;
      RECT 357.500000 313.590000 399.500000 314.410000 ;
      RECT 307.500000 313.590000 349.500000 314.410000 ;
      RECT 257.500000 313.590000 299.500000 314.410000 ;
      RECT 207.500000 313.590000 249.500000 314.410000 ;
      RECT 157.500000 313.590000 199.500000 314.410000 ;
      RECT 107.500000 313.590000 149.500000 314.410000 ;
      RECT 57.500000 313.590000 99.500000 314.410000 ;
      RECT 15.500000 313.590000 49.500000 314.410000 ;
      RECT 1183.500000 312.410000 1186.000000 315.590000 ;
      RECT 1169.500000 312.410000 1170.500000 313.590000 ;
      RECT 1116.500000 312.410000 1149.500000 313.590000 ;
      RECT 1107.500000 312.410000 1108.500000 313.590000 ;
      RECT 1066.500000 312.410000 1099.500000 313.590000 ;
      RECT 1057.500000 312.410000 1058.500000 313.590000 ;
      RECT 1016.500000 312.410000 1049.500000 313.590000 ;
      RECT 1007.500000 312.410000 1008.500000 313.590000 ;
      RECT 966.500000 312.410000 999.500000 313.590000 ;
      RECT 957.500000 312.410000 958.500000 313.590000 ;
      RECT 916.500000 312.410000 949.500000 313.590000 ;
      RECT 907.500000 312.410000 908.500000 313.590000 ;
      RECT 866.500000 312.410000 899.500000 313.590000 ;
      RECT 857.500000 312.410000 858.500000 313.590000 ;
      RECT 816.500000 312.410000 849.500000 313.590000 ;
      RECT 807.500000 312.410000 808.500000 313.590000 ;
      RECT 766.500000 312.410000 799.500000 313.590000 ;
      RECT 757.500000 312.410000 758.500000 313.590000 ;
      RECT 716.500000 312.410000 749.500000 313.590000 ;
      RECT 707.500000 312.410000 708.500000 313.590000 ;
      RECT 666.500000 312.410000 699.500000 313.590000 ;
      RECT 657.500000 312.410000 658.500000 313.590000 ;
      RECT 616.500000 312.410000 649.500000 313.590000 ;
      RECT 607.500000 312.410000 608.500000 313.590000 ;
      RECT 566.500000 312.410000 599.500000 313.590000 ;
      RECT 557.500000 312.410000 558.500000 313.590000 ;
      RECT 516.500000 312.410000 549.500000 313.590000 ;
      RECT 507.500000 312.410000 508.500000 313.590000 ;
      RECT 416.500000 312.410000 499.500000 313.590000 ;
      RECT 407.500000 312.410000 408.500000 313.590000 ;
      RECT 366.500000 312.410000 399.500000 313.590000 ;
      RECT 357.500000 312.410000 358.500000 313.590000 ;
      RECT 316.500000 312.410000 349.500000 313.590000 ;
      RECT 307.500000 312.410000 308.500000 313.590000 ;
      RECT 266.500000 312.410000 299.500000 313.590000 ;
      RECT 257.500000 312.410000 258.500000 313.590000 ;
      RECT 216.500000 312.410000 249.500000 313.590000 ;
      RECT 207.500000 312.410000 208.500000 313.590000 ;
      RECT 166.500000 312.410000 199.500000 313.590000 ;
      RECT 157.500000 312.410000 158.500000 313.590000 ;
      RECT 116.500000 312.410000 149.500000 313.590000 ;
      RECT 107.500000 312.410000 108.500000 313.590000 ;
      RECT 66.500000 312.410000 99.500000 313.590000 ;
      RECT 57.500000 312.410000 58.500000 313.590000 ;
      RECT 29.500000 312.410000 49.500000 313.590000 ;
      RECT 15.500000 312.410000 16.500000 313.590000 ;
      RECT 0.000000 312.410000 2.500000 315.590000 ;
      RECT 1169.500000 311.590000 1186.000000 312.410000 ;
      RECT 1116.500000 311.590000 1156.500000 312.410000 ;
      RECT 1066.500000 311.590000 1108.500000 312.410000 ;
      RECT 1016.500000 311.590000 1058.500000 312.410000 ;
      RECT 966.500000 311.590000 1008.500000 312.410000 ;
      RECT 916.500000 311.590000 958.500000 312.410000 ;
      RECT 866.500000 311.590000 908.500000 312.410000 ;
      RECT 816.500000 311.590000 858.500000 312.410000 ;
      RECT 766.500000 311.590000 808.500000 312.410000 ;
      RECT 716.500000 311.590000 758.500000 312.410000 ;
      RECT 666.500000 311.590000 708.500000 312.410000 ;
      RECT 616.500000 311.590000 658.500000 312.410000 ;
      RECT 566.500000 311.590000 608.500000 312.410000 ;
      RECT 516.500000 311.590000 558.500000 312.410000 ;
      RECT 416.500000 311.590000 508.500000 312.410000 ;
      RECT 366.500000 311.590000 408.500000 312.410000 ;
      RECT 316.500000 311.590000 358.500000 312.410000 ;
      RECT 266.500000 311.590000 308.500000 312.410000 ;
      RECT 216.500000 311.590000 258.500000 312.410000 ;
      RECT 166.500000 311.590000 208.500000 312.410000 ;
      RECT 116.500000 311.590000 158.500000 312.410000 ;
      RECT 66.500000 311.590000 108.500000 312.410000 ;
      RECT 29.500000 311.590000 58.500000 312.410000 ;
      RECT 0.000000 311.590000 16.500000 312.410000 ;
      RECT 0.000000 311.170000 2.500000 311.590000 ;
      RECT 1183.500000 311.165000 1186.000000 311.590000 ;
      RECT 1169.500000 310.410000 1170.500000 311.590000 ;
      RECT 1116.500000 310.410000 1149.500000 311.590000 ;
      RECT 1107.500000 310.410000 1108.500000 311.590000 ;
      RECT 1066.500000 310.410000 1099.500000 311.590000 ;
      RECT 1057.500000 310.410000 1058.500000 311.590000 ;
      RECT 1016.500000 310.410000 1049.500000 311.590000 ;
      RECT 1007.500000 310.410000 1008.500000 311.590000 ;
      RECT 966.500000 310.410000 999.500000 311.590000 ;
      RECT 957.500000 310.410000 958.500000 311.590000 ;
      RECT 916.500000 310.410000 949.500000 311.590000 ;
      RECT 907.500000 310.410000 908.500000 311.590000 ;
      RECT 866.500000 310.410000 899.500000 311.590000 ;
      RECT 857.500000 310.410000 858.500000 311.590000 ;
      RECT 816.500000 310.410000 849.500000 311.590000 ;
      RECT 807.500000 310.410000 808.500000 311.590000 ;
      RECT 766.500000 310.410000 799.500000 311.590000 ;
      RECT 757.500000 310.410000 758.500000 311.590000 ;
      RECT 716.500000 310.410000 749.500000 311.590000 ;
      RECT 707.500000 310.410000 708.500000 311.590000 ;
      RECT 666.500000 310.410000 699.500000 311.590000 ;
      RECT 657.500000 310.410000 658.500000 311.590000 ;
      RECT 616.500000 310.410000 649.500000 311.590000 ;
      RECT 607.500000 310.410000 608.500000 311.590000 ;
      RECT 566.500000 310.410000 599.500000 311.590000 ;
      RECT 557.500000 310.410000 558.500000 311.590000 ;
      RECT 516.500000 310.410000 549.500000 311.590000 ;
      RECT 507.500000 310.410000 508.500000 311.590000 ;
      RECT 416.500000 310.410000 499.500000 311.590000 ;
      RECT 407.500000 310.410000 408.500000 311.590000 ;
      RECT 366.500000 310.410000 399.500000 311.590000 ;
      RECT 357.500000 310.410000 358.500000 311.590000 ;
      RECT 316.500000 310.410000 349.500000 311.590000 ;
      RECT 307.500000 310.410000 308.500000 311.590000 ;
      RECT 266.500000 310.410000 299.500000 311.590000 ;
      RECT 257.500000 310.410000 258.500000 311.590000 ;
      RECT 216.500000 310.410000 249.500000 311.590000 ;
      RECT 207.500000 310.410000 208.500000 311.590000 ;
      RECT 166.500000 310.410000 199.500000 311.590000 ;
      RECT 157.500000 310.410000 158.500000 311.590000 ;
      RECT 116.500000 310.410000 149.500000 311.590000 ;
      RECT 107.500000 310.410000 108.500000 311.590000 ;
      RECT 66.500000 310.410000 99.500000 311.590000 ;
      RECT 57.500000 310.410000 58.500000 311.590000 ;
      RECT 29.500000 310.410000 49.500000 311.590000 ;
      RECT 15.500000 310.410000 16.500000 311.590000 ;
      RECT 1157.500000 309.590000 1170.500000 310.410000 ;
      RECT 1107.500000 309.590000 1149.500000 310.410000 ;
      RECT 1057.500000 309.590000 1099.500000 310.410000 ;
      RECT 1007.500000 309.590000 1049.500000 310.410000 ;
      RECT 957.500000 309.590000 999.500000 310.410000 ;
      RECT 907.500000 309.590000 949.500000 310.410000 ;
      RECT 857.500000 309.590000 899.500000 310.410000 ;
      RECT 807.500000 309.590000 849.500000 310.410000 ;
      RECT 757.500000 309.590000 799.500000 310.410000 ;
      RECT 707.500000 309.590000 749.500000 310.410000 ;
      RECT 657.500000 309.590000 699.500000 310.410000 ;
      RECT 607.500000 309.590000 649.500000 310.410000 ;
      RECT 557.500000 309.590000 599.500000 310.410000 ;
      RECT 507.500000 309.590000 549.500000 310.410000 ;
      RECT 407.500000 309.590000 499.500000 310.410000 ;
      RECT 357.500000 309.590000 399.500000 310.410000 ;
      RECT 307.500000 309.590000 349.500000 310.410000 ;
      RECT 257.500000 309.590000 299.500000 310.410000 ;
      RECT 207.500000 309.590000 249.500000 310.410000 ;
      RECT 157.500000 309.590000 199.500000 310.410000 ;
      RECT 107.500000 309.590000 149.500000 310.410000 ;
      RECT 57.500000 309.590000 99.500000 310.410000 ;
      RECT 15.500000 309.590000 49.500000 310.410000 ;
      RECT 1183.500000 308.410000 1183.980000 311.165000 ;
      RECT 1169.500000 308.410000 1170.500000 309.590000 ;
      RECT 1116.500000 308.410000 1149.500000 309.590000 ;
      RECT 1107.500000 308.410000 1108.500000 309.590000 ;
      RECT 1066.500000 308.410000 1099.500000 309.590000 ;
      RECT 1057.500000 308.410000 1058.500000 309.590000 ;
      RECT 1016.500000 308.410000 1049.500000 309.590000 ;
      RECT 1007.500000 308.410000 1008.500000 309.590000 ;
      RECT 966.500000 308.410000 999.500000 309.590000 ;
      RECT 957.500000 308.410000 958.500000 309.590000 ;
      RECT 916.500000 308.410000 949.500000 309.590000 ;
      RECT 907.500000 308.410000 908.500000 309.590000 ;
      RECT 866.500000 308.410000 899.500000 309.590000 ;
      RECT 857.500000 308.410000 858.500000 309.590000 ;
      RECT 816.500000 308.410000 849.500000 309.590000 ;
      RECT 807.500000 308.410000 808.500000 309.590000 ;
      RECT 766.500000 308.410000 799.500000 309.590000 ;
      RECT 757.500000 308.410000 758.500000 309.590000 ;
      RECT 716.500000 308.410000 749.500000 309.590000 ;
      RECT 707.500000 308.410000 708.500000 309.590000 ;
      RECT 666.500000 308.410000 699.500000 309.590000 ;
      RECT 657.500000 308.410000 658.500000 309.590000 ;
      RECT 616.500000 308.410000 649.500000 309.590000 ;
      RECT 607.500000 308.410000 608.500000 309.590000 ;
      RECT 566.500000 308.410000 599.500000 309.590000 ;
      RECT 557.500000 308.410000 558.500000 309.590000 ;
      RECT 516.500000 308.410000 549.500000 309.590000 ;
      RECT 507.500000 308.410000 508.500000 309.590000 ;
      RECT 416.500000 308.410000 499.500000 309.590000 ;
      RECT 407.500000 308.410000 408.500000 309.590000 ;
      RECT 366.500000 308.410000 399.500000 309.590000 ;
      RECT 357.500000 308.410000 358.500000 309.590000 ;
      RECT 316.500000 308.410000 349.500000 309.590000 ;
      RECT 307.500000 308.410000 308.500000 309.590000 ;
      RECT 266.500000 308.410000 299.500000 309.590000 ;
      RECT 257.500000 308.410000 258.500000 309.590000 ;
      RECT 216.500000 308.410000 249.500000 309.590000 ;
      RECT 207.500000 308.410000 208.500000 309.590000 ;
      RECT 166.500000 308.410000 199.500000 309.590000 ;
      RECT 157.500000 308.410000 158.500000 309.590000 ;
      RECT 116.500000 308.410000 149.500000 309.590000 ;
      RECT 107.500000 308.410000 108.500000 309.590000 ;
      RECT 66.500000 308.410000 99.500000 309.590000 ;
      RECT 57.500000 308.410000 58.500000 309.590000 ;
      RECT 29.500000 308.410000 49.500000 309.590000 ;
      RECT 15.500000 308.410000 16.500000 309.590000 ;
      RECT 2.020000 308.410000 2.500000 311.170000 ;
      RECT 2.020000 308.070000 16.500000 308.410000 ;
      RECT 1169.500000 308.065000 1183.980000 308.410000 ;
      RECT 1169.500000 307.590000 1186.000000 308.065000 ;
      RECT 1116.500000 307.590000 1156.500000 308.410000 ;
      RECT 1066.500000 307.590000 1108.500000 308.410000 ;
      RECT 1016.500000 307.590000 1058.500000 308.410000 ;
      RECT 966.500000 307.590000 1008.500000 308.410000 ;
      RECT 916.500000 307.590000 958.500000 308.410000 ;
      RECT 866.500000 307.590000 908.500000 308.410000 ;
      RECT 816.500000 307.590000 858.500000 308.410000 ;
      RECT 766.500000 307.590000 808.500000 308.410000 ;
      RECT 716.500000 307.590000 758.500000 308.410000 ;
      RECT 666.500000 307.590000 708.500000 308.410000 ;
      RECT 616.500000 307.590000 658.500000 308.410000 ;
      RECT 566.500000 307.590000 608.500000 308.410000 ;
      RECT 516.500000 307.590000 558.500000 308.410000 ;
      RECT 416.500000 307.590000 508.500000 308.410000 ;
      RECT 366.500000 307.590000 408.500000 308.410000 ;
      RECT 316.500000 307.590000 358.500000 308.410000 ;
      RECT 266.500000 307.590000 308.500000 308.410000 ;
      RECT 216.500000 307.590000 258.500000 308.410000 ;
      RECT 166.500000 307.590000 208.500000 308.410000 ;
      RECT 116.500000 307.590000 158.500000 308.410000 ;
      RECT 66.500000 307.590000 108.500000 308.410000 ;
      RECT 29.500000 307.590000 58.500000 308.410000 ;
      RECT 0.000000 307.590000 16.500000 308.070000 ;
      RECT 1169.500000 306.410000 1170.500000 307.590000 ;
      RECT 1116.500000 306.410000 1149.500000 307.590000 ;
      RECT 1107.500000 306.410000 1108.500000 307.590000 ;
      RECT 1066.500000 306.410000 1099.500000 307.590000 ;
      RECT 1057.500000 306.410000 1058.500000 307.590000 ;
      RECT 1016.500000 306.410000 1049.500000 307.590000 ;
      RECT 1007.500000 306.410000 1008.500000 307.590000 ;
      RECT 966.500000 306.410000 999.500000 307.590000 ;
      RECT 957.500000 306.410000 958.500000 307.590000 ;
      RECT 916.500000 306.410000 949.500000 307.590000 ;
      RECT 907.500000 306.410000 908.500000 307.590000 ;
      RECT 866.500000 306.410000 899.500000 307.590000 ;
      RECT 857.500000 306.410000 858.500000 307.590000 ;
      RECT 816.500000 306.410000 849.500000 307.590000 ;
      RECT 807.500000 306.410000 808.500000 307.590000 ;
      RECT 766.500000 306.410000 799.500000 307.590000 ;
      RECT 757.500000 306.410000 758.500000 307.590000 ;
      RECT 716.500000 306.410000 749.500000 307.590000 ;
      RECT 707.500000 306.410000 708.500000 307.590000 ;
      RECT 666.500000 306.410000 699.500000 307.590000 ;
      RECT 657.500000 306.410000 658.500000 307.590000 ;
      RECT 616.500000 306.410000 649.500000 307.590000 ;
      RECT 607.500000 306.410000 608.500000 307.590000 ;
      RECT 566.500000 306.410000 599.500000 307.590000 ;
      RECT 557.500000 306.410000 558.500000 307.590000 ;
      RECT 516.500000 306.410000 549.500000 307.590000 ;
      RECT 507.500000 306.410000 508.500000 307.590000 ;
      RECT 416.500000 306.410000 499.500000 307.590000 ;
      RECT 407.500000 306.410000 408.500000 307.590000 ;
      RECT 366.500000 306.410000 399.500000 307.590000 ;
      RECT 357.500000 306.410000 358.500000 307.590000 ;
      RECT 316.500000 306.410000 349.500000 307.590000 ;
      RECT 307.500000 306.410000 308.500000 307.590000 ;
      RECT 266.500000 306.410000 299.500000 307.590000 ;
      RECT 257.500000 306.410000 258.500000 307.590000 ;
      RECT 216.500000 306.410000 249.500000 307.590000 ;
      RECT 207.500000 306.410000 208.500000 307.590000 ;
      RECT 166.500000 306.410000 199.500000 307.590000 ;
      RECT 157.500000 306.410000 158.500000 307.590000 ;
      RECT 116.500000 306.410000 149.500000 307.590000 ;
      RECT 107.500000 306.410000 108.500000 307.590000 ;
      RECT 66.500000 306.410000 99.500000 307.590000 ;
      RECT 57.500000 306.410000 58.500000 307.590000 ;
      RECT 29.500000 306.410000 49.500000 307.590000 ;
      RECT 15.500000 306.410000 16.500000 307.590000 ;
      RECT 1157.500000 305.590000 1170.500000 306.410000 ;
      RECT 1107.500000 305.590000 1149.500000 306.410000 ;
      RECT 1057.500000 305.590000 1099.500000 306.410000 ;
      RECT 1007.500000 305.590000 1049.500000 306.410000 ;
      RECT 957.500000 305.590000 999.500000 306.410000 ;
      RECT 907.500000 305.590000 949.500000 306.410000 ;
      RECT 857.500000 305.590000 899.500000 306.410000 ;
      RECT 807.500000 305.590000 849.500000 306.410000 ;
      RECT 757.500000 305.590000 799.500000 306.410000 ;
      RECT 707.500000 305.590000 749.500000 306.410000 ;
      RECT 657.500000 305.590000 699.500000 306.410000 ;
      RECT 607.500000 305.590000 649.500000 306.410000 ;
      RECT 557.500000 305.590000 599.500000 306.410000 ;
      RECT 507.500000 305.590000 549.500000 306.410000 ;
      RECT 407.500000 305.590000 499.500000 306.410000 ;
      RECT 357.500000 305.590000 399.500000 306.410000 ;
      RECT 307.500000 305.590000 349.500000 306.410000 ;
      RECT 257.500000 305.590000 299.500000 306.410000 ;
      RECT 207.500000 305.590000 249.500000 306.410000 ;
      RECT 157.500000 305.590000 199.500000 306.410000 ;
      RECT 107.500000 305.590000 149.500000 306.410000 ;
      RECT 57.500000 305.590000 99.500000 306.410000 ;
      RECT 15.500000 305.590000 49.500000 306.410000 ;
      RECT 1183.500000 305.485000 1186.000000 307.590000 ;
      RECT 1183.500000 304.410000 1183.980000 305.485000 ;
      RECT 1169.500000 304.410000 1170.500000 305.590000 ;
      RECT 1116.500000 304.410000 1149.500000 305.590000 ;
      RECT 1107.500000 304.410000 1108.500000 305.590000 ;
      RECT 1066.500000 304.410000 1099.500000 305.590000 ;
      RECT 1057.500000 304.410000 1058.500000 305.590000 ;
      RECT 1016.500000 304.410000 1049.500000 305.590000 ;
      RECT 1007.500000 304.410000 1008.500000 305.590000 ;
      RECT 966.500000 304.410000 999.500000 305.590000 ;
      RECT 957.500000 304.410000 958.500000 305.590000 ;
      RECT 916.500000 304.410000 949.500000 305.590000 ;
      RECT 907.500000 304.410000 908.500000 305.590000 ;
      RECT 866.500000 304.410000 899.500000 305.590000 ;
      RECT 857.500000 304.410000 858.500000 305.590000 ;
      RECT 816.500000 304.410000 849.500000 305.590000 ;
      RECT 807.500000 304.410000 808.500000 305.590000 ;
      RECT 766.500000 304.410000 799.500000 305.590000 ;
      RECT 757.500000 304.410000 758.500000 305.590000 ;
      RECT 716.500000 304.410000 749.500000 305.590000 ;
      RECT 707.500000 304.410000 708.500000 305.590000 ;
      RECT 666.500000 304.410000 699.500000 305.590000 ;
      RECT 657.500000 304.410000 658.500000 305.590000 ;
      RECT 616.500000 304.410000 649.500000 305.590000 ;
      RECT 607.500000 304.410000 608.500000 305.590000 ;
      RECT 566.500000 304.410000 599.500000 305.590000 ;
      RECT 557.500000 304.410000 558.500000 305.590000 ;
      RECT 516.500000 304.410000 549.500000 305.590000 ;
      RECT 507.500000 304.410000 508.500000 305.590000 ;
      RECT 416.500000 304.410000 499.500000 305.590000 ;
      RECT 407.500000 304.410000 408.500000 305.590000 ;
      RECT 366.500000 304.410000 399.500000 305.590000 ;
      RECT 357.500000 304.410000 358.500000 305.590000 ;
      RECT 316.500000 304.410000 349.500000 305.590000 ;
      RECT 307.500000 304.410000 308.500000 305.590000 ;
      RECT 266.500000 304.410000 299.500000 305.590000 ;
      RECT 257.500000 304.410000 258.500000 305.590000 ;
      RECT 216.500000 304.410000 249.500000 305.590000 ;
      RECT 207.500000 304.410000 208.500000 305.590000 ;
      RECT 166.500000 304.410000 199.500000 305.590000 ;
      RECT 157.500000 304.410000 158.500000 305.590000 ;
      RECT 116.500000 304.410000 149.500000 305.590000 ;
      RECT 107.500000 304.410000 108.500000 305.590000 ;
      RECT 66.500000 304.410000 99.500000 305.590000 ;
      RECT 57.500000 304.410000 58.500000 305.590000 ;
      RECT 29.500000 304.410000 49.500000 305.590000 ;
      RECT 15.500000 304.410000 16.500000 305.590000 ;
      RECT 0.000000 304.410000 2.500000 307.590000 ;
      RECT 1169.500000 303.590000 1183.980000 304.410000 ;
      RECT 1116.500000 303.590000 1156.500000 304.410000 ;
      RECT 1066.500000 303.590000 1108.500000 304.410000 ;
      RECT 1016.500000 303.590000 1058.500000 304.410000 ;
      RECT 966.500000 303.590000 1008.500000 304.410000 ;
      RECT 916.500000 303.590000 958.500000 304.410000 ;
      RECT 866.500000 303.590000 908.500000 304.410000 ;
      RECT 816.500000 303.590000 858.500000 304.410000 ;
      RECT 766.500000 303.590000 808.500000 304.410000 ;
      RECT 716.500000 303.590000 758.500000 304.410000 ;
      RECT 666.500000 303.590000 708.500000 304.410000 ;
      RECT 616.500000 303.590000 658.500000 304.410000 ;
      RECT 566.500000 303.590000 608.500000 304.410000 ;
      RECT 516.500000 303.590000 558.500000 304.410000 ;
      RECT 416.500000 303.590000 508.500000 304.410000 ;
      RECT 366.500000 303.590000 408.500000 304.410000 ;
      RECT 316.500000 303.590000 358.500000 304.410000 ;
      RECT 266.500000 303.590000 308.500000 304.410000 ;
      RECT 216.500000 303.590000 258.500000 304.410000 ;
      RECT 166.500000 303.590000 208.500000 304.410000 ;
      RECT 116.500000 303.590000 158.500000 304.410000 ;
      RECT 66.500000 303.590000 108.500000 304.410000 ;
      RECT 29.500000 303.590000 58.500000 304.410000 ;
      RECT 0.000000 303.590000 16.500000 304.410000 ;
      RECT 1169.500000 302.410000 1170.500000 303.590000 ;
      RECT 1116.500000 302.410000 1149.500000 303.590000 ;
      RECT 1107.500000 302.410000 1108.500000 303.590000 ;
      RECT 1066.500000 302.410000 1099.500000 303.590000 ;
      RECT 1057.500000 302.410000 1058.500000 303.590000 ;
      RECT 1016.500000 302.410000 1049.500000 303.590000 ;
      RECT 1007.500000 302.410000 1008.500000 303.590000 ;
      RECT 966.500000 302.410000 999.500000 303.590000 ;
      RECT 957.500000 302.410000 958.500000 303.590000 ;
      RECT 916.500000 302.410000 949.500000 303.590000 ;
      RECT 907.500000 302.410000 908.500000 303.590000 ;
      RECT 866.500000 302.410000 899.500000 303.590000 ;
      RECT 857.500000 302.410000 858.500000 303.590000 ;
      RECT 816.500000 302.410000 849.500000 303.590000 ;
      RECT 807.500000 302.410000 808.500000 303.590000 ;
      RECT 766.500000 302.410000 799.500000 303.590000 ;
      RECT 757.500000 302.410000 758.500000 303.590000 ;
      RECT 716.500000 302.410000 749.500000 303.590000 ;
      RECT 707.500000 302.410000 708.500000 303.590000 ;
      RECT 666.500000 302.410000 699.500000 303.590000 ;
      RECT 657.500000 302.410000 658.500000 303.590000 ;
      RECT 616.500000 302.410000 649.500000 303.590000 ;
      RECT 607.500000 302.410000 608.500000 303.590000 ;
      RECT 566.500000 302.410000 599.500000 303.590000 ;
      RECT 557.500000 302.410000 558.500000 303.590000 ;
      RECT 516.500000 302.410000 549.500000 303.590000 ;
      RECT 507.500000 302.410000 508.500000 303.590000 ;
      RECT 416.500000 302.410000 499.500000 303.590000 ;
      RECT 407.500000 302.410000 408.500000 303.590000 ;
      RECT 366.500000 302.410000 399.500000 303.590000 ;
      RECT 357.500000 302.410000 358.500000 303.590000 ;
      RECT 316.500000 302.410000 349.500000 303.590000 ;
      RECT 307.500000 302.410000 308.500000 303.590000 ;
      RECT 266.500000 302.410000 299.500000 303.590000 ;
      RECT 257.500000 302.410000 258.500000 303.590000 ;
      RECT 216.500000 302.410000 249.500000 303.590000 ;
      RECT 207.500000 302.410000 208.500000 303.590000 ;
      RECT 166.500000 302.410000 199.500000 303.590000 ;
      RECT 157.500000 302.410000 158.500000 303.590000 ;
      RECT 116.500000 302.410000 149.500000 303.590000 ;
      RECT 107.500000 302.410000 108.500000 303.590000 ;
      RECT 66.500000 302.410000 99.500000 303.590000 ;
      RECT 57.500000 302.410000 58.500000 303.590000 ;
      RECT 29.500000 302.410000 49.500000 303.590000 ;
      RECT 15.500000 302.410000 16.500000 303.590000 ;
      RECT 1183.500000 302.385000 1183.980000 303.590000 ;
      RECT 1157.500000 301.590000 1170.500000 302.410000 ;
      RECT 1107.500000 301.590000 1149.500000 302.410000 ;
      RECT 1057.500000 301.590000 1099.500000 302.410000 ;
      RECT 1007.500000 301.590000 1049.500000 302.410000 ;
      RECT 957.500000 301.590000 999.500000 302.410000 ;
      RECT 907.500000 301.590000 949.500000 302.410000 ;
      RECT 857.500000 301.590000 899.500000 302.410000 ;
      RECT 807.500000 301.590000 849.500000 302.410000 ;
      RECT 757.500000 301.590000 799.500000 302.410000 ;
      RECT 707.500000 301.590000 749.500000 302.410000 ;
      RECT 657.500000 301.590000 699.500000 302.410000 ;
      RECT 607.500000 301.590000 649.500000 302.410000 ;
      RECT 557.500000 301.590000 599.500000 302.410000 ;
      RECT 507.500000 301.590000 549.500000 302.410000 ;
      RECT 407.500000 301.590000 499.500000 302.410000 ;
      RECT 357.500000 301.590000 399.500000 302.410000 ;
      RECT 307.500000 301.590000 349.500000 302.410000 ;
      RECT 257.500000 301.590000 299.500000 302.410000 ;
      RECT 207.500000 301.590000 249.500000 302.410000 ;
      RECT 157.500000 301.590000 199.500000 302.410000 ;
      RECT 107.500000 301.590000 149.500000 302.410000 ;
      RECT 57.500000 301.590000 99.500000 302.410000 ;
      RECT 15.500000 301.590000 49.500000 302.410000 ;
      RECT 1183.500000 301.525000 1186.000000 302.385000 ;
      RECT 0.000000 300.575000 2.500000 303.590000 ;
      RECT 1183.500000 300.410000 1183.980000 301.525000 ;
      RECT 1169.500000 300.410000 1170.500000 301.590000 ;
      RECT 1116.500000 300.410000 1149.500000 301.590000 ;
      RECT 1107.500000 300.410000 1108.500000 301.590000 ;
      RECT 1066.500000 300.410000 1099.500000 301.590000 ;
      RECT 1057.500000 300.410000 1058.500000 301.590000 ;
      RECT 1016.500000 300.410000 1049.500000 301.590000 ;
      RECT 1007.500000 300.410000 1008.500000 301.590000 ;
      RECT 966.500000 300.410000 999.500000 301.590000 ;
      RECT 957.500000 300.410000 958.500000 301.590000 ;
      RECT 916.500000 300.410000 949.500000 301.590000 ;
      RECT 907.500000 300.410000 908.500000 301.590000 ;
      RECT 866.500000 300.410000 899.500000 301.590000 ;
      RECT 857.500000 300.410000 858.500000 301.590000 ;
      RECT 816.500000 300.410000 849.500000 301.590000 ;
      RECT 807.500000 300.410000 808.500000 301.590000 ;
      RECT 766.500000 300.410000 799.500000 301.590000 ;
      RECT 757.500000 300.410000 758.500000 301.590000 ;
      RECT 716.500000 300.410000 749.500000 301.590000 ;
      RECT 707.500000 300.410000 708.500000 301.590000 ;
      RECT 666.500000 300.410000 699.500000 301.590000 ;
      RECT 657.500000 300.410000 658.500000 301.590000 ;
      RECT 616.500000 300.410000 649.500000 301.590000 ;
      RECT 607.500000 300.410000 608.500000 301.590000 ;
      RECT 566.500000 300.410000 599.500000 301.590000 ;
      RECT 557.500000 300.410000 558.500000 301.590000 ;
      RECT 516.500000 300.410000 549.500000 301.590000 ;
      RECT 507.500000 300.410000 508.500000 301.590000 ;
      RECT 416.500000 300.410000 499.500000 301.590000 ;
      RECT 407.500000 300.410000 408.500000 301.590000 ;
      RECT 366.500000 300.410000 399.500000 301.590000 ;
      RECT 357.500000 300.410000 358.500000 301.590000 ;
      RECT 316.500000 300.410000 349.500000 301.590000 ;
      RECT 307.500000 300.410000 308.500000 301.590000 ;
      RECT 266.500000 300.410000 299.500000 301.590000 ;
      RECT 257.500000 300.410000 258.500000 301.590000 ;
      RECT 216.500000 300.410000 249.500000 301.590000 ;
      RECT 207.500000 300.410000 208.500000 301.590000 ;
      RECT 166.500000 300.410000 199.500000 301.590000 ;
      RECT 157.500000 300.410000 158.500000 301.590000 ;
      RECT 116.500000 300.410000 149.500000 301.590000 ;
      RECT 107.500000 300.410000 108.500000 301.590000 ;
      RECT 66.500000 300.410000 99.500000 301.590000 ;
      RECT 57.500000 300.410000 58.500000 301.590000 ;
      RECT 29.500000 300.410000 49.500000 301.590000 ;
      RECT 15.500000 300.410000 16.500000 301.590000 ;
      RECT 2.020000 300.410000 2.500000 300.575000 ;
      RECT 1169.500000 299.590000 1183.980000 300.410000 ;
      RECT 1116.500000 299.590000 1156.500000 300.410000 ;
      RECT 1066.500000 299.590000 1108.500000 300.410000 ;
      RECT 1016.500000 299.590000 1058.500000 300.410000 ;
      RECT 966.500000 299.590000 1008.500000 300.410000 ;
      RECT 916.500000 299.590000 958.500000 300.410000 ;
      RECT 866.500000 299.590000 908.500000 300.410000 ;
      RECT 816.500000 299.590000 858.500000 300.410000 ;
      RECT 766.500000 299.590000 808.500000 300.410000 ;
      RECT 716.500000 299.590000 758.500000 300.410000 ;
      RECT 666.500000 299.590000 708.500000 300.410000 ;
      RECT 616.500000 299.590000 658.500000 300.410000 ;
      RECT 566.500000 299.590000 608.500000 300.410000 ;
      RECT 516.500000 299.590000 558.500000 300.410000 ;
      RECT 416.500000 299.590000 508.500000 300.410000 ;
      RECT 366.500000 299.590000 408.500000 300.410000 ;
      RECT 316.500000 299.590000 358.500000 300.410000 ;
      RECT 266.500000 299.590000 308.500000 300.410000 ;
      RECT 216.500000 299.590000 258.500000 300.410000 ;
      RECT 166.500000 299.590000 208.500000 300.410000 ;
      RECT 116.500000 299.590000 158.500000 300.410000 ;
      RECT 66.500000 299.590000 108.500000 300.410000 ;
      RECT 29.500000 299.590000 58.500000 300.410000 ;
      RECT 2.020000 299.590000 16.500000 300.410000 ;
      RECT 1183.500000 298.425000 1183.980000 299.590000 ;
      RECT 1169.500000 298.410000 1170.500000 299.590000 ;
      RECT 1116.500000 298.410000 1149.500000 299.590000 ;
      RECT 1107.500000 298.410000 1108.500000 299.590000 ;
      RECT 1066.500000 298.410000 1099.500000 299.590000 ;
      RECT 1057.500000 298.410000 1058.500000 299.590000 ;
      RECT 1016.500000 298.410000 1049.500000 299.590000 ;
      RECT 1007.500000 298.410000 1008.500000 299.590000 ;
      RECT 966.500000 298.410000 999.500000 299.590000 ;
      RECT 957.500000 298.410000 958.500000 299.590000 ;
      RECT 916.500000 298.410000 949.500000 299.590000 ;
      RECT 907.500000 298.410000 908.500000 299.590000 ;
      RECT 866.500000 298.410000 899.500000 299.590000 ;
      RECT 857.500000 298.410000 858.500000 299.590000 ;
      RECT 816.500000 298.410000 849.500000 299.590000 ;
      RECT 807.500000 298.410000 808.500000 299.590000 ;
      RECT 766.500000 298.410000 799.500000 299.590000 ;
      RECT 757.500000 298.410000 758.500000 299.590000 ;
      RECT 716.500000 298.410000 749.500000 299.590000 ;
      RECT 707.500000 298.410000 708.500000 299.590000 ;
      RECT 666.500000 298.410000 699.500000 299.590000 ;
      RECT 657.500000 298.410000 658.500000 299.590000 ;
      RECT 616.500000 298.410000 649.500000 299.590000 ;
      RECT 607.500000 298.410000 608.500000 299.590000 ;
      RECT 566.500000 298.410000 599.500000 299.590000 ;
      RECT 557.500000 298.410000 558.500000 299.590000 ;
      RECT 516.500000 298.410000 549.500000 299.590000 ;
      RECT 507.500000 298.410000 508.500000 299.590000 ;
      RECT 416.500000 298.410000 449.500000 299.590000 ;
      RECT 407.500000 298.410000 408.500000 299.590000 ;
      RECT 366.500000 298.410000 399.500000 299.590000 ;
      RECT 357.500000 298.410000 358.500000 299.590000 ;
      RECT 316.500000 298.410000 349.500000 299.590000 ;
      RECT 307.500000 298.410000 308.500000 299.590000 ;
      RECT 266.500000 298.410000 299.500000 299.590000 ;
      RECT 257.500000 298.410000 258.500000 299.590000 ;
      RECT 216.500000 298.410000 249.500000 299.590000 ;
      RECT 207.500000 298.410000 208.500000 299.590000 ;
      RECT 166.500000 298.410000 199.500000 299.590000 ;
      RECT 157.500000 298.410000 158.500000 299.590000 ;
      RECT 116.500000 298.410000 149.500000 299.590000 ;
      RECT 107.500000 298.410000 108.500000 299.590000 ;
      RECT 66.500000 298.410000 99.500000 299.590000 ;
      RECT 57.500000 298.410000 58.500000 299.590000 ;
      RECT 29.500000 298.410000 49.500000 299.590000 ;
      RECT 15.500000 298.410000 16.500000 299.590000 ;
      RECT 1157.500000 297.590000 1170.500000 298.410000 ;
      RECT 1107.500000 297.590000 1149.500000 298.410000 ;
      RECT 1057.500000 297.590000 1099.500000 298.410000 ;
      RECT 1007.500000 297.590000 1049.500000 298.410000 ;
      RECT 957.500000 297.590000 999.500000 298.410000 ;
      RECT 907.500000 297.590000 949.500000 298.410000 ;
      RECT 857.500000 297.590000 899.500000 298.410000 ;
      RECT 807.500000 297.590000 849.500000 298.410000 ;
      RECT 757.500000 297.590000 799.500000 298.410000 ;
      RECT 707.500000 297.590000 749.500000 298.410000 ;
      RECT 657.500000 297.590000 699.500000 298.410000 ;
      RECT 607.500000 297.590000 649.500000 298.410000 ;
      RECT 557.500000 297.590000 599.500000 298.410000 ;
      RECT 507.500000 297.590000 549.500000 298.410000 ;
      RECT 457.500000 297.590000 499.500000 299.590000 ;
      RECT 407.500000 297.590000 449.500000 298.410000 ;
      RECT 357.500000 297.590000 399.500000 298.410000 ;
      RECT 307.500000 297.590000 349.500000 298.410000 ;
      RECT 257.500000 297.590000 299.500000 298.410000 ;
      RECT 207.500000 297.590000 249.500000 298.410000 ;
      RECT 157.500000 297.590000 199.500000 298.410000 ;
      RECT 107.500000 297.590000 149.500000 298.410000 ;
      RECT 57.500000 297.590000 99.500000 298.410000 ;
      RECT 15.500000 297.590000 49.500000 298.410000 ;
      RECT 2.020000 297.475000 2.500000 299.590000 ;
      RECT 0.000000 296.615000 2.500000 297.475000 ;
      RECT 1183.500000 296.410000 1186.000000 298.425000 ;
      RECT 1169.500000 296.410000 1170.500000 297.590000 ;
      RECT 1116.500000 296.410000 1149.500000 297.590000 ;
      RECT 1107.500000 296.410000 1108.500000 297.590000 ;
      RECT 1066.500000 296.410000 1099.500000 297.590000 ;
      RECT 1057.500000 296.410000 1058.500000 297.590000 ;
      RECT 1016.500000 296.410000 1049.500000 297.590000 ;
      RECT 1007.500000 296.410000 1008.500000 297.590000 ;
      RECT 966.500000 296.410000 999.500000 297.590000 ;
      RECT 957.500000 296.410000 958.500000 297.590000 ;
      RECT 916.500000 296.410000 949.500000 297.590000 ;
      RECT 907.500000 296.410000 908.500000 297.590000 ;
      RECT 866.500000 296.410000 899.500000 297.590000 ;
      RECT 857.500000 296.410000 858.500000 297.590000 ;
      RECT 816.500000 296.410000 849.500000 297.590000 ;
      RECT 807.500000 296.410000 808.500000 297.590000 ;
      RECT 766.500000 296.410000 799.500000 297.590000 ;
      RECT 757.500000 296.410000 758.500000 297.590000 ;
      RECT 716.500000 296.410000 749.500000 297.590000 ;
      RECT 707.500000 296.410000 708.500000 297.590000 ;
      RECT 666.500000 296.410000 699.500000 297.590000 ;
      RECT 657.500000 296.410000 658.500000 297.590000 ;
      RECT 616.500000 296.410000 649.500000 297.590000 ;
      RECT 607.500000 296.410000 608.500000 297.590000 ;
      RECT 566.500000 296.410000 599.500000 297.590000 ;
      RECT 557.500000 296.410000 558.500000 297.590000 ;
      RECT 516.500000 296.410000 549.500000 297.590000 ;
      RECT 507.500000 296.410000 508.500000 297.590000 ;
      RECT 466.500000 296.410000 499.500000 297.590000 ;
      RECT 457.500000 296.410000 458.500000 297.590000 ;
      RECT 416.500000 296.410000 449.500000 297.590000 ;
      RECT 407.500000 296.410000 408.500000 297.590000 ;
      RECT 366.500000 296.410000 399.500000 297.590000 ;
      RECT 357.500000 296.410000 358.500000 297.590000 ;
      RECT 316.500000 296.410000 349.500000 297.590000 ;
      RECT 307.500000 296.410000 308.500000 297.590000 ;
      RECT 266.500000 296.410000 299.500000 297.590000 ;
      RECT 257.500000 296.410000 258.500000 297.590000 ;
      RECT 216.500000 296.410000 249.500000 297.590000 ;
      RECT 207.500000 296.410000 208.500000 297.590000 ;
      RECT 166.500000 296.410000 199.500000 297.590000 ;
      RECT 157.500000 296.410000 158.500000 297.590000 ;
      RECT 116.500000 296.410000 149.500000 297.590000 ;
      RECT 107.500000 296.410000 108.500000 297.590000 ;
      RECT 66.500000 296.410000 99.500000 297.590000 ;
      RECT 57.500000 296.410000 58.500000 297.590000 ;
      RECT 29.500000 296.410000 49.500000 297.590000 ;
      RECT 15.500000 296.410000 16.500000 297.590000 ;
      RECT 2.020000 296.410000 2.500000 296.615000 ;
      RECT 1169.500000 295.590000 1186.000000 296.410000 ;
      RECT 1116.500000 295.590000 1156.500000 296.410000 ;
      RECT 1066.500000 295.590000 1108.500000 296.410000 ;
      RECT 1016.500000 295.590000 1058.500000 296.410000 ;
      RECT 966.500000 295.590000 1008.500000 296.410000 ;
      RECT 916.500000 295.590000 958.500000 296.410000 ;
      RECT 866.500000 295.590000 908.500000 296.410000 ;
      RECT 816.500000 295.590000 858.500000 296.410000 ;
      RECT 766.500000 295.590000 808.500000 296.410000 ;
      RECT 716.500000 295.590000 758.500000 296.410000 ;
      RECT 666.500000 295.590000 708.500000 296.410000 ;
      RECT 616.500000 295.590000 658.500000 296.410000 ;
      RECT 566.500000 295.590000 608.500000 296.410000 ;
      RECT 516.500000 295.590000 558.500000 296.410000 ;
      RECT 466.500000 295.590000 508.500000 296.410000 ;
      RECT 416.500000 295.590000 458.500000 296.410000 ;
      RECT 366.500000 295.590000 408.500000 296.410000 ;
      RECT 316.500000 295.590000 358.500000 296.410000 ;
      RECT 266.500000 295.590000 308.500000 296.410000 ;
      RECT 216.500000 295.590000 258.500000 296.410000 ;
      RECT 166.500000 295.590000 208.500000 296.410000 ;
      RECT 116.500000 295.590000 158.500000 296.410000 ;
      RECT 66.500000 295.590000 108.500000 296.410000 ;
      RECT 29.500000 295.590000 58.500000 296.410000 ;
      RECT 2.020000 295.590000 16.500000 296.410000 ;
      RECT 1169.500000 294.410000 1170.500000 295.590000 ;
      RECT 1116.500000 294.410000 1149.500000 295.590000 ;
      RECT 1107.500000 294.410000 1108.500000 295.590000 ;
      RECT 1066.500000 294.410000 1099.500000 295.590000 ;
      RECT 1057.500000 294.410000 1058.500000 295.590000 ;
      RECT 1016.500000 294.410000 1049.500000 295.590000 ;
      RECT 1007.500000 294.410000 1008.500000 295.590000 ;
      RECT 966.500000 294.410000 999.500000 295.590000 ;
      RECT 957.500000 294.410000 958.500000 295.590000 ;
      RECT 916.500000 294.410000 949.500000 295.590000 ;
      RECT 907.500000 294.410000 908.500000 295.590000 ;
      RECT 866.500000 294.410000 899.500000 295.590000 ;
      RECT 857.500000 294.410000 858.500000 295.590000 ;
      RECT 816.500000 294.410000 849.500000 295.590000 ;
      RECT 807.500000 294.410000 808.500000 295.590000 ;
      RECT 766.500000 294.410000 799.500000 295.590000 ;
      RECT 757.500000 294.410000 758.500000 295.590000 ;
      RECT 716.500000 294.410000 749.500000 295.590000 ;
      RECT 707.500000 294.410000 708.500000 295.590000 ;
      RECT 666.500000 294.410000 699.500000 295.590000 ;
      RECT 657.500000 294.410000 658.500000 295.590000 ;
      RECT 616.500000 294.410000 649.500000 295.590000 ;
      RECT 607.500000 294.410000 608.500000 295.590000 ;
      RECT 566.500000 294.410000 599.500000 295.590000 ;
      RECT 557.500000 294.410000 558.500000 295.590000 ;
      RECT 516.500000 294.410000 549.500000 295.590000 ;
      RECT 507.500000 294.410000 508.500000 295.590000 ;
      RECT 466.500000 294.410000 499.500000 295.590000 ;
      RECT 457.500000 294.410000 458.500000 295.590000 ;
      RECT 416.500000 294.410000 449.500000 295.590000 ;
      RECT 407.500000 294.410000 408.500000 295.590000 ;
      RECT 366.500000 294.410000 399.500000 295.590000 ;
      RECT 357.500000 294.410000 358.500000 295.590000 ;
      RECT 316.500000 294.410000 349.500000 295.590000 ;
      RECT 307.500000 294.410000 308.500000 295.590000 ;
      RECT 266.500000 294.410000 299.500000 295.590000 ;
      RECT 257.500000 294.410000 258.500000 295.590000 ;
      RECT 216.500000 294.410000 249.500000 295.590000 ;
      RECT 207.500000 294.410000 208.500000 295.590000 ;
      RECT 166.500000 294.410000 199.500000 295.590000 ;
      RECT 157.500000 294.410000 158.500000 295.590000 ;
      RECT 116.500000 294.410000 149.500000 295.590000 ;
      RECT 107.500000 294.410000 108.500000 295.590000 ;
      RECT 66.500000 294.410000 99.500000 295.590000 ;
      RECT 57.500000 294.410000 58.500000 295.590000 ;
      RECT 29.500000 294.410000 49.500000 295.590000 ;
      RECT 15.500000 294.410000 16.500000 295.590000 ;
      RECT 1157.500000 293.590000 1170.500000 294.410000 ;
      RECT 1107.500000 293.590000 1149.500000 294.410000 ;
      RECT 1057.500000 293.590000 1099.500000 294.410000 ;
      RECT 1007.500000 293.590000 1049.500000 294.410000 ;
      RECT 957.500000 293.590000 999.500000 294.410000 ;
      RECT 907.500000 293.590000 949.500000 294.410000 ;
      RECT 857.500000 293.590000 899.500000 294.410000 ;
      RECT 807.500000 293.590000 849.500000 294.410000 ;
      RECT 757.500000 293.590000 799.500000 294.410000 ;
      RECT 707.500000 293.590000 749.500000 294.410000 ;
      RECT 657.500000 293.590000 699.500000 294.410000 ;
      RECT 607.500000 293.590000 649.500000 294.410000 ;
      RECT 557.500000 293.590000 599.500000 294.410000 ;
      RECT 507.500000 293.590000 549.500000 294.410000 ;
      RECT 457.500000 293.590000 499.500000 294.410000 ;
      RECT 407.500000 293.590000 449.500000 294.410000 ;
      RECT 357.500000 293.590000 399.500000 294.410000 ;
      RECT 307.500000 293.590000 349.500000 294.410000 ;
      RECT 257.500000 293.590000 299.500000 294.410000 ;
      RECT 207.500000 293.590000 249.500000 294.410000 ;
      RECT 157.500000 293.590000 199.500000 294.410000 ;
      RECT 107.500000 293.590000 149.500000 294.410000 ;
      RECT 57.500000 293.590000 99.500000 294.410000 ;
      RECT 15.500000 293.590000 49.500000 294.410000 ;
      RECT 2.020000 293.515000 2.500000 295.590000 ;
      RECT 1183.500000 292.410000 1186.000000 295.590000 ;
      RECT 1169.500000 292.410000 1170.500000 293.590000 ;
      RECT 1116.500000 292.410000 1149.500000 293.590000 ;
      RECT 1107.500000 292.410000 1108.500000 293.590000 ;
      RECT 1066.500000 292.410000 1099.500000 293.590000 ;
      RECT 1057.500000 292.410000 1058.500000 293.590000 ;
      RECT 1016.500000 292.410000 1049.500000 293.590000 ;
      RECT 1007.500000 292.410000 1008.500000 293.590000 ;
      RECT 966.500000 292.410000 999.500000 293.590000 ;
      RECT 957.500000 292.410000 958.500000 293.590000 ;
      RECT 916.500000 292.410000 949.500000 293.590000 ;
      RECT 907.500000 292.410000 908.500000 293.590000 ;
      RECT 866.500000 292.410000 899.500000 293.590000 ;
      RECT 857.500000 292.410000 858.500000 293.590000 ;
      RECT 816.500000 292.410000 849.500000 293.590000 ;
      RECT 807.500000 292.410000 808.500000 293.590000 ;
      RECT 766.500000 292.410000 799.500000 293.590000 ;
      RECT 757.500000 292.410000 758.500000 293.590000 ;
      RECT 716.500000 292.410000 749.500000 293.590000 ;
      RECT 707.500000 292.410000 708.500000 293.590000 ;
      RECT 666.500000 292.410000 699.500000 293.590000 ;
      RECT 657.500000 292.410000 658.500000 293.590000 ;
      RECT 616.500000 292.410000 649.500000 293.590000 ;
      RECT 607.500000 292.410000 608.500000 293.590000 ;
      RECT 566.500000 292.410000 599.500000 293.590000 ;
      RECT 557.500000 292.410000 558.500000 293.590000 ;
      RECT 516.500000 292.410000 549.500000 293.590000 ;
      RECT 507.500000 292.410000 508.500000 293.590000 ;
      RECT 466.500000 292.410000 499.500000 293.590000 ;
      RECT 457.500000 292.410000 458.500000 293.590000 ;
      RECT 416.500000 292.410000 449.500000 293.590000 ;
      RECT 407.500000 292.410000 408.500000 293.590000 ;
      RECT 366.500000 292.410000 399.500000 293.590000 ;
      RECT 357.500000 292.410000 358.500000 293.590000 ;
      RECT 316.500000 292.410000 349.500000 293.590000 ;
      RECT 307.500000 292.410000 308.500000 293.590000 ;
      RECT 266.500000 292.410000 299.500000 293.590000 ;
      RECT 257.500000 292.410000 258.500000 293.590000 ;
      RECT 216.500000 292.410000 249.500000 293.590000 ;
      RECT 207.500000 292.410000 208.500000 293.590000 ;
      RECT 166.500000 292.410000 199.500000 293.590000 ;
      RECT 157.500000 292.410000 158.500000 293.590000 ;
      RECT 116.500000 292.410000 149.500000 293.590000 ;
      RECT 107.500000 292.410000 108.500000 293.590000 ;
      RECT 66.500000 292.410000 99.500000 293.590000 ;
      RECT 57.500000 292.410000 58.500000 293.590000 ;
      RECT 29.500000 292.410000 49.500000 293.590000 ;
      RECT 15.500000 292.410000 16.500000 293.590000 ;
      RECT 0.000000 292.410000 2.500000 293.515000 ;
      RECT 1169.500000 291.590000 1186.000000 292.410000 ;
      RECT 1116.500000 291.590000 1156.500000 292.410000 ;
      RECT 1066.500000 291.590000 1108.500000 292.410000 ;
      RECT 1016.500000 291.590000 1058.500000 292.410000 ;
      RECT 966.500000 291.590000 1008.500000 292.410000 ;
      RECT 916.500000 291.590000 958.500000 292.410000 ;
      RECT 866.500000 291.590000 908.500000 292.410000 ;
      RECT 816.500000 291.590000 858.500000 292.410000 ;
      RECT 766.500000 291.590000 808.500000 292.410000 ;
      RECT 716.500000 291.590000 758.500000 292.410000 ;
      RECT 666.500000 291.590000 708.500000 292.410000 ;
      RECT 616.500000 291.590000 658.500000 292.410000 ;
      RECT 566.500000 291.590000 608.500000 292.410000 ;
      RECT 516.500000 291.590000 558.500000 292.410000 ;
      RECT 466.500000 291.590000 508.500000 292.410000 ;
      RECT 416.500000 291.590000 458.500000 292.410000 ;
      RECT 366.500000 291.590000 408.500000 292.410000 ;
      RECT 316.500000 291.590000 358.500000 292.410000 ;
      RECT 266.500000 291.590000 308.500000 292.410000 ;
      RECT 216.500000 291.590000 258.500000 292.410000 ;
      RECT 166.500000 291.590000 208.500000 292.410000 ;
      RECT 116.500000 291.590000 158.500000 292.410000 ;
      RECT 66.500000 291.590000 108.500000 292.410000 ;
      RECT 29.500000 291.590000 58.500000 292.410000 ;
      RECT 0.000000 291.590000 16.500000 292.410000 ;
      RECT 0.000000 290.935000 2.500000 291.590000 ;
      RECT 1183.500000 290.930000 1186.000000 291.590000 ;
      RECT 1169.500000 290.410000 1170.500000 291.590000 ;
      RECT 1116.500000 290.410000 1149.500000 291.590000 ;
      RECT 1107.500000 290.410000 1108.500000 291.590000 ;
      RECT 1066.500000 290.410000 1099.500000 291.590000 ;
      RECT 1057.500000 290.410000 1058.500000 291.590000 ;
      RECT 1016.500000 290.410000 1049.500000 291.590000 ;
      RECT 1007.500000 290.410000 1008.500000 291.590000 ;
      RECT 966.500000 290.410000 999.500000 291.590000 ;
      RECT 957.500000 290.410000 958.500000 291.590000 ;
      RECT 916.500000 290.410000 949.500000 291.590000 ;
      RECT 907.500000 290.410000 908.500000 291.590000 ;
      RECT 866.500000 290.410000 899.500000 291.590000 ;
      RECT 857.500000 290.410000 858.500000 291.590000 ;
      RECT 816.500000 290.410000 849.500000 291.590000 ;
      RECT 807.500000 290.410000 808.500000 291.590000 ;
      RECT 766.500000 290.410000 799.500000 291.590000 ;
      RECT 757.500000 290.410000 758.500000 291.590000 ;
      RECT 716.500000 290.410000 749.500000 291.590000 ;
      RECT 707.500000 290.410000 708.500000 291.590000 ;
      RECT 666.500000 290.410000 699.500000 291.590000 ;
      RECT 657.500000 290.410000 658.500000 291.590000 ;
      RECT 616.500000 290.410000 649.500000 291.590000 ;
      RECT 607.500000 290.410000 608.500000 291.590000 ;
      RECT 566.500000 290.410000 599.500000 291.590000 ;
      RECT 557.500000 290.410000 558.500000 291.590000 ;
      RECT 516.500000 290.410000 549.500000 291.590000 ;
      RECT 507.500000 290.410000 508.500000 291.590000 ;
      RECT 466.500000 290.410000 499.500000 291.590000 ;
      RECT 457.500000 290.410000 458.500000 291.590000 ;
      RECT 416.500000 290.410000 449.500000 291.590000 ;
      RECT 407.500000 290.410000 408.500000 291.590000 ;
      RECT 366.500000 290.410000 399.500000 291.590000 ;
      RECT 357.500000 290.410000 358.500000 291.590000 ;
      RECT 316.500000 290.410000 349.500000 291.590000 ;
      RECT 307.500000 290.410000 308.500000 291.590000 ;
      RECT 266.500000 290.410000 299.500000 291.590000 ;
      RECT 257.500000 290.410000 258.500000 291.590000 ;
      RECT 216.500000 290.410000 249.500000 291.590000 ;
      RECT 207.500000 290.410000 208.500000 291.590000 ;
      RECT 166.500000 290.410000 199.500000 291.590000 ;
      RECT 157.500000 290.410000 158.500000 291.590000 ;
      RECT 116.500000 290.410000 149.500000 291.590000 ;
      RECT 107.500000 290.410000 108.500000 291.590000 ;
      RECT 66.500000 290.410000 99.500000 291.590000 ;
      RECT 57.500000 290.410000 58.500000 291.590000 ;
      RECT 29.500000 290.410000 49.500000 291.590000 ;
      RECT 15.500000 290.410000 16.500000 291.590000 ;
      RECT 1157.500000 289.590000 1170.500000 290.410000 ;
      RECT 1107.500000 289.590000 1149.500000 290.410000 ;
      RECT 1057.500000 289.590000 1099.500000 290.410000 ;
      RECT 1007.500000 289.590000 1049.500000 290.410000 ;
      RECT 957.500000 289.590000 999.500000 290.410000 ;
      RECT 907.500000 289.590000 949.500000 290.410000 ;
      RECT 857.500000 289.590000 899.500000 290.410000 ;
      RECT 807.500000 289.590000 849.500000 290.410000 ;
      RECT 757.500000 289.590000 799.500000 290.410000 ;
      RECT 707.500000 289.590000 749.500000 290.410000 ;
      RECT 657.500000 289.590000 699.500000 290.410000 ;
      RECT 607.500000 289.590000 649.500000 290.410000 ;
      RECT 557.500000 289.590000 599.500000 290.410000 ;
      RECT 507.500000 289.590000 549.500000 290.410000 ;
      RECT 457.500000 289.590000 499.500000 290.410000 ;
      RECT 407.500000 289.590000 449.500000 290.410000 ;
      RECT 357.500000 289.590000 399.500000 290.410000 ;
      RECT 307.500000 289.590000 349.500000 290.410000 ;
      RECT 257.500000 289.590000 299.500000 290.410000 ;
      RECT 207.500000 289.590000 249.500000 290.410000 ;
      RECT 157.500000 289.590000 199.500000 290.410000 ;
      RECT 107.500000 289.590000 149.500000 290.410000 ;
      RECT 57.500000 289.590000 99.500000 290.410000 ;
      RECT 15.500000 289.590000 49.500000 290.410000 ;
      RECT 1183.500000 288.410000 1183.980000 290.930000 ;
      RECT 1169.500000 288.410000 1170.500000 289.590000 ;
      RECT 1116.500000 288.410000 1149.500000 289.590000 ;
      RECT 1107.500000 288.410000 1108.500000 289.590000 ;
      RECT 1066.500000 288.410000 1099.500000 289.590000 ;
      RECT 1057.500000 288.410000 1058.500000 289.590000 ;
      RECT 1016.500000 288.410000 1049.500000 289.590000 ;
      RECT 1007.500000 288.410000 1008.500000 289.590000 ;
      RECT 966.500000 288.410000 999.500000 289.590000 ;
      RECT 957.500000 288.410000 958.500000 289.590000 ;
      RECT 916.500000 288.410000 949.500000 289.590000 ;
      RECT 907.500000 288.410000 908.500000 289.590000 ;
      RECT 866.500000 288.410000 899.500000 289.590000 ;
      RECT 857.500000 288.410000 858.500000 289.590000 ;
      RECT 816.500000 288.410000 849.500000 289.590000 ;
      RECT 807.500000 288.410000 808.500000 289.590000 ;
      RECT 766.500000 288.410000 799.500000 289.590000 ;
      RECT 757.500000 288.410000 758.500000 289.590000 ;
      RECT 716.500000 288.410000 749.500000 289.590000 ;
      RECT 707.500000 288.410000 708.500000 289.590000 ;
      RECT 666.500000 288.410000 699.500000 289.590000 ;
      RECT 657.500000 288.410000 658.500000 289.590000 ;
      RECT 616.500000 288.410000 649.500000 289.590000 ;
      RECT 607.500000 288.410000 608.500000 289.590000 ;
      RECT 566.500000 288.410000 599.500000 289.590000 ;
      RECT 557.500000 288.410000 558.500000 289.590000 ;
      RECT 516.500000 288.410000 549.500000 289.590000 ;
      RECT 507.500000 288.410000 508.500000 289.590000 ;
      RECT 466.500000 288.410000 499.500000 289.590000 ;
      RECT 457.500000 288.410000 458.500000 289.590000 ;
      RECT 416.500000 288.410000 449.500000 289.590000 ;
      RECT 407.500000 288.410000 408.500000 289.590000 ;
      RECT 366.500000 288.410000 399.500000 289.590000 ;
      RECT 357.500000 288.410000 358.500000 289.590000 ;
      RECT 316.500000 288.410000 349.500000 289.590000 ;
      RECT 307.500000 288.410000 308.500000 289.590000 ;
      RECT 266.500000 288.410000 299.500000 289.590000 ;
      RECT 257.500000 288.410000 258.500000 289.590000 ;
      RECT 216.500000 288.410000 249.500000 289.590000 ;
      RECT 207.500000 288.410000 208.500000 289.590000 ;
      RECT 166.500000 288.410000 199.500000 289.590000 ;
      RECT 157.500000 288.410000 158.500000 289.590000 ;
      RECT 116.500000 288.410000 149.500000 289.590000 ;
      RECT 107.500000 288.410000 108.500000 289.590000 ;
      RECT 66.500000 288.410000 99.500000 289.590000 ;
      RECT 57.500000 288.410000 58.500000 289.590000 ;
      RECT 29.500000 288.410000 49.500000 289.590000 ;
      RECT 15.500000 288.410000 16.500000 289.590000 ;
      RECT 2.020000 288.410000 2.500000 290.935000 ;
      RECT 2.020000 287.835000 16.500000 288.410000 ;
      RECT 1169.500000 287.830000 1183.980000 288.410000 ;
      RECT 1169.500000 287.590000 1186.000000 287.830000 ;
      RECT 1116.500000 287.590000 1156.500000 288.410000 ;
      RECT 1066.500000 287.590000 1108.500000 288.410000 ;
      RECT 1016.500000 287.590000 1058.500000 288.410000 ;
      RECT 966.500000 287.590000 1008.500000 288.410000 ;
      RECT 916.500000 287.590000 958.500000 288.410000 ;
      RECT 866.500000 287.590000 908.500000 288.410000 ;
      RECT 816.500000 287.590000 858.500000 288.410000 ;
      RECT 766.500000 287.590000 808.500000 288.410000 ;
      RECT 716.500000 287.590000 758.500000 288.410000 ;
      RECT 666.500000 287.590000 708.500000 288.410000 ;
      RECT 616.500000 287.590000 658.500000 288.410000 ;
      RECT 566.500000 287.590000 608.500000 288.410000 ;
      RECT 516.500000 287.590000 558.500000 288.410000 ;
      RECT 466.500000 287.590000 508.500000 288.410000 ;
      RECT 416.500000 287.590000 458.500000 288.410000 ;
      RECT 366.500000 287.590000 408.500000 288.410000 ;
      RECT 316.500000 287.590000 358.500000 288.410000 ;
      RECT 266.500000 287.590000 308.500000 288.410000 ;
      RECT 216.500000 287.590000 258.500000 288.410000 ;
      RECT 166.500000 287.590000 208.500000 288.410000 ;
      RECT 116.500000 287.590000 158.500000 288.410000 ;
      RECT 66.500000 287.590000 108.500000 288.410000 ;
      RECT 29.500000 287.590000 58.500000 288.410000 ;
      RECT 0.000000 287.590000 16.500000 287.835000 ;
      RECT 1169.500000 286.410000 1170.500000 287.590000 ;
      RECT 1116.500000 286.410000 1149.500000 287.590000 ;
      RECT 1107.500000 286.410000 1108.500000 287.590000 ;
      RECT 1066.500000 286.410000 1099.500000 287.590000 ;
      RECT 1057.500000 286.410000 1058.500000 287.590000 ;
      RECT 1016.500000 286.410000 1049.500000 287.590000 ;
      RECT 1007.500000 286.410000 1008.500000 287.590000 ;
      RECT 966.500000 286.410000 999.500000 287.590000 ;
      RECT 957.500000 286.410000 958.500000 287.590000 ;
      RECT 916.500000 286.410000 949.500000 287.590000 ;
      RECT 907.500000 286.410000 908.500000 287.590000 ;
      RECT 866.500000 286.410000 899.500000 287.590000 ;
      RECT 857.500000 286.410000 858.500000 287.590000 ;
      RECT 816.500000 286.410000 849.500000 287.590000 ;
      RECT 807.500000 286.410000 808.500000 287.590000 ;
      RECT 766.500000 286.410000 799.500000 287.590000 ;
      RECT 757.500000 286.410000 758.500000 287.590000 ;
      RECT 716.500000 286.410000 749.500000 287.590000 ;
      RECT 707.500000 286.410000 708.500000 287.590000 ;
      RECT 666.500000 286.410000 699.500000 287.590000 ;
      RECT 657.500000 286.410000 658.500000 287.590000 ;
      RECT 616.500000 286.410000 649.500000 287.590000 ;
      RECT 607.500000 286.410000 608.500000 287.590000 ;
      RECT 566.500000 286.410000 599.500000 287.590000 ;
      RECT 557.500000 286.410000 558.500000 287.590000 ;
      RECT 516.500000 286.410000 549.500000 287.590000 ;
      RECT 507.500000 286.410000 508.500000 287.590000 ;
      RECT 466.500000 286.410000 499.500000 287.590000 ;
      RECT 457.500000 286.410000 458.500000 287.590000 ;
      RECT 416.500000 286.410000 449.500000 287.590000 ;
      RECT 407.500000 286.410000 408.500000 287.590000 ;
      RECT 366.500000 286.410000 399.500000 287.590000 ;
      RECT 357.500000 286.410000 358.500000 287.590000 ;
      RECT 316.500000 286.410000 349.500000 287.590000 ;
      RECT 307.500000 286.410000 308.500000 287.590000 ;
      RECT 266.500000 286.410000 299.500000 287.590000 ;
      RECT 257.500000 286.410000 258.500000 287.590000 ;
      RECT 216.500000 286.410000 249.500000 287.590000 ;
      RECT 207.500000 286.410000 208.500000 287.590000 ;
      RECT 166.500000 286.410000 199.500000 287.590000 ;
      RECT 157.500000 286.410000 158.500000 287.590000 ;
      RECT 116.500000 286.410000 149.500000 287.590000 ;
      RECT 107.500000 286.410000 108.500000 287.590000 ;
      RECT 66.500000 286.410000 99.500000 287.590000 ;
      RECT 57.500000 286.410000 58.500000 287.590000 ;
      RECT 29.500000 286.410000 49.500000 287.590000 ;
      RECT 15.500000 286.410000 16.500000 287.590000 ;
      RECT 1157.500000 285.590000 1170.500000 286.410000 ;
      RECT 1107.500000 285.590000 1149.500000 286.410000 ;
      RECT 1057.500000 285.590000 1099.500000 286.410000 ;
      RECT 1007.500000 285.590000 1049.500000 286.410000 ;
      RECT 957.500000 285.590000 999.500000 286.410000 ;
      RECT 907.500000 285.590000 949.500000 286.410000 ;
      RECT 857.500000 285.590000 899.500000 286.410000 ;
      RECT 807.500000 285.590000 849.500000 286.410000 ;
      RECT 757.500000 285.590000 799.500000 286.410000 ;
      RECT 707.500000 285.590000 749.500000 286.410000 ;
      RECT 657.500000 285.590000 699.500000 286.410000 ;
      RECT 607.500000 285.590000 649.500000 286.410000 ;
      RECT 557.500000 285.590000 599.500000 286.410000 ;
      RECT 507.500000 285.590000 549.500000 286.410000 ;
      RECT 457.500000 285.590000 499.500000 286.410000 ;
      RECT 407.500000 285.590000 449.500000 286.410000 ;
      RECT 357.500000 285.590000 399.500000 286.410000 ;
      RECT 307.500000 285.590000 349.500000 286.410000 ;
      RECT 257.500000 285.590000 299.500000 286.410000 ;
      RECT 207.500000 285.590000 249.500000 286.410000 ;
      RECT 157.500000 285.590000 199.500000 286.410000 ;
      RECT 107.500000 285.590000 149.500000 286.410000 ;
      RECT 57.500000 285.590000 99.500000 286.410000 ;
      RECT 15.500000 285.590000 49.500000 286.410000 ;
      RECT 1183.500000 284.410000 1186.000000 287.590000 ;
      RECT 1169.500000 284.410000 1170.500000 285.590000 ;
      RECT 1116.500000 284.410000 1149.500000 285.590000 ;
      RECT 1107.500000 284.410000 1108.500000 285.590000 ;
      RECT 1066.500000 284.410000 1099.500000 285.590000 ;
      RECT 1057.500000 284.410000 1058.500000 285.590000 ;
      RECT 1016.500000 284.410000 1049.500000 285.590000 ;
      RECT 1007.500000 284.410000 1008.500000 285.590000 ;
      RECT 966.500000 284.410000 999.500000 285.590000 ;
      RECT 957.500000 284.410000 958.500000 285.590000 ;
      RECT 916.500000 284.410000 949.500000 285.590000 ;
      RECT 907.500000 284.410000 908.500000 285.590000 ;
      RECT 866.500000 284.410000 899.500000 285.590000 ;
      RECT 857.500000 284.410000 858.500000 285.590000 ;
      RECT 816.500000 284.410000 849.500000 285.590000 ;
      RECT 807.500000 284.410000 808.500000 285.590000 ;
      RECT 766.500000 284.410000 799.500000 285.590000 ;
      RECT 757.500000 284.410000 758.500000 285.590000 ;
      RECT 716.500000 284.410000 749.500000 285.590000 ;
      RECT 707.500000 284.410000 708.500000 285.590000 ;
      RECT 666.500000 284.410000 699.500000 285.590000 ;
      RECT 657.500000 284.410000 658.500000 285.590000 ;
      RECT 616.500000 284.410000 649.500000 285.590000 ;
      RECT 607.500000 284.410000 608.500000 285.590000 ;
      RECT 566.500000 284.410000 599.500000 285.590000 ;
      RECT 557.500000 284.410000 558.500000 285.590000 ;
      RECT 516.500000 284.410000 549.500000 285.590000 ;
      RECT 507.500000 284.410000 508.500000 285.590000 ;
      RECT 466.500000 284.410000 499.500000 285.590000 ;
      RECT 457.500000 284.410000 458.500000 285.590000 ;
      RECT 416.500000 284.410000 449.500000 285.590000 ;
      RECT 407.500000 284.410000 408.500000 285.590000 ;
      RECT 366.500000 284.410000 399.500000 285.590000 ;
      RECT 357.500000 284.410000 358.500000 285.590000 ;
      RECT 316.500000 284.410000 349.500000 285.590000 ;
      RECT 307.500000 284.410000 308.500000 285.590000 ;
      RECT 266.500000 284.410000 299.500000 285.590000 ;
      RECT 257.500000 284.410000 258.500000 285.590000 ;
      RECT 216.500000 284.410000 249.500000 285.590000 ;
      RECT 207.500000 284.410000 208.500000 285.590000 ;
      RECT 166.500000 284.410000 199.500000 285.590000 ;
      RECT 157.500000 284.410000 158.500000 285.590000 ;
      RECT 116.500000 284.410000 149.500000 285.590000 ;
      RECT 107.500000 284.410000 108.500000 285.590000 ;
      RECT 66.500000 284.410000 99.500000 285.590000 ;
      RECT 57.500000 284.410000 58.500000 285.590000 ;
      RECT 29.500000 284.410000 49.500000 285.590000 ;
      RECT 15.500000 284.410000 16.500000 285.590000 ;
      RECT 0.000000 284.410000 2.500000 287.590000 ;
      RECT 1169.500000 283.590000 1186.000000 284.410000 ;
      RECT 1116.500000 283.590000 1156.500000 284.410000 ;
      RECT 1066.500000 283.590000 1108.500000 284.410000 ;
      RECT 1016.500000 283.590000 1058.500000 284.410000 ;
      RECT 966.500000 283.590000 1008.500000 284.410000 ;
      RECT 916.500000 283.590000 958.500000 284.410000 ;
      RECT 866.500000 283.590000 908.500000 284.410000 ;
      RECT 816.500000 283.590000 858.500000 284.410000 ;
      RECT 766.500000 283.590000 808.500000 284.410000 ;
      RECT 716.500000 283.590000 758.500000 284.410000 ;
      RECT 666.500000 283.590000 708.500000 284.410000 ;
      RECT 616.500000 283.590000 658.500000 284.410000 ;
      RECT 566.500000 283.590000 608.500000 284.410000 ;
      RECT 516.500000 283.590000 558.500000 284.410000 ;
      RECT 466.500000 283.590000 508.500000 284.410000 ;
      RECT 416.500000 283.590000 458.500000 284.410000 ;
      RECT 366.500000 283.590000 408.500000 284.410000 ;
      RECT 316.500000 283.590000 358.500000 284.410000 ;
      RECT 266.500000 283.590000 308.500000 284.410000 ;
      RECT 216.500000 283.590000 258.500000 284.410000 ;
      RECT 166.500000 283.590000 208.500000 284.410000 ;
      RECT 116.500000 283.590000 158.500000 284.410000 ;
      RECT 66.500000 283.590000 108.500000 284.410000 ;
      RECT 29.500000 283.590000 58.500000 284.410000 ;
      RECT 0.000000 283.590000 16.500000 284.410000 ;
      RECT 1169.500000 282.410000 1170.500000 283.590000 ;
      RECT 1116.500000 282.410000 1149.500000 283.590000 ;
      RECT 1107.500000 282.410000 1108.500000 283.590000 ;
      RECT 1066.500000 282.410000 1099.500000 283.590000 ;
      RECT 1057.500000 282.410000 1058.500000 283.590000 ;
      RECT 1016.500000 282.410000 1049.500000 283.590000 ;
      RECT 1007.500000 282.410000 1008.500000 283.590000 ;
      RECT 966.500000 282.410000 999.500000 283.590000 ;
      RECT 957.500000 282.410000 958.500000 283.590000 ;
      RECT 916.500000 282.410000 949.500000 283.590000 ;
      RECT 907.500000 282.410000 908.500000 283.590000 ;
      RECT 866.500000 282.410000 899.500000 283.590000 ;
      RECT 857.500000 282.410000 858.500000 283.590000 ;
      RECT 816.500000 282.410000 849.500000 283.590000 ;
      RECT 807.500000 282.410000 808.500000 283.590000 ;
      RECT 766.500000 282.410000 799.500000 283.590000 ;
      RECT 757.500000 282.410000 758.500000 283.590000 ;
      RECT 716.500000 282.410000 749.500000 283.590000 ;
      RECT 707.500000 282.410000 708.500000 283.590000 ;
      RECT 666.500000 282.410000 699.500000 283.590000 ;
      RECT 657.500000 282.410000 658.500000 283.590000 ;
      RECT 616.500000 282.410000 649.500000 283.590000 ;
      RECT 607.500000 282.410000 608.500000 283.590000 ;
      RECT 566.500000 282.410000 599.500000 283.590000 ;
      RECT 557.500000 282.410000 558.500000 283.590000 ;
      RECT 516.500000 282.410000 549.500000 283.590000 ;
      RECT 507.500000 282.410000 508.500000 283.590000 ;
      RECT 466.500000 282.410000 499.500000 283.590000 ;
      RECT 457.500000 282.410000 458.500000 283.590000 ;
      RECT 416.500000 282.410000 449.500000 283.590000 ;
      RECT 407.500000 282.410000 408.500000 283.590000 ;
      RECT 366.500000 282.410000 399.500000 283.590000 ;
      RECT 357.500000 282.410000 358.500000 283.590000 ;
      RECT 316.500000 282.410000 349.500000 283.590000 ;
      RECT 307.500000 282.410000 308.500000 283.590000 ;
      RECT 266.500000 282.410000 299.500000 283.590000 ;
      RECT 257.500000 282.410000 258.500000 283.590000 ;
      RECT 216.500000 282.410000 249.500000 283.590000 ;
      RECT 207.500000 282.410000 208.500000 283.590000 ;
      RECT 166.500000 282.410000 199.500000 283.590000 ;
      RECT 157.500000 282.410000 158.500000 283.590000 ;
      RECT 116.500000 282.410000 149.500000 283.590000 ;
      RECT 107.500000 282.410000 108.500000 283.590000 ;
      RECT 66.500000 282.410000 99.500000 283.590000 ;
      RECT 57.500000 282.410000 58.500000 283.590000 ;
      RECT 29.500000 282.410000 49.500000 283.590000 ;
      RECT 15.500000 282.410000 16.500000 283.590000 ;
      RECT 1157.500000 281.590000 1170.500000 282.410000 ;
      RECT 1107.500000 281.590000 1149.500000 282.410000 ;
      RECT 1057.500000 281.590000 1099.500000 282.410000 ;
      RECT 1007.500000 281.590000 1049.500000 282.410000 ;
      RECT 957.500000 281.590000 999.500000 282.410000 ;
      RECT 907.500000 281.590000 949.500000 282.410000 ;
      RECT 857.500000 281.590000 899.500000 282.410000 ;
      RECT 807.500000 281.590000 849.500000 282.410000 ;
      RECT 757.500000 281.590000 799.500000 282.410000 ;
      RECT 707.500000 281.590000 749.500000 282.410000 ;
      RECT 657.500000 281.590000 699.500000 282.410000 ;
      RECT 607.500000 281.590000 649.500000 282.410000 ;
      RECT 557.500000 281.590000 599.500000 282.410000 ;
      RECT 507.500000 281.590000 549.500000 282.410000 ;
      RECT 457.500000 281.590000 499.500000 282.410000 ;
      RECT 407.500000 281.590000 449.500000 282.410000 ;
      RECT 357.500000 281.590000 399.500000 282.410000 ;
      RECT 307.500000 281.590000 349.500000 282.410000 ;
      RECT 257.500000 281.590000 299.500000 282.410000 ;
      RECT 207.500000 281.590000 249.500000 282.410000 ;
      RECT 157.500000 281.590000 199.500000 282.410000 ;
      RECT 107.500000 281.590000 149.500000 282.410000 ;
      RECT 57.500000 281.590000 99.500000 282.410000 ;
      RECT 15.500000 281.590000 49.500000 282.410000 ;
      RECT 1183.500000 280.410000 1186.000000 283.590000 ;
      RECT 1169.500000 280.410000 1170.500000 281.590000 ;
      RECT 1116.500000 280.410000 1149.500000 281.590000 ;
      RECT 1107.500000 280.410000 1108.500000 281.590000 ;
      RECT 1066.500000 280.410000 1099.500000 281.590000 ;
      RECT 1057.500000 280.410000 1058.500000 281.590000 ;
      RECT 1016.500000 280.410000 1049.500000 281.590000 ;
      RECT 1007.500000 280.410000 1008.500000 281.590000 ;
      RECT 966.500000 280.410000 999.500000 281.590000 ;
      RECT 957.500000 280.410000 958.500000 281.590000 ;
      RECT 916.500000 280.410000 949.500000 281.590000 ;
      RECT 907.500000 280.410000 908.500000 281.590000 ;
      RECT 866.500000 280.410000 899.500000 281.590000 ;
      RECT 857.500000 280.410000 858.500000 281.590000 ;
      RECT 816.500000 280.410000 849.500000 281.590000 ;
      RECT 807.500000 280.410000 808.500000 281.590000 ;
      RECT 766.500000 280.410000 799.500000 281.590000 ;
      RECT 757.500000 280.410000 758.500000 281.590000 ;
      RECT 716.500000 280.410000 749.500000 281.590000 ;
      RECT 707.500000 280.410000 708.500000 281.590000 ;
      RECT 666.500000 280.410000 699.500000 281.590000 ;
      RECT 657.500000 280.410000 658.500000 281.590000 ;
      RECT 616.500000 280.410000 649.500000 281.590000 ;
      RECT 607.500000 280.410000 608.500000 281.590000 ;
      RECT 566.500000 280.410000 599.500000 281.590000 ;
      RECT 557.500000 280.410000 558.500000 281.590000 ;
      RECT 516.500000 280.410000 549.500000 281.590000 ;
      RECT 507.500000 280.410000 508.500000 281.590000 ;
      RECT 466.500000 280.410000 499.500000 281.590000 ;
      RECT 457.500000 280.410000 458.500000 281.590000 ;
      RECT 416.500000 280.410000 449.500000 281.590000 ;
      RECT 407.500000 280.410000 408.500000 281.590000 ;
      RECT 366.500000 280.410000 399.500000 281.590000 ;
      RECT 357.500000 280.410000 358.500000 281.590000 ;
      RECT 316.500000 280.410000 349.500000 281.590000 ;
      RECT 307.500000 280.410000 308.500000 281.590000 ;
      RECT 266.500000 280.410000 299.500000 281.590000 ;
      RECT 257.500000 280.410000 258.500000 281.590000 ;
      RECT 216.500000 280.410000 249.500000 281.590000 ;
      RECT 207.500000 280.410000 208.500000 281.590000 ;
      RECT 166.500000 280.410000 199.500000 281.590000 ;
      RECT 157.500000 280.410000 158.500000 281.590000 ;
      RECT 116.500000 280.410000 149.500000 281.590000 ;
      RECT 107.500000 280.410000 108.500000 281.590000 ;
      RECT 66.500000 280.410000 99.500000 281.590000 ;
      RECT 57.500000 280.410000 58.500000 281.590000 ;
      RECT 29.500000 280.410000 49.500000 281.590000 ;
      RECT 15.500000 280.410000 16.500000 281.590000 ;
      RECT 0.000000 280.410000 2.500000 283.590000 ;
      RECT 1169.500000 279.590000 1186.000000 280.410000 ;
      RECT 1116.500000 279.590000 1156.500000 280.410000 ;
      RECT 1066.500000 279.590000 1108.500000 280.410000 ;
      RECT 1016.500000 279.590000 1058.500000 280.410000 ;
      RECT 966.500000 279.590000 1008.500000 280.410000 ;
      RECT 916.500000 279.590000 958.500000 280.410000 ;
      RECT 866.500000 279.590000 908.500000 280.410000 ;
      RECT 816.500000 279.590000 858.500000 280.410000 ;
      RECT 766.500000 279.590000 808.500000 280.410000 ;
      RECT 716.500000 279.590000 758.500000 280.410000 ;
      RECT 666.500000 279.590000 708.500000 280.410000 ;
      RECT 616.500000 279.590000 658.500000 280.410000 ;
      RECT 566.500000 279.590000 608.500000 280.410000 ;
      RECT 516.500000 279.590000 558.500000 280.410000 ;
      RECT 466.500000 279.590000 508.500000 280.410000 ;
      RECT 416.500000 279.590000 458.500000 280.410000 ;
      RECT 366.500000 279.590000 408.500000 280.410000 ;
      RECT 316.500000 279.590000 358.500000 280.410000 ;
      RECT 266.500000 279.590000 308.500000 280.410000 ;
      RECT 216.500000 279.590000 258.500000 280.410000 ;
      RECT 166.500000 279.590000 208.500000 280.410000 ;
      RECT 116.500000 279.590000 158.500000 280.410000 ;
      RECT 66.500000 279.590000 108.500000 280.410000 ;
      RECT 29.500000 279.590000 58.500000 280.410000 ;
      RECT 0.000000 279.590000 16.500000 280.410000 ;
      RECT 1169.500000 278.410000 1170.500000 279.590000 ;
      RECT 1116.500000 278.410000 1149.500000 279.590000 ;
      RECT 1107.500000 278.410000 1108.500000 279.590000 ;
      RECT 1066.500000 278.410000 1099.500000 279.590000 ;
      RECT 1057.500000 278.410000 1058.500000 279.590000 ;
      RECT 1016.500000 278.410000 1049.500000 279.590000 ;
      RECT 1007.500000 278.410000 1008.500000 279.590000 ;
      RECT 966.500000 278.410000 999.500000 279.590000 ;
      RECT 957.500000 278.410000 958.500000 279.590000 ;
      RECT 916.500000 278.410000 949.500000 279.590000 ;
      RECT 907.500000 278.410000 908.500000 279.590000 ;
      RECT 866.500000 278.410000 899.500000 279.590000 ;
      RECT 857.500000 278.410000 858.500000 279.590000 ;
      RECT 816.500000 278.410000 849.500000 279.590000 ;
      RECT 807.500000 278.410000 808.500000 279.590000 ;
      RECT 766.500000 278.410000 799.500000 279.590000 ;
      RECT 757.500000 278.410000 758.500000 279.590000 ;
      RECT 716.500000 278.410000 749.500000 279.590000 ;
      RECT 707.500000 278.410000 708.500000 279.590000 ;
      RECT 666.500000 278.410000 699.500000 279.590000 ;
      RECT 657.500000 278.410000 658.500000 279.590000 ;
      RECT 616.500000 278.410000 649.500000 279.590000 ;
      RECT 607.500000 278.410000 608.500000 279.590000 ;
      RECT 566.500000 278.410000 599.500000 279.590000 ;
      RECT 557.500000 278.410000 558.500000 279.590000 ;
      RECT 516.500000 278.410000 549.500000 279.590000 ;
      RECT 507.500000 278.410000 508.500000 279.590000 ;
      RECT 466.500000 278.410000 499.500000 279.590000 ;
      RECT 457.500000 278.410000 458.500000 279.590000 ;
      RECT 416.500000 278.410000 449.500000 279.590000 ;
      RECT 407.500000 278.410000 408.500000 279.590000 ;
      RECT 366.500000 278.410000 399.500000 279.590000 ;
      RECT 357.500000 278.410000 358.500000 279.590000 ;
      RECT 316.500000 278.410000 349.500000 279.590000 ;
      RECT 307.500000 278.410000 308.500000 279.590000 ;
      RECT 266.500000 278.410000 299.500000 279.590000 ;
      RECT 257.500000 278.410000 258.500000 279.590000 ;
      RECT 216.500000 278.410000 249.500000 279.590000 ;
      RECT 207.500000 278.410000 208.500000 279.590000 ;
      RECT 166.500000 278.410000 199.500000 279.590000 ;
      RECT 157.500000 278.410000 158.500000 279.590000 ;
      RECT 116.500000 278.410000 149.500000 279.590000 ;
      RECT 107.500000 278.410000 108.500000 279.590000 ;
      RECT 66.500000 278.410000 99.500000 279.590000 ;
      RECT 57.500000 278.410000 58.500000 279.590000 ;
      RECT 29.500000 278.410000 49.500000 279.590000 ;
      RECT 15.500000 278.410000 16.500000 279.590000 ;
      RECT 1157.500000 277.590000 1170.500000 278.410000 ;
      RECT 1107.500000 277.590000 1149.500000 278.410000 ;
      RECT 1057.500000 277.590000 1099.500000 278.410000 ;
      RECT 1007.500000 277.590000 1049.500000 278.410000 ;
      RECT 957.500000 277.590000 999.500000 278.410000 ;
      RECT 907.500000 277.590000 949.500000 278.410000 ;
      RECT 857.500000 277.590000 899.500000 278.410000 ;
      RECT 807.500000 277.590000 849.500000 278.410000 ;
      RECT 757.500000 277.590000 799.500000 278.410000 ;
      RECT 707.500000 277.590000 749.500000 278.410000 ;
      RECT 657.500000 277.590000 699.500000 278.410000 ;
      RECT 607.500000 277.590000 649.500000 278.410000 ;
      RECT 557.500000 277.590000 599.500000 278.410000 ;
      RECT 507.500000 277.590000 549.500000 278.410000 ;
      RECT 457.500000 277.590000 499.500000 278.410000 ;
      RECT 407.500000 277.590000 449.500000 278.410000 ;
      RECT 357.500000 277.590000 399.500000 278.410000 ;
      RECT 307.500000 277.590000 349.500000 278.410000 ;
      RECT 257.500000 277.590000 299.500000 278.410000 ;
      RECT 207.500000 277.590000 249.500000 278.410000 ;
      RECT 157.500000 277.590000 199.500000 278.410000 ;
      RECT 107.500000 277.590000 149.500000 278.410000 ;
      RECT 57.500000 277.590000 99.500000 278.410000 ;
      RECT 15.500000 277.590000 49.500000 278.410000 ;
      RECT 1183.500000 276.410000 1186.000000 279.590000 ;
      RECT 1169.500000 276.410000 1170.500000 277.590000 ;
      RECT 1116.500000 276.410000 1149.500000 277.590000 ;
      RECT 1107.500000 276.410000 1108.500000 277.590000 ;
      RECT 1066.500000 276.410000 1099.500000 277.590000 ;
      RECT 1057.500000 276.410000 1058.500000 277.590000 ;
      RECT 1016.500000 276.410000 1049.500000 277.590000 ;
      RECT 1007.500000 276.410000 1008.500000 277.590000 ;
      RECT 966.500000 276.410000 999.500000 277.590000 ;
      RECT 957.500000 276.410000 958.500000 277.590000 ;
      RECT 916.500000 276.410000 949.500000 277.590000 ;
      RECT 907.500000 276.410000 908.500000 277.590000 ;
      RECT 866.500000 276.410000 899.500000 277.590000 ;
      RECT 857.500000 276.410000 858.500000 277.590000 ;
      RECT 816.500000 276.410000 849.500000 277.590000 ;
      RECT 807.500000 276.410000 808.500000 277.590000 ;
      RECT 766.500000 276.410000 799.500000 277.590000 ;
      RECT 757.500000 276.410000 758.500000 277.590000 ;
      RECT 716.500000 276.410000 749.500000 277.590000 ;
      RECT 707.500000 276.410000 708.500000 277.590000 ;
      RECT 666.500000 276.410000 699.500000 277.590000 ;
      RECT 657.500000 276.410000 658.500000 277.590000 ;
      RECT 616.500000 276.410000 649.500000 277.590000 ;
      RECT 607.500000 276.410000 608.500000 277.590000 ;
      RECT 566.500000 276.410000 599.500000 277.590000 ;
      RECT 557.500000 276.410000 558.500000 277.590000 ;
      RECT 516.500000 276.410000 549.500000 277.590000 ;
      RECT 507.500000 276.410000 508.500000 277.590000 ;
      RECT 466.500000 276.410000 499.500000 277.590000 ;
      RECT 457.500000 276.410000 458.500000 277.590000 ;
      RECT 416.500000 276.410000 449.500000 277.590000 ;
      RECT 407.500000 276.410000 408.500000 277.590000 ;
      RECT 366.500000 276.410000 399.500000 277.590000 ;
      RECT 357.500000 276.410000 358.500000 277.590000 ;
      RECT 316.500000 276.410000 349.500000 277.590000 ;
      RECT 307.500000 276.410000 308.500000 277.590000 ;
      RECT 266.500000 276.410000 299.500000 277.590000 ;
      RECT 257.500000 276.410000 258.500000 277.590000 ;
      RECT 216.500000 276.410000 249.500000 277.590000 ;
      RECT 207.500000 276.410000 208.500000 277.590000 ;
      RECT 166.500000 276.410000 199.500000 277.590000 ;
      RECT 157.500000 276.410000 158.500000 277.590000 ;
      RECT 116.500000 276.410000 149.500000 277.590000 ;
      RECT 107.500000 276.410000 108.500000 277.590000 ;
      RECT 66.500000 276.410000 99.500000 277.590000 ;
      RECT 57.500000 276.410000 58.500000 277.590000 ;
      RECT 29.500000 276.410000 49.500000 277.590000 ;
      RECT 15.500000 276.410000 16.500000 277.590000 ;
      RECT 0.000000 276.410000 2.500000 279.590000 ;
      RECT 1169.500000 275.590000 1186.000000 276.410000 ;
      RECT 1116.500000 275.590000 1156.500000 276.410000 ;
      RECT 1066.500000 275.590000 1108.500000 276.410000 ;
      RECT 1016.500000 275.590000 1058.500000 276.410000 ;
      RECT 966.500000 275.590000 1008.500000 276.410000 ;
      RECT 916.500000 275.590000 958.500000 276.410000 ;
      RECT 866.500000 275.590000 908.500000 276.410000 ;
      RECT 816.500000 275.590000 858.500000 276.410000 ;
      RECT 766.500000 275.590000 808.500000 276.410000 ;
      RECT 716.500000 275.590000 758.500000 276.410000 ;
      RECT 666.500000 275.590000 708.500000 276.410000 ;
      RECT 616.500000 275.590000 658.500000 276.410000 ;
      RECT 566.500000 275.590000 608.500000 276.410000 ;
      RECT 516.500000 275.590000 558.500000 276.410000 ;
      RECT 466.500000 275.590000 508.500000 276.410000 ;
      RECT 416.500000 275.590000 458.500000 276.410000 ;
      RECT 366.500000 275.590000 408.500000 276.410000 ;
      RECT 316.500000 275.590000 358.500000 276.410000 ;
      RECT 266.500000 275.590000 308.500000 276.410000 ;
      RECT 216.500000 275.590000 258.500000 276.410000 ;
      RECT 166.500000 275.590000 208.500000 276.410000 ;
      RECT 116.500000 275.590000 158.500000 276.410000 ;
      RECT 66.500000 275.590000 108.500000 276.410000 ;
      RECT 29.500000 275.590000 58.500000 276.410000 ;
      RECT 0.000000 275.590000 16.500000 276.410000 ;
      RECT 1169.500000 274.410000 1170.500000 275.590000 ;
      RECT 1116.500000 274.410000 1149.500000 275.590000 ;
      RECT 1107.500000 274.410000 1108.500000 275.590000 ;
      RECT 1066.500000 274.410000 1099.500000 275.590000 ;
      RECT 1057.500000 274.410000 1058.500000 275.590000 ;
      RECT 1016.500000 274.410000 1049.500000 275.590000 ;
      RECT 1007.500000 274.410000 1008.500000 275.590000 ;
      RECT 966.500000 274.410000 999.500000 275.590000 ;
      RECT 957.500000 274.410000 958.500000 275.590000 ;
      RECT 916.500000 274.410000 949.500000 275.590000 ;
      RECT 907.500000 274.410000 908.500000 275.590000 ;
      RECT 866.500000 274.410000 899.500000 275.590000 ;
      RECT 857.500000 274.410000 858.500000 275.590000 ;
      RECT 816.500000 274.410000 849.500000 275.590000 ;
      RECT 807.500000 274.410000 808.500000 275.590000 ;
      RECT 766.500000 274.410000 799.500000 275.590000 ;
      RECT 757.500000 274.410000 758.500000 275.590000 ;
      RECT 716.500000 274.410000 749.500000 275.590000 ;
      RECT 707.500000 274.410000 708.500000 275.590000 ;
      RECT 666.500000 274.410000 699.500000 275.590000 ;
      RECT 657.500000 274.410000 658.500000 275.590000 ;
      RECT 616.500000 274.410000 649.500000 275.590000 ;
      RECT 607.500000 274.410000 608.500000 275.590000 ;
      RECT 566.500000 274.410000 599.500000 275.590000 ;
      RECT 557.500000 274.410000 558.500000 275.590000 ;
      RECT 516.500000 274.410000 549.500000 275.590000 ;
      RECT 507.500000 274.410000 508.500000 275.590000 ;
      RECT 466.500000 274.410000 499.500000 275.590000 ;
      RECT 457.500000 274.410000 458.500000 275.590000 ;
      RECT 416.500000 274.410000 449.500000 275.590000 ;
      RECT 407.500000 274.410000 408.500000 275.590000 ;
      RECT 366.500000 274.410000 399.500000 275.590000 ;
      RECT 357.500000 274.410000 358.500000 275.590000 ;
      RECT 316.500000 274.410000 349.500000 275.590000 ;
      RECT 307.500000 274.410000 308.500000 275.590000 ;
      RECT 266.500000 274.410000 299.500000 275.590000 ;
      RECT 257.500000 274.410000 258.500000 275.590000 ;
      RECT 216.500000 274.410000 249.500000 275.590000 ;
      RECT 207.500000 274.410000 208.500000 275.590000 ;
      RECT 166.500000 274.410000 199.500000 275.590000 ;
      RECT 157.500000 274.410000 158.500000 275.590000 ;
      RECT 116.500000 274.410000 149.500000 275.590000 ;
      RECT 107.500000 274.410000 108.500000 275.590000 ;
      RECT 66.500000 274.410000 99.500000 275.590000 ;
      RECT 57.500000 274.410000 58.500000 275.590000 ;
      RECT 29.500000 274.410000 49.500000 275.590000 ;
      RECT 15.500000 274.410000 16.500000 275.590000 ;
      RECT 1157.500000 273.590000 1170.500000 274.410000 ;
      RECT 1107.500000 273.590000 1149.500000 274.410000 ;
      RECT 1057.500000 273.590000 1099.500000 274.410000 ;
      RECT 1007.500000 273.590000 1049.500000 274.410000 ;
      RECT 957.500000 273.590000 999.500000 274.410000 ;
      RECT 907.500000 273.590000 949.500000 274.410000 ;
      RECT 857.500000 273.590000 899.500000 274.410000 ;
      RECT 807.500000 273.590000 849.500000 274.410000 ;
      RECT 757.500000 273.590000 799.500000 274.410000 ;
      RECT 707.500000 273.590000 749.500000 274.410000 ;
      RECT 657.500000 273.590000 699.500000 274.410000 ;
      RECT 607.500000 273.590000 649.500000 274.410000 ;
      RECT 557.500000 273.590000 599.500000 274.410000 ;
      RECT 507.500000 273.590000 549.500000 274.410000 ;
      RECT 457.500000 273.590000 499.500000 274.410000 ;
      RECT 407.500000 273.590000 449.500000 274.410000 ;
      RECT 357.500000 273.590000 399.500000 274.410000 ;
      RECT 307.500000 273.590000 349.500000 274.410000 ;
      RECT 257.500000 273.590000 299.500000 274.410000 ;
      RECT 207.500000 273.590000 249.500000 274.410000 ;
      RECT 157.500000 273.590000 199.500000 274.410000 ;
      RECT 107.500000 273.590000 149.500000 274.410000 ;
      RECT 57.500000 273.590000 99.500000 274.410000 ;
      RECT 15.500000 273.590000 49.500000 274.410000 ;
      RECT 1183.500000 272.410000 1186.000000 275.590000 ;
      RECT 1169.500000 272.410000 1170.500000 273.590000 ;
      RECT 1116.500000 272.410000 1149.500000 273.590000 ;
      RECT 1107.500000 272.410000 1108.500000 273.590000 ;
      RECT 1066.500000 272.410000 1099.500000 273.590000 ;
      RECT 1057.500000 272.410000 1058.500000 273.590000 ;
      RECT 1016.500000 272.410000 1049.500000 273.590000 ;
      RECT 1007.500000 272.410000 1008.500000 273.590000 ;
      RECT 966.500000 272.410000 999.500000 273.590000 ;
      RECT 957.500000 272.410000 958.500000 273.590000 ;
      RECT 916.500000 272.410000 949.500000 273.590000 ;
      RECT 907.500000 272.410000 908.500000 273.590000 ;
      RECT 866.500000 272.410000 899.500000 273.590000 ;
      RECT 857.500000 272.410000 858.500000 273.590000 ;
      RECT 816.500000 272.410000 849.500000 273.590000 ;
      RECT 807.500000 272.410000 808.500000 273.590000 ;
      RECT 766.500000 272.410000 799.500000 273.590000 ;
      RECT 757.500000 272.410000 758.500000 273.590000 ;
      RECT 716.500000 272.410000 749.500000 273.590000 ;
      RECT 707.500000 272.410000 708.500000 273.590000 ;
      RECT 666.500000 272.410000 699.500000 273.590000 ;
      RECT 657.500000 272.410000 658.500000 273.590000 ;
      RECT 616.500000 272.410000 649.500000 273.590000 ;
      RECT 607.500000 272.410000 608.500000 273.590000 ;
      RECT 566.500000 272.410000 599.500000 273.590000 ;
      RECT 557.500000 272.410000 558.500000 273.590000 ;
      RECT 516.500000 272.410000 549.500000 273.590000 ;
      RECT 507.500000 272.410000 508.500000 273.590000 ;
      RECT 466.500000 272.410000 499.500000 273.590000 ;
      RECT 457.500000 272.410000 458.500000 273.590000 ;
      RECT 416.500000 272.410000 449.500000 273.590000 ;
      RECT 407.500000 272.410000 408.500000 273.590000 ;
      RECT 366.500000 272.410000 399.500000 273.590000 ;
      RECT 357.500000 272.410000 358.500000 273.590000 ;
      RECT 316.500000 272.410000 349.500000 273.590000 ;
      RECT 307.500000 272.410000 308.500000 273.590000 ;
      RECT 266.500000 272.410000 299.500000 273.590000 ;
      RECT 257.500000 272.410000 258.500000 273.590000 ;
      RECT 216.500000 272.410000 249.500000 273.590000 ;
      RECT 207.500000 272.410000 208.500000 273.590000 ;
      RECT 166.500000 272.410000 199.500000 273.590000 ;
      RECT 157.500000 272.410000 158.500000 273.590000 ;
      RECT 116.500000 272.410000 149.500000 273.590000 ;
      RECT 107.500000 272.410000 108.500000 273.590000 ;
      RECT 66.500000 272.410000 99.500000 273.590000 ;
      RECT 57.500000 272.410000 58.500000 273.590000 ;
      RECT 29.500000 272.410000 49.500000 273.590000 ;
      RECT 15.500000 272.410000 16.500000 273.590000 ;
      RECT 0.000000 272.410000 2.500000 275.590000 ;
      RECT 1169.500000 271.590000 1186.000000 272.410000 ;
      RECT 1116.500000 271.590000 1156.500000 272.410000 ;
      RECT 1066.500000 271.590000 1108.500000 272.410000 ;
      RECT 1016.500000 271.590000 1058.500000 272.410000 ;
      RECT 966.500000 271.590000 1008.500000 272.410000 ;
      RECT 916.500000 271.590000 958.500000 272.410000 ;
      RECT 866.500000 271.590000 908.500000 272.410000 ;
      RECT 816.500000 271.590000 858.500000 272.410000 ;
      RECT 766.500000 271.590000 808.500000 272.410000 ;
      RECT 716.500000 271.590000 758.500000 272.410000 ;
      RECT 666.500000 271.590000 708.500000 272.410000 ;
      RECT 616.500000 271.590000 658.500000 272.410000 ;
      RECT 566.500000 271.590000 608.500000 272.410000 ;
      RECT 516.500000 271.590000 558.500000 272.410000 ;
      RECT 466.500000 271.590000 508.500000 272.410000 ;
      RECT 416.500000 271.590000 458.500000 272.410000 ;
      RECT 366.500000 271.590000 408.500000 272.410000 ;
      RECT 316.500000 271.590000 358.500000 272.410000 ;
      RECT 266.500000 271.590000 308.500000 272.410000 ;
      RECT 216.500000 271.590000 258.500000 272.410000 ;
      RECT 166.500000 271.590000 208.500000 272.410000 ;
      RECT 116.500000 271.590000 158.500000 272.410000 ;
      RECT 66.500000 271.590000 108.500000 272.410000 ;
      RECT 29.500000 271.590000 58.500000 272.410000 ;
      RECT 0.000000 271.590000 16.500000 272.410000 ;
      RECT 1169.500000 270.410000 1170.500000 271.590000 ;
      RECT 1116.500000 270.410000 1149.500000 271.590000 ;
      RECT 1107.500000 270.410000 1108.500000 271.590000 ;
      RECT 1066.500000 270.410000 1099.500000 271.590000 ;
      RECT 1057.500000 270.410000 1058.500000 271.590000 ;
      RECT 1016.500000 270.410000 1049.500000 271.590000 ;
      RECT 1007.500000 270.410000 1008.500000 271.590000 ;
      RECT 966.500000 270.410000 999.500000 271.590000 ;
      RECT 957.500000 270.410000 958.500000 271.590000 ;
      RECT 916.500000 270.410000 949.500000 271.590000 ;
      RECT 907.500000 270.410000 908.500000 271.590000 ;
      RECT 866.500000 270.410000 899.500000 271.590000 ;
      RECT 857.500000 270.410000 858.500000 271.590000 ;
      RECT 816.500000 270.410000 849.500000 271.590000 ;
      RECT 807.500000 270.410000 808.500000 271.590000 ;
      RECT 766.500000 270.410000 799.500000 271.590000 ;
      RECT 757.500000 270.410000 758.500000 271.590000 ;
      RECT 716.500000 270.410000 749.500000 271.590000 ;
      RECT 707.500000 270.410000 708.500000 271.590000 ;
      RECT 666.500000 270.410000 699.500000 271.590000 ;
      RECT 657.500000 270.410000 658.500000 271.590000 ;
      RECT 616.500000 270.410000 649.500000 271.590000 ;
      RECT 607.500000 270.410000 608.500000 271.590000 ;
      RECT 566.500000 270.410000 599.500000 271.590000 ;
      RECT 557.500000 270.410000 558.500000 271.590000 ;
      RECT 516.500000 270.410000 549.500000 271.590000 ;
      RECT 507.500000 270.410000 508.500000 271.590000 ;
      RECT 466.500000 270.410000 499.500000 271.590000 ;
      RECT 457.500000 270.410000 458.500000 271.590000 ;
      RECT 416.500000 270.410000 449.500000 271.590000 ;
      RECT 407.500000 270.410000 408.500000 271.590000 ;
      RECT 366.500000 270.410000 399.500000 271.590000 ;
      RECT 357.500000 270.410000 358.500000 271.590000 ;
      RECT 316.500000 270.410000 349.500000 271.590000 ;
      RECT 307.500000 270.410000 308.500000 271.590000 ;
      RECT 266.500000 270.410000 299.500000 271.590000 ;
      RECT 257.500000 270.410000 258.500000 271.590000 ;
      RECT 216.500000 270.410000 249.500000 271.590000 ;
      RECT 207.500000 270.410000 208.500000 271.590000 ;
      RECT 166.500000 270.410000 199.500000 271.590000 ;
      RECT 157.500000 270.410000 158.500000 271.590000 ;
      RECT 116.500000 270.410000 149.500000 271.590000 ;
      RECT 107.500000 270.410000 108.500000 271.590000 ;
      RECT 66.500000 270.410000 99.500000 271.590000 ;
      RECT 57.500000 270.410000 58.500000 271.590000 ;
      RECT 29.500000 270.410000 49.500000 271.590000 ;
      RECT 15.500000 270.410000 16.500000 271.590000 ;
      RECT 1157.500000 269.590000 1170.500000 270.410000 ;
      RECT 1107.500000 269.590000 1149.500000 270.410000 ;
      RECT 1057.500000 269.590000 1099.500000 270.410000 ;
      RECT 1007.500000 269.590000 1049.500000 270.410000 ;
      RECT 957.500000 269.590000 999.500000 270.410000 ;
      RECT 907.500000 269.590000 949.500000 270.410000 ;
      RECT 857.500000 269.590000 899.500000 270.410000 ;
      RECT 807.500000 269.590000 849.500000 270.410000 ;
      RECT 757.500000 269.590000 799.500000 270.410000 ;
      RECT 707.500000 269.590000 749.500000 270.410000 ;
      RECT 657.500000 269.590000 699.500000 270.410000 ;
      RECT 607.500000 269.590000 649.500000 270.410000 ;
      RECT 557.500000 269.590000 599.500000 270.410000 ;
      RECT 507.500000 269.590000 549.500000 270.410000 ;
      RECT 457.500000 269.590000 499.500000 270.410000 ;
      RECT 407.500000 269.590000 449.500000 270.410000 ;
      RECT 357.500000 269.590000 399.500000 270.410000 ;
      RECT 307.500000 269.590000 349.500000 270.410000 ;
      RECT 257.500000 269.590000 299.500000 270.410000 ;
      RECT 207.500000 269.590000 249.500000 270.410000 ;
      RECT 157.500000 269.590000 199.500000 270.410000 ;
      RECT 107.500000 269.590000 149.500000 270.410000 ;
      RECT 57.500000 269.590000 99.500000 270.410000 ;
      RECT 15.500000 269.590000 49.500000 270.410000 ;
      RECT 1183.500000 268.410000 1186.000000 271.590000 ;
      RECT 1169.500000 268.410000 1170.500000 269.590000 ;
      RECT 1116.500000 268.410000 1149.500000 269.590000 ;
      RECT 1107.500000 268.410000 1108.500000 269.590000 ;
      RECT 1066.500000 268.410000 1099.500000 269.590000 ;
      RECT 1057.500000 268.410000 1058.500000 269.590000 ;
      RECT 1016.500000 268.410000 1049.500000 269.590000 ;
      RECT 1007.500000 268.410000 1008.500000 269.590000 ;
      RECT 966.500000 268.410000 999.500000 269.590000 ;
      RECT 957.500000 268.410000 958.500000 269.590000 ;
      RECT 916.500000 268.410000 949.500000 269.590000 ;
      RECT 907.500000 268.410000 908.500000 269.590000 ;
      RECT 866.500000 268.410000 899.500000 269.590000 ;
      RECT 857.500000 268.410000 858.500000 269.590000 ;
      RECT 816.500000 268.410000 849.500000 269.590000 ;
      RECT 807.500000 268.410000 808.500000 269.590000 ;
      RECT 766.500000 268.410000 799.500000 269.590000 ;
      RECT 757.500000 268.410000 758.500000 269.590000 ;
      RECT 716.500000 268.410000 749.500000 269.590000 ;
      RECT 707.500000 268.410000 708.500000 269.590000 ;
      RECT 666.500000 268.410000 699.500000 269.590000 ;
      RECT 657.500000 268.410000 658.500000 269.590000 ;
      RECT 616.500000 268.410000 649.500000 269.590000 ;
      RECT 607.500000 268.410000 608.500000 269.590000 ;
      RECT 566.500000 268.410000 599.500000 269.590000 ;
      RECT 557.500000 268.410000 558.500000 269.590000 ;
      RECT 516.500000 268.410000 549.500000 269.590000 ;
      RECT 507.500000 268.410000 508.500000 269.590000 ;
      RECT 466.500000 268.410000 499.500000 269.590000 ;
      RECT 457.500000 268.410000 458.500000 269.590000 ;
      RECT 416.500000 268.410000 449.500000 269.590000 ;
      RECT 407.500000 268.410000 408.500000 269.590000 ;
      RECT 366.500000 268.410000 399.500000 269.590000 ;
      RECT 357.500000 268.410000 358.500000 269.590000 ;
      RECT 316.500000 268.410000 349.500000 269.590000 ;
      RECT 307.500000 268.410000 308.500000 269.590000 ;
      RECT 266.500000 268.410000 299.500000 269.590000 ;
      RECT 257.500000 268.410000 258.500000 269.590000 ;
      RECT 216.500000 268.410000 249.500000 269.590000 ;
      RECT 207.500000 268.410000 208.500000 269.590000 ;
      RECT 166.500000 268.410000 199.500000 269.590000 ;
      RECT 157.500000 268.410000 158.500000 269.590000 ;
      RECT 116.500000 268.410000 149.500000 269.590000 ;
      RECT 107.500000 268.410000 108.500000 269.590000 ;
      RECT 66.500000 268.410000 99.500000 269.590000 ;
      RECT 57.500000 268.410000 58.500000 269.590000 ;
      RECT 29.500000 268.410000 49.500000 269.590000 ;
      RECT 15.500000 268.410000 16.500000 269.590000 ;
      RECT 0.000000 268.410000 2.500000 271.590000 ;
      RECT 1169.500000 267.590000 1186.000000 268.410000 ;
      RECT 1116.500000 267.590000 1156.500000 268.410000 ;
      RECT 1066.500000 267.590000 1108.500000 268.410000 ;
      RECT 1016.500000 267.590000 1058.500000 268.410000 ;
      RECT 966.500000 267.590000 1008.500000 268.410000 ;
      RECT 916.500000 267.590000 958.500000 268.410000 ;
      RECT 866.500000 267.590000 908.500000 268.410000 ;
      RECT 816.500000 267.590000 858.500000 268.410000 ;
      RECT 766.500000 267.590000 808.500000 268.410000 ;
      RECT 716.500000 267.590000 758.500000 268.410000 ;
      RECT 666.500000 267.590000 708.500000 268.410000 ;
      RECT 616.500000 267.590000 658.500000 268.410000 ;
      RECT 566.500000 267.590000 608.500000 268.410000 ;
      RECT 516.500000 267.590000 558.500000 268.410000 ;
      RECT 466.500000 267.590000 508.500000 268.410000 ;
      RECT 416.500000 267.590000 458.500000 268.410000 ;
      RECT 366.500000 267.590000 408.500000 268.410000 ;
      RECT 316.500000 267.590000 358.500000 268.410000 ;
      RECT 266.500000 267.590000 308.500000 268.410000 ;
      RECT 216.500000 267.590000 258.500000 268.410000 ;
      RECT 166.500000 267.590000 208.500000 268.410000 ;
      RECT 116.500000 267.590000 158.500000 268.410000 ;
      RECT 66.500000 267.590000 108.500000 268.410000 ;
      RECT 29.500000 267.590000 58.500000 268.410000 ;
      RECT 0.000000 267.590000 16.500000 268.410000 ;
      RECT 1169.500000 266.410000 1170.500000 267.590000 ;
      RECT 1116.500000 266.410000 1149.500000 267.590000 ;
      RECT 1107.500000 266.410000 1108.500000 267.590000 ;
      RECT 1066.500000 266.410000 1099.500000 267.590000 ;
      RECT 1057.500000 266.410000 1058.500000 267.590000 ;
      RECT 1016.500000 266.410000 1049.500000 267.590000 ;
      RECT 1007.500000 266.410000 1008.500000 267.590000 ;
      RECT 966.500000 266.410000 999.500000 267.590000 ;
      RECT 957.500000 266.410000 958.500000 267.590000 ;
      RECT 916.500000 266.410000 949.500000 267.590000 ;
      RECT 907.500000 266.410000 908.500000 267.590000 ;
      RECT 866.500000 266.410000 899.500000 267.590000 ;
      RECT 857.500000 266.410000 858.500000 267.590000 ;
      RECT 816.500000 266.410000 849.500000 267.590000 ;
      RECT 807.500000 266.410000 808.500000 267.590000 ;
      RECT 766.500000 266.410000 799.500000 267.590000 ;
      RECT 757.500000 266.410000 758.500000 267.590000 ;
      RECT 716.500000 266.410000 749.500000 267.590000 ;
      RECT 707.500000 266.410000 708.500000 267.590000 ;
      RECT 666.500000 266.410000 699.500000 267.590000 ;
      RECT 657.500000 266.410000 658.500000 267.590000 ;
      RECT 616.500000 266.410000 649.500000 267.590000 ;
      RECT 607.500000 266.410000 608.500000 267.590000 ;
      RECT 566.500000 266.410000 599.500000 267.590000 ;
      RECT 557.500000 266.410000 558.500000 267.590000 ;
      RECT 516.500000 266.410000 549.500000 267.590000 ;
      RECT 507.500000 266.410000 508.500000 267.590000 ;
      RECT 466.500000 266.410000 499.500000 267.590000 ;
      RECT 457.500000 266.410000 458.500000 267.590000 ;
      RECT 416.500000 266.410000 449.500000 267.590000 ;
      RECT 407.500000 266.410000 408.500000 267.590000 ;
      RECT 366.500000 266.410000 399.500000 267.590000 ;
      RECT 357.500000 266.410000 358.500000 267.590000 ;
      RECT 316.500000 266.410000 349.500000 267.590000 ;
      RECT 307.500000 266.410000 308.500000 267.590000 ;
      RECT 266.500000 266.410000 299.500000 267.590000 ;
      RECT 257.500000 266.410000 258.500000 267.590000 ;
      RECT 216.500000 266.410000 249.500000 267.590000 ;
      RECT 207.500000 266.410000 208.500000 267.590000 ;
      RECT 166.500000 266.410000 199.500000 267.590000 ;
      RECT 157.500000 266.410000 158.500000 267.590000 ;
      RECT 116.500000 266.410000 149.500000 267.590000 ;
      RECT 107.500000 266.410000 108.500000 267.590000 ;
      RECT 66.500000 266.410000 99.500000 267.590000 ;
      RECT 57.500000 266.410000 58.500000 267.590000 ;
      RECT 29.500000 266.410000 49.500000 267.590000 ;
      RECT 15.500000 266.410000 16.500000 267.590000 ;
      RECT 1157.500000 265.590000 1170.500000 266.410000 ;
      RECT 1107.500000 265.590000 1149.500000 266.410000 ;
      RECT 1057.500000 265.590000 1099.500000 266.410000 ;
      RECT 1007.500000 265.590000 1049.500000 266.410000 ;
      RECT 957.500000 265.590000 999.500000 266.410000 ;
      RECT 907.500000 265.590000 949.500000 266.410000 ;
      RECT 857.500000 265.590000 899.500000 266.410000 ;
      RECT 807.500000 265.590000 849.500000 266.410000 ;
      RECT 757.500000 265.590000 799.500000 266.410000 ;
      RECT 707.500000 265.590000 749.500000 266.410000 ;
      RECT 657.500000 265.590000 699.500000 266.410000 ;
      RECT 607.500000 265.590000 649.500000 266.410000 ;
      RECT 557.500000 265.590000 599.500000 266.410000 ;
      RECT 507.500000 265.590000 549.500000 266.410000 ;
      RECT 457.500000 265.590000 499.500000 266.410000 ;
      RECT 407.500000 265.590000 449.500000 266.410000 ;
      RECT 357.500000 265.590000 399.500000 266.410000 ;
      RECT 307.500000 265.590000 349.500000 266.410000 ;
      RECT 257.500000 265.590000 299.500000 266.410000 ;
      RECT 207.500000 265.590000 249.500000 266.410000 ;
      RECT 157.500000 265.590000 199.500000 266.410000 ;
      RECT 107.500000 265.590000 149.500000 266.410000 ;
      RECT 57.500000 265.590000 99.500000 266.410000 ;
      RECT 15.500000 265.590000 49.500000 266.410000 ;
      RECT 1183.500000 264.410000 1186.000000 267.590000 ;
      RECT 1169.500000 264.410000 1170.500000 265.590000 ;
      RECT 1116.500000 264.410000 1149.500000 265.590000 ;
      RECT 1107.500000 264.410000 1108.500000 265.590000 ;
      RECT 1066.500000 264.410000 1099.500000 265.590000 ;
      RECT 1057.500000 264.410000 1058.500000 265.590000 ;
      RECT 1016.500000 264.410000 1049.500000 265.590000 ;
      RECT 1007.500000 264.410000 1008.500000 265.590000 ;
      RECT 966.500000 264.410000 999.500000 265.590000 ;
      RECT 957.500000 264.410000 958.500000 265.590000 ;
      RECT 916.500000 264.410000 949.500000 265.590000 ;
      RECT 907.500000 264.410000 908.500000 265.590000 ;
      RECT 866.500000 264.410000 899.500000 265.590000 ;
      RECT 857.500000 264.410000 858.500000 265.590000 ;
      RECT 816.500000 264.410000 849.500000 265.590000 ;
      RECT 807.500000 264.410000 808.500000 265.590000 ;
      RECT 766.500000 264.410000 799.500000 265.590000 ;
      RECT 757.500000 264.410000 758.500000 265.590000 ;
      RECT 716.500000 264.410000 749.500000 265.590000 ;
      RECT 707.500000 264.410000 708.500000 265.590000 ;
      RECT 666.500000 264.410000 699.500000 265.590000 ;
      RECT 657.500000 264.410000 658.500000 265.590000 ;
      RECT 616.500000 264.410000 649.500000 265.590000 ;
      RECT 607.500000 264.410000 608.500000 265.590000 ;
      RECT 566.500000 264.410000 599.500000 265.590000 ;
      RECT 557.500000 264.410000 558.500000 265.590000 ;
      RECT 516.500000 264.410000 549.500000 265.590000 ;
      RECT 507.500000 264.410000 508.500000 265.590000 ;
      RECT 466.500000 264.410000 499.500000 265.590000 ;
      RECT 457.500000 264.410000 458.500000 265.590000 ;
      RECT 416.500000 264.410000 449.500000 265.590000 ;
      RECT 407.500000 264.410000 408.500000 265.590000 ;
      RECT 366.500000 264.410000 399.500000 265.590000 ;
      RECT 357.500000 264.410000 358.500000 265.590000 ;
      RECT 316.500000 264.410000 349.500000 265.590000 ;
      RECT 307.500000 264.410000 308.500000 265.590000 ;
      RECT 266.500000 264.410000 299.500000 265.590000 ;
      RECT 257.500000 264.410000 258.500000 265.590000 ;
      RECT 216.500000 264.410000 249.500000 265.590000 ;
      RECT 207.500000 264.410000 208.500000 265.590000 ;
      RECT 166.500000 264.410000 199.500000 265.590000 ;
      RECT 157.500000 264.410000 158.500000 265.590000 ;
      RECT 116.500000 264.410000 149.500000 265.590000 ;
      RECT 107.500000 264.410000 108.500000 265.590000 ;
      RECT 66.500000 264.410000 99.500000 265.590000 ;
      RECT 57.500000 264.410000 58.500000 265.590000 ;
      RECT 29.500000 264.410000 49.500000 265.590000 ;
      RECT 15.500000 264.410000 16.500000 265.590000 ;
      RECT 0.000000 264.410000 2.500000 267.590000 ;
      RECT 1169.500000 263.590000 1186.000000 264.410000 ;
      RECT 1116.500000 263.590000 1156.500000 264.410000 ;
      RECT 1066.500000 263.590000 1108.500000 264.410000 ;
      RECT 1016.500000 263.590000 1058.500000 264.410000 ;
      RECT 966.500000 263.590000 1008.500000 264.410000 ;
      RECT 916.500000 263.590000 958.500000 264.410000 ;
      RECT 866.500000 263.590000 908.500000 264.410000 ;
      RECT 816.500000 263.590000 858.500000 264.410000 ;
      RECT 766.500000 263.590000 808.500000 264.410000 ;
      RECT 716.500000 263.590000 758.500000 264.410000 ;
      RECT 666.500000 263.590000 708.500000 264.410000 ;
      RECT 616.500000 263.590000 658.500000 264.410000 ;
      RECT 566.500000 263.590000 608.500000 264.410000 ;
      RECT 516.500000 263.590000 558.500000 264.410000 ;
      RECT 466.500000 263.590000 508.500000 264.410000 ;
      RECT 416.500000 263.590000 458.500000 264.410000 ;
      RECT 366.500000 263.590000 408.500000 264.410000 ;
      RECT 316.500000 263.590000 358.500000 264.410000 ;
      RECT 266.500000 263.590000 308.500000 264.410000 ;
      RECT 216.500000 263.590000 258.500000 264.410000 ;
      RECT 166.500000 263.590000 208.500000 264.410000 ;
      RECT 116.500000 263.590000 158.500000 264.410000 ;
      RECT 66.500000 263.590000 108.500000 264.410000 ;
      RECT 29.500000 263.590000 58.500000 264.410000 ;
      RECT 0.000000 263.590000 16.500000 264.410000 ;
      RECT 1169.500000 262.410000 1170.500000 263.590000 ;
      RECT 1116.500000 262.410000 1149.500000 263.590000 ;
      RECT 1107.500000 262.410000 1108.500000 263.590000 ;
      RECT 1066.500000 262.410000 1099.500000 263.590000 ;
      RECT 1057.500000 262.410000 1058.500000 263.590000 ;
      RECT 1016.500000 262.410000 1049.500000 263.590000 ;
      RECT 1007.500000 262.410000 1008.500000 263.590000 ;
      RECT 966.500000 262.410000 999.500000 263.590000 ;
      RECT 957.500000 262.410000 958.500000 263.590000 ;
      RECT 916.500000 262.410000 949.500000 263.590000 ;
      RECT 907.500000 262.410000 908.500000 263.590000 ;
      RECT 866.500000 262.410000 899.500000 263.590000 ;
      RECT 857.500000 262.410000 858.500000 263.590000 ;
      RECT 816.500000 262.410000 849.500000 263.590000 ;
      RECT 807.500000 262.410000 808.500000 263.590000 ;
      RECT 766.500000 262.410000 799.500000 263.590000 ;
      RECT 757.500000 262.410000 758.500000 263.590000 ;
      RECT 716.500000 262.410000 749.500000 263.590000 ;
      RECT 707.500000 262.410000 708.500000 263.590000 ;
      RECT 666.500000 262.410000 699.500000 263.590000 ;
      RECT 657.500000 262.410000 658.500000 263.590000 ;
      RECT 616.500000 262.410000 649.500000 263.590000 ;
      RECT 607.500000 262.410000 608.500000 263.590000 ;
      RECT 566.500000 262.410000 599.500000 263.590000 ;
      RECT 557.500000 262.410000 558.500000 263.590000 ;
      RECT 516.500000 262.410000 549.500000 263.590000 ;
      RECT 507.500000 262.410000 508.500000 263.590000 ;
      RECT 466.500000 262.410000 499.500000 263.590000 ;
      RECT 457.500000 262.410000 458.500000 263.590000 ;
      RECT 416.500000 262.410000 449.500000 263.590000 ;
      RECT 407.500000 262.410000 408.500000 263.590000 ;
      RECT 366.500000 262.410000 399.500000 263.590000 ;
      RECT 357.500000 262.410000 358.500000 263.590000 ;
      RECT 316.500000 262.410000 349.500000 263.590000 ;
      RECT 307.500000 262.410000 308.500000 263.590000 ;
      RECT 266.500000 262.410000 299.500000 263.590000 ;
      RECT 257.500000 262.410000 258.500000 263.590000 ;
      RECT 216.500000 262.410000 249.500000 263.590000 ;
      RECT 207.500000 262.410000 208.500000 263.590000 ;
      RECT 166.500000 262.410000 199.500000 263.590000 ;
      RECT 157.500000 262.410000 158.500000 263.590000 ;
      RECT 116.500000 262.410000 149.500000 263.590000 ;
      RECT 107.500000 262.410000 108.500000 263.590000 ;
      RECT 66.500000 262.410000 99.500000 263.590000 ;
      RECT 57.500000 262.410000 58.500000 263.590000 ;
      RECT 29.500000 262.410000 49.500000 263.590000 ;
      RECT 15.500000 262.410000 16.500000 263.590000 ;
      RECT 1157.500000 261.590000 1170.500000 262.410000 ;
      RECT 1107.500000 261.590000 1149.500000 262.410000 ;
      RECT 1057.500000 261.590000 1099.500000 262.410000 ;
      RECT 1007.500000 261.590000 1049.500000 262.410000 ;
      RECT 957.500000 261.590000 999.500000 262.410000 ;
      RECT 907.500000 261.590000 949.500000 262.410000 ;
      RECT 857.500000 261.590000 899.500000 262.410000 ;
      RECT 807.500000 261.590000 849.500000 262.410000 ;
      RECT 757.500000 261.590000 799.500000 262.410000 ;
      RECT 707.500000 261.590000 749.500000 262.410000 ;
      RECT 657.500000 261.590000 699.500000 262.410000 ;
      RECT 607.500000 261.590000 649.500000 262.410000 ;
      RECT 557.500000 261.590000 599.500000 262.410000 ;
      RECT 507.500000 261.590000 549.500000 262.410000 ;
      RECT 457.500000 261.590000 499.500000 262.410000 ;
      RECT 407.500000 261.590000 449.500000 262.410000 ;
      RECT 357.500000 261.590000 399.500000 262.410000 ;
      RECT 307.500000 261.590000 349.500000 262.410000 ;
      RECT 257.500000 261.590000 299.500000 262.410000 ;
      RECT 207.500000 261.590000 249.500000 262.410000 ;
      RECT 157.500000 261.590000 199.500000 262.410000 ;
      RECT 107.500000 261.590000 149.500000 262.410000 ;
      RECT 57.500000 261.590000 99.500000 262.410000 ;
      RECT 15.500000 261.590000 49.500000 262.410000 ;
      RECT 1183.500000 260.410000 1186.000000 263.590000 ;
      RECT 1169.500000 260.410000 1170.500000 261.590000 ;
      RECT 1116.500000 260.410000 1149.500000 261.590000 ;
      RECT 1107.500000 260.410000 1108.500000 261.590000 ;
      RECT 1066.500000 260.410000 1099.500000 261.590000 ;
      RECT 1057.500000 260.410000 1058.500000 261.590000 ;
      RECT 1016.500000 260.410000 1049.500000 261.590000 ;
      RECT 1007.500000 260.410000 1008.500000 261.590000 ;
      RECT 966.500000 260.410000 999.500000 261.590000 ;
      RECT 957.500000 260.410000 958.500000 261.590000 ;
      RECT 916.500000 260.410000 949.500000 261.590000 ;
      RECT 907.500000 260.410000 908.500000 261.590000 ;
      RECT 866.500000 260.410000 899.500000 261.590000 ;
      RECT 857.500000 260.410000 858.500000 261.590000 ;
      RECT 816.500000 260.410000 849.500000 261.590000 ;
      RECT 807.500000 260.410000 808.500000 261.590000 ;
      RECT 766.500000 260.410000 799.500000 261.590000 ;
      RECT 757.500000 260.410000 758.500000 261.590000 ;
      RECT 716.500000 260.410000 749.500000 261.590000 ;
      RECT 707.500000 260.410000 708.500000 261.590000 ;
      RECT 666.500000 260.410000 699.500000 261.590000 ;
      RECT 657.500000 260.410000 658.500000 261.590000 ;
      RECT 616.500000 260.410000 649.500000 261.590000 ;
      RECT 607.500000 260.410000 608.500000 261.590000 ;
      RECT 566.500000 260.410000 599.500000 261.590000 ;
      RECT 557.500000 260.410000 558.500000 261.590000 ;
      RECT 516.500000 260.410000 549.500000 261.590000 ;
      RECT 507.500000 260.410000 508.500000 261.590000 ;
      RECT 466.500000 260.410000 499.500000 261.590000 ;
      RECT 457.500000 260.410000 458.500000 261.590000 ;
      RECT 416.500000 260.410000 449.500000 261.590000 ;
      RECT 407.500000 260.410000 408.500000 261.590000 ;
      RECT 366.500000 260.410000 399.500000 261.590000 ;
      RECT 357.500000 260.410000 358.500000 261.590000 ;
      RECT 316.500000 260.410000 349.500000 261.590000 ;
      RECT 307.500000 260.410000 308.500000 261.590000 ;
      RECT 266.500000 260.410000 299.500000 261.590000 ;
      RECT 257.500000 260.410000 258.500000 261.590000 ;
      RECT 216.500000 260.410000 249.500000 261.590000 ;
      RECT 207.500000 260.410000 208.500000 261.590000 ;
      RECT 166.500000 260.410000 199.500000 261.590000 ;
      RECT 157.500000 260.410000 158.500000 261.590000 ;
      RECT 116.500000 260.410000 149.500000 261.590000 ;
      RECT 107.500000 260.410000 108.500000 261.590000 ;
      RECT 66.500000 260.410000 99.500000 261.590000 ;
      RECT 57.500000 260.410000 58.500000 261.590000 ;
      RECT 29.500000 260.410000 49.500000 261.590000 ;
      RECT 15.500000 260.410000 16.500000 261.590000 ;
      RECT 0.000000 260.410000 2.500000 263.590000 ;
      RECT 1169.500000 259.590000 1186.000000 260.410000 ;
      RECT 1116.500000 259.590000 1156.500000 260.410000 ;
      RECT 1169.500000 258.410000 1170.500000 259.590000 ;
      RECT 1116.500000 258.410000 1149.500000 259.590000 ;
      RECT 1066.500000 258.410000 1108.500000 260.410000 ;
      RECT 1016.500000 258.410000 1058.500000 260.410000 ;
      RECT 966.500000 258.410000 1008.500000 260.410000 ;
      RECT 916.500000 258.410000 958.500000 260.410000 ;
      RECT 866.500000 258.410000 908.500000 260.410000 ;
      RECT 816.500000 258.410000 858.500000 260.410000 ;
      RECT 766.500000 258.410000 808.500000 260.410000 ;
      RECT 716.500000 258.410000 758.500000 260.410000 ;
      RECT 666.500000 258.410000 708.500000 260.410000 ;
      RECT 616.500000 258.410000 658.500000 260.410000 ;
      RECT 566.500000 258.410000 608.500000 260.410000 ;
      RECT 516.500000 258.410000 558.500000 260.410000 ;
      RECT 466.500000 258.410000 508.500000 260.410000 ;
      RECT 416.500000 258.410000 458.500000 260.410000 ;
      RECT 366.500000 258.410000 408.500000 260.410000 ;
      RECT 316.500000 258.410000 358.500000 260.410000 ;
      RECT 266.500000 258.410000 308.500000 260.410000 ;
      RECT 216.500000 258.410000 258.500000 260.410000 ;
      RECT 166.500000 258.410000 208.500000 260.410000 ;
      RECT 116.500000 258.410000 158.500000 260.410000 ;
      RECT 66.500000 258.410000 108.500000 260.410000 ;
      RECT 29.500000 258.410000 58.500000 260.410000 ;
      RECT 0.000000 258.410000 16.500000 260.410000 ;
      RECT 1157.500000 257.590000 1170.500000 258.410000 ;
      RECT 1183.500000 256.410000 1186.000000 259.590000 ;
      RECT 1169.500000 256.410000 1170.500000 257.590000 ;
      RECT 0.000000 256.410000 1149.500000 258.410000 ;
      RECT 1169.500000 255.590000 1186.000000 256.410000 ;
      RECT 1169.500000 254.410000 1170.500000 255.590000 ;
      RECT 0.000000 254.410000 1156.500000 256.410000 ;
      RECT 0.000000 253.590000 1170.500000 254.410000 ;
      RECT 1183.500000 252.410000 1186.000000 255.590000 ;
      RECT 1169.500000 252.410000 1170.500000 253.590000 ;
      RECT 1169.500000 251.590000 1186.000000 252.410000 ;
      RECT 1169.500000 250.410000 1170.500000 251.590000 ;
      RECT 0.000000 250.410000 1156.500000 253.590000 ;
      RECT 0.000000 249.590000 1170.500000 250.410000 ;
      RECT 1183.500000 248.410000 1186.000000 251.590000 ;
      RECT 1169.500000 248.410000 1170.500000 249.590000 ;
      RECT 1169.500000 247.590000 1186.000000 248.410000 ;
      RECT 1169.500000 246.410000 1170.500000 247.590000 ;
      RECT 0.000000 246.410000 1156.500000 249.590000 ;
      RECT 0.000000 245.590000 1170.500000 246.410000 ;
      RECT 1183.500000 244.410000 1186.000000 247.590000 ;
      RECT 1169.500000 244.410000 1170.500000 245.590000 ;
      RECT 1169.500000 243.590000 1186.000000 244.410000 ;
      RECT 1169.500000 242.410000 1170.500000 243.590000 ;
      RECT 0.000000 242.410000 1156.500000 245.590000 ;
      RECT 0.000000 241.590000 1170.500000 242.410000 ;
      RECT 1183.500000 240.410000 1186.000000 243.590000 ;
      RECT 1169.500000 240.410000 1170.500000 241.590000 ;
      RECT 1169.500000 239.590000 1186.000000 240.410000 ;
      RECT 1169.500000 238.410000 1170.500000 239.590000 ;
      RECT 0.000000 238.410000 1156.500000 241.590000 ;
      RECT 0.000000 237.590000 1170.500000 238.410000 ;
      RECT 1183.500000 236.410000 1186.000000 239.590000 ;
      RECT 1169.500000 236.410000 1170.500000 237.590000 ;
      RECT 1169.500000 235.590000 1186.000000 236.410000 ;
      RECT 1169.500000 234.410000 1170.500000 235.590000 ;
      RECT 0.000000 234.410000 1156.500000 237.590000 ;
      RECT 0.000000 233.590000 1170.500000 234.410000 ;
      RECT 1183.500000 232.410000 1186.000000 235.590000 ;
      RECT 1169.500000 232.410000 1170.500000 233.590000 ;
      RECT 1169.500000 231.590000 1186.000000 232.410000 ;
      RECT 1169.500000 230.410000 1170.500000 231.590000 ;
      RECT 0.000000 230.410000 1156.500000 233.590000 ;
      RECT 0.000000 229.590000 1170.500000 230.410000 ;
      RECT 1183.500000 228.410000 1186.000000 231.590000 ;
      RECT 1169.500000 228.410000 1170.500000 229.590000 ;
      RECT 1169.500000 227.590000 1186.000000 228.410000 ;
      RECT 1169.500000 226.410000 1170.500000 227.590000 ;
      RECT 0.000000 226.410000 1156.500000 229.590000 ;
      RECT 0.000000 225.590000 1170.500000 226.410000 ;
      RECT 1183.500000 224.410000 1186.000000 227.590000 ;
      RECT 1169.500000 224.410000 1170.500000 225.590000 ;
      RECT 1169.500000 223.590000 1186.000000 224.410000 ;
      RECT 0.000000 223.170000 1156.500000 225.590000 ;
      RECT 1183.500000 223.165000 1186.000000 223.590000 ;
      RECT 1169.500000 222.410000 1170.500000 223.590000 ;
      RECT 2.020000 222.410000 1156.500000 223.170000 ;
      RECT 2.020000 221.590000 1170.500000 222.410000 ;
      RECT 1183.500000 220.410000 1183.980000 223.165000 ;
      RECT 1169.500000 220.410000 1170.500000 221.590000 ;
      RECT 2.020000 220.070000 1156.500000 221.590000 ;
      RECT 1169.500000 220.065000 1183.980000 220.410000 ;
      RECT 1169.500000 219.590000 1186.000000 220.065000 ;
      RECT 1169.500000 218.410000 1170.500000 219.590000 ;
      RECT 0.000000 218.410000 1156.500000 220.070000 ;
      RECT 0.000000 217.590000 1170.500000 218.410000 ;
      RECT 1183.500000 217.485000 1186.000000 219.590000 ;
      RECT 1183.500000 216.410000 1183.980000 217.485000 ;
      RECT 1169.500000 216.410000 1170.500000 217.590000 ;
      RECT 1169.500000 215.590000 1183.980000 216.410000 ;
      RECT 1169.500000 214.410000 1170.500000 215.590000 ;
      RECT 0.000000 214.410000 1156.500000 217.590000 ;
      RECT 1183.500000 214.385000 1183.980000 215.590000 ;
      RECT 0.000000 213.590000 1170.500000 214.410000 ;
      RECT 1183.500000 213.525000 1186.000000 214.385000 ;
      RECT 0.000000 212.575000 1156.500000 213.590000 ;
      RECT 1183.500000 212.410000 1183.980000 213.525000 ;
      RECT 1169.500000 212.410000 1170.500000 213.590000 ;
      RECT 1169.500000 211.590000 1183.980000 212.410000 ;
      RECT 1183.500000 210.425000 1183.980000 211.590000 ;
      RECT 1169.500000 210.410000 1170.500000 211.590000 ;
      RECT 2.020000 210.410000 1156.500000 212.575000 ;
      RECT 2.020000 209.590000 1170.500000 210.410000 ;
      RECT 2.020000 209.475000 1156.500000 209.590000 ;
      RECT 0.000000 208.615000 1156.500000 209.475000 ;
      RECT 1183.500000 208.410000 1186.000000 210.425000 ;
      RECT 1169.500000 208.410000 1170.500000 209.590000 ;
      RECT 1169.500000 207.590000 1186.000000 208.410000 ;
      RECT 1169.500000 206.410000 1170.500000 207.590000 ;
      RECT 2.020000 206.410000 1156.500000 208.615000 ;
      RECT 2.020000 205.590000 1170.500000 206.410000 ;
      RECT 2.020000 205.515000 1156.500000 205.590000 ;
      RECT 1183.500000 204.410000 1186.000000 207.590000 ;
      RECT 1169.500000 204.410000 1170.500000 205.590000 ;
      RECT 1169.500000 203.590000 1186.000000 204.410000 ;
      RECT 0.000000 202.935000 1156.500000 205.515000 ;
      RECT 1183.500000 202.930000 1186.000000 203.590000 ;
      RECT 1169.500000 202.410000 1170.500000 203.590000 ;
      RECT 2.020000 202.410000 1156.500000 202.935000 ;
      RECT 2.020000 201.590000 1170.500000 202.410000 ;
      RECT 1183.500000 200.410000 1183.980000 202.930000 ;
      RECT 1169.500000 200.410000 1170.500000 201.590000 ;
      RECT 2.020000 199.835000 1156.500000 201.590000 ;
      RECT 1169.500000 199.830000 1183.980000 200.410000 ;
      RECT 1169.500000 199.590000 1186.000000 199.830000 ;
      RECT 1169.500000 198.410000 1170.500000 199.590000 ;
      RECT 0.000000 198.410000 1156.500000 199.835000 ;
      RECT 0.000000 197.590000 1170.500000 198.410000 ;
      RECT 1183.500000 196.410000 1186.000000 199.590000 ;
      RECT 1169.500000 196.410000 1170.500000 197.590000 ;
      RECT 1169.500000 195.590000 1186.000000 196.410000 ;
      RECT 1169.500000 194.410000 1170.500000 195.590000 ;
      RECT 0.000000 194.410000 1156.500000 197.590000 ;
      RECT 0.000000 193.590000 1170.500000 194.410000 ;
      RECT 1183.500000 192.410000 1186.000000 195.590000 ;
      RECT 1169.500000 192.410000 1170.500000 193.590000 ;
      RECT 1169.500000 191.590000 1186.000000 192.410000 ;
      RECT 1169.500000 190.410000 1170.500000 191.590000 ;
      RECT 0.000000 190.410000 1156.500000 193.590000 ;
      RECT 0.000000 189.590000 1170.500000 190.410000 ;
      RECT 1183.500000 188.410000 1186.000000 191.590000 ;
      RECT 1169.500000 188.410000 1170.500000 189.590000 ;
      RECT 1169.500000 187.590000 1186.000000 188.410000 ;
      RECT 1169.500000 186.410000 1170.500000 187.590000 ;
      RECT 0.000000 186.410000 1156.500000 189.590000 ;
      RECT 0.000000 185.590000 1170.500000 186.410000 ;
      RECT 1183.500000 184.410000 1186.000000 187.590000 ;
      RECT 1169.500000 184.410000 1170.500000 185.590000 ;
      RECT 1169.500000 183.590000 1186.000000 184.410000 ;
      RECT 1169.500000 182.410000 1170.500000 183.590000 ;
      RECT 0.000000 182.410000 1156.500000 185.590000 ;
      RECT 0.000000 181.590000 1170.500000 182.410000 ;
      RECT 1183.500000 180.410000 1186.000000 183.590000 ;
      RECT 1169.500000 180.410000 1170.500000 181.590000 ;
      RECT 1169.500000 179.590000 1186.000000 180.410000 ;
      RECT 1169.500000 178.410000 1170.500000 179.590000 ;
      RECT 0.000000 178.410000 1156.500000 181.590000 ;
      RECT 0.000000 177.590000 1170.500000 178.410000 ;
      RECT 1183.500000 176.410000 1186.000000 179.590000 ;
      RECT 1169.500000 176.410000 1170.500000 177.590000 ;
      RECT 1169.500000 175.590000 1186.000000 176.410000 ;
      RECT 1169.500000 174.410000 1170.500000 175.590000 ;
      RECT 0.000000 174.410000 1156.500000 177.590000 ;
      RECT 0.000000 173.590000 1170.500000 174.410000 ;
      RECT 1183.500000 172.410000 1186.000000 175.590000 ;
      RECT 1169.500000 172.410000 1170.500000 173.590000 ;
      RECT 1169.500000 171.590000 1186.000000 172.410000 ;
      RECT 1169.500000 170.410000 1170.500000 171.590000 ;
      RECT 0.000000 170.410000 1156.500000 173.590000 ;
      RECT 0.000000 169.590000 1170.500000 170.410000 ;
      RECT 1183.500000 168.410000 1186.000000 171.590000 ;
      RECT 1169.500000 168.410000 1170.500000 169.590000 ;
      RECT 1169.500000 167.590000 1186.000000 168.410000 ;
      RECT 1169.500000 166.410000 1170.500000 167.590000 ;
      RECT 0.000000 166.410000 1156.500000 169.590000 ;
      RECT 0.000000 165.590000 1170.500000 166.410000 ;
      RECT 1183.500000 164.410000 1186.000000 167.590000 ;
      RECT 1169.500000 164.410000 1170.500000 165.590000 ;
      RECT 1169.500000 163.590000 1186.000000 164.410000 ;
      RECT 1169.500000 162.410000 1170.500000 163.590000 ;
      RECT 0.000000 162.410000 1156.500000 165.590000 ;
      RECT 0.000000 161.590000 1170.500000 162.410000 ;
      RECT 1183.500000 160.410000 1186.000000 163.590000 ;
      RECT 1169.500000 160.410000 1170.500000 161.590000 ;
      RECT 1169.500000 159.590000 1186.000000 160.410000 ;
      RECT 1169.500000 158.410000 1170.500000 159.590000 ;
      RECT 0.000000 158.410000 1156.500000 161.590000 ;
      RECT 0.000000 157.590000 1170.500000 158.410000 ;
      RECT 1183.500000 156.410000 1186.000000 159.590000 ;
      RECT 1169.500000 156.410000 1170.500000 157.590000 ;
      RECT 1169.500000 155.590000 1186.000000 156.410000 ;
      RECT 1169.500000 154.410000 1170.500000 155.590000 ;
      RECT 0.000000 154.410000 1156.500000 157.590000 ;
      RECT 0.000000 153.590000 1170.500000 154.410000 ;
      RECT 1183.500000 152.410000 1186.000000 155.590000 ;
      RECT 1169.500000 152.410000 1170.500000 153.590000 ;
      RECT 1169.500000 151.590000 1186.000000 152.410000 ;
      RECT 1169.500000 150.410000 1170.500000 151.590000 ;
      RECT 0.000000 150.410000 1156.500000 153.590000 ;
      RECT 0.000000 149.590000 1170.500000 150.410000 ;
      RECT 1183.500000 148.410000 1186.000000 151.590000 ;
      RECT 1169.500000 148.410000 1170.500000 149.590000 ;
      RECT 1169.500000 147.590000 1186.000000 148.410000 ;
      RECT 1169.500000 146.410000 1170.500000 147.590000 ;
      RECT 0.000000 146.410000 1156.500000 149.590000 ;
      RECT 0.000000 145.590000 1170.500000 146.410000 ;
      RECT 1183.500000 144.410000 1186.000000 147.590000 ;
      RECT 1169.500000 144.410000 1170.500000 145.590000 ;
      RECT 1169.500000 143.590000 1186.000000 144.410000 ;
      RECT 1169.500000 142.410000 1170.500000 143.590000 ;
      RECT 0.000000 142.410000 1156.500000 145.590000 ;
      RECT 0.000000 141.590000 1170.500000 142.410000 ;
      RECT 1183.500000 140.410000 1186.000000 143.590000 ;
      RECT 1169.500000 140.410000 1170.500000 141.590000 ;
      RECT 1169.500000 139.590000 1186.000000 140.410000 ;
      RECT 1169.500000 138.410000 1170.500000 139.590000 ;
      RECT 0.000000 138.410000 1156.500000 141.590000 ;
      RECT 0.000000 137.590000 1170.500000 138.410000 ;
      RECT 1183.500000 136.410000 1186.000000 139.590000 ;
      RECT 1169.500000 136.410000 1170.500000 137.590000 ;
      RECT 1169.500000 135.590000 1186.000000 136.410000 ;
      RECT 0.000000 135.590000 1156.500000 137.590000 ;
      RECT 0.000000 135.170000 1149.500000 135.590000 ;
      RECT 1183.500000 135.165000 1186.000000 135.590000 ;
      RECT 1169.500000 134.410000 1170.500000 135.590000 ;
      RECT 1157.500000 133.590000 1170.500000 134.410000 ;
      RECT 1183.500000 132.410000 1183.980000 135.165000 ;
      RECT 1169.500000 132.410000 1170.500000 133.590000 ;
      RECT 2.020000 132.410000 1149.500000 135.170000 ;
      RECT 2.020000 132.070000 1156.500000 132.410000 ;
      RECT 1169.500000 132.065000 1183.980000 132.410000 ;
      RECT 1169.500000 131.590000 1186.000000 132.065000 ;
      RECT 1169.500000 130.410000 1170.500000 131.590000 ;
      RECT 0.000000 130.410000 1156.500000 132.070000 ;
      RECT 0.000000 129.590000 1170.500000 130.410000 ;
      RECT 1183.500000 129.485000 1186.000000 131.590000 ;
      RECT 1183.500000 128.410000 1183.980000 129.485000 ;
      RECT 1169.500000 128.410000 1170.500000 129.590000 ;
      RECT 1169.500000 127.590000 1183.980000 128.410000 ;
      RECT 1169.500000 126.410000 1170.500000 127.590000 ;
      RECT 0.000000 126.410000 1156.500000 129.590000 ;
      RECT 1183.500000 126.385000 1183.980000 127.590000 ;
      RECT 0.000000 125.590000 1170.500000 126.410000 ;
      RECT 1183.500000 125.525000 1186.000000 126.385000 ;
      RECT 0.000000 124.575000 1156.500000 125.590000 ;
      RECT 1183.500000 124.410000 1183.980000 125.525000 ;
      RECT 1169.500000 124.410000 1170.500000 125.590000 ;
      RECT 1169.500000 123.590000 1183.980000 124.410000 ;
      RECT 1183.500000 122.425000 1183.980000 123.590000 ;
      RECT 1169.500000 122.410000 1170.500000 123.590000 ;
      RECT 2.020000 122.410000 1156.500000 124.575000 ;
      RECT 2.020000 121.590000 1170.500000 122.410000 ;
      RECT 2.020000 121.475000 1156.500000 121.590000 ;
      RECT 0.000000 120.615000 1156.500000 121.475000 ;
      RECT 1183.500000 120.410000 1186.000000 122.425000 ;
      RECT 1169.500000 120.410000 1170.500000 121.590000 ;
      RECT 1169.500000 119.590000 1186.000000 120.410000 ;
      RECT 1169.500000 118.410000 1170.500000 119.590000 ;
      RECT 2.020000 118.410000 1156.500000 120.615000 ;
      RECT 2.020000 117.590000 1170.500000 118.410000 ;
      RECT 2.020000 117.515000 1156.500000 117.590000 ;
      RECT 1183.500000 116.410000 1186.000000 119.590000 ;
      RECT 1169.500000 116.410000 1170.500000 117.590000 ;
      RECT 1169.500000 115.590000 1186.000000 116.410000 ;
      RECT 0.000000 114.935000 1156.500000 117.515000 ;
      RECT 1183.500000 114.930000 1186.000000 115.590000 ;
      RECT 1169.500000 114.410000 1170.500000 115.590000 ;
      RECT 2.020000 114.410000 1156.500000 114.935000 ;
      RECT 2.020000 113.590000 1170.500000 114.410000 ;
      RECT 1183.500000 112.410000 1183.980000 114.930000 ;
      RECT 1169.500000 112.410000 1170.500000 113.590000 ;
      RECT 2.020000 111.835000 1156.500000 113.590000 ;
      RECT 1169.500000 111.830000 1183.980000 112.410000 ;
      RECT 1169.500000 111.590000 1186.000000 111.830000 ;
      RECT 1169.500000 110.410000 1170.500000 111.590000 ;
      RECT 0.000000 110.410000 1156.500000 111.835000 ;
      RECT 0.000000 109.590000 1170.500000 110.410000 ;
      RECT 1183.500000 108.410000 1186.000000 111.590000 ;
      RECT 1169.500000 108.410000 1170.500000 109.590000 ;
      RECT 1169.500000 107.590000 1186.000000 108.410000 ;
      RECT 1169.500000 106.410000 1170.500000 107.590000 ;
      RECT 0.000000 106.410000 1156.500000 109.590000 ;
      RECT 0.000000 105.590000 1170.500000 106.410000 ;
      RECT 1183.500000 104.410000 1186.000000 107.590000 ;
      RECT 1169.500000 104.410000 1170.500000 105.590000 ;
      RECT 1169.500000 103.590000 1186.000000 104.410000 ;
      RECT 1169.500000 102.410000 1170.500000 103.590000 ;
      RECT 0.000000 102.410000 1156.500000 105.590000 ;
      RECT 0.000000 101.590000 1170.500000 102.410000 ;
      RECT 1183.500000 100.410000 1186.000000 103.590000 ;
      RECT 1169.500000 100.410000 1170.500000 101.590000 ;
      RECT 1169.500000 99.590000 1186.000000 100.410000 ;
      RECT 1169.500000 98.410000 1170.500000 99.590000 ;
      RECT 0.000000 98.410000 1156.500000 101.590000 ;
      RECT 0.000000 97.590000 1170.500000 98.410000 ;
      RECT 1183.500000 96.410000 1186.000000 99.590000 ;
      RECT 1169.500000 96.410000 1170.500000 97.590000 ;
      RECT 1169.500000 95.590000 1186.000000 96.410000 ;
      RECT 1169.500000 94.410000 1170.500000 95.590000 ;
      RECT 0.000000 94.410000 1156.500000 97.590000 ;
      RECT 0.000000 93.590000 1170.500000 94.410000 ;
      RECT 1183.500000 92.410000 1186.000000 95.590000 ;
      RECT 1169.500000 92.410000 1170.500000 93.590000 ;
      RECT 1169.500000 91.590000 1186.000000 92.410000 ;
      RECT 1169.500000 90.410000 1170.500000 91.590000 ;
      RECT 0.000000 90.410000 1156.500000 93.590000 ;
      RECT 0.000000 89.590000 1170.500000 90.410000 ;
      RECT 1183.500000 88.410000 1186.000000 91.590000 ;
      RECT 1169.500000 88.410000 1170.500000 89.590000 ;
      RECT 1169.500000 87.590000 1186.000000 88.410000 ;
      RECT 1169.500000 86.410000 1170.500000 87.590000 ;
      RECT 0.000000 86.410000 1156.500000 89.590000 ;
      RECT 0.000000 85.590000 1170.500000 86.410000 ;
      RECT 1183.500000 84.410000 1186.000000 87.590000 ;
      RECT 1169.500000 84.410000 1170.500000 85.590000 ;
      RECT 1169.500000 83.590000 1186.000000 84.410000 ;
      RECT 1169.500000 82.410000 1170.500000 83.590000 ;
      RECT 0.000000 82.410000 1156.500000 85.590000 ;
      RECT 0.000000 81.590000 1170.500000 82.410000 ;
      RECT 1183.500000 80.410000 1186.000000 83.590000 ;
      RECT 1169.500000 80.410000 1170.500000 81.590000 ;
      RECT 1169.500000 79.590000 1186.000000 80.410000 ;
      RECT 1169.500000 78.410000 1170.500000 79.590000 ;
      RECT 0.000000 78.410000 1156.500000 81.590000 ;
      RECT 0.000000 77.590000 1170.500000 78.410000 ;
      RECT 1183.500000 76.410000 1186.000000 79.590000 ;
      RECT 1169.500000 76.410000 1170.500000 77.590000 ;
      RECT 1169.500000 75.590000 1186.000000 76.410000 ;
      RECT 1169.500000 74.410000 1170.500000 75.590000 ;
      RECT 0.000000 74.410000 1156.500000 77.590000 ;
      RECT 0.000000 73.590000 1170.500000 74.410000 ;
      RECT 1183.500000 72.410000 1186.000000 75.590000 ;
      RECT 1169.500000 72.410000 1170.500000 73.590000 ;
      RECT 1169.500000 71.590000 1186.000000 72.410000 ;
      RECT 1169.500000 70.410000 1170.500000 71.590000 ;
      RECT 0.000000 70.410000 1156.500000 73.590000 ;
      RECT 0.000000 69.590000 1170.500000 70.410000 ;
      RECT 1183.500000 68.410000 1186.000000 71.590000 ;
      RECT 1169.500000 68.410000 1170.500000 69.590000 ;
      RECT 1169.500000 67.590000 1186.000000 68.410000 ;
      RECT 1169.500000 66.410000 1170.500000 67.590000 ;
      RECT 0.000000 66.410000 1156.500000 69.590000 ;
      RECT 0.000000 65.590000 1170.500000 66.410000 ;
      RECT 1183.500000 64.410000 1186.000000 67.590000 ;
      RECT 1169.500000 64.410000 1170.500000 65.590000 ;
      RECT 1169.500000 63.590000 1186.000000 64.410000 ;
      RECT 1169.500000 62.410000 1170.500000 63.590000 ;
      RECT 0.000000 62.410000 1156.500000 65.590000 ;
      RECT 0.000000 61.590000 1170.500000 62.410000 ;
      RECT 1183.500000 60.410000 1186.000000 63.590000 ;
      RECT 1169.500000 60.410000 1170.500000 61.590000 ;
      RECT 1169.500000 59.590000 1186.000000 60.410000 ;
      RECT 1169.500000 58.410000 1170.500000 59.590000 ;
      RECT 0.000000 58.410000 1156.500000 61.590000 ;
      RECT 0.000000 57.590000 1170.500000 58.410000 ;
      RECT 1183.500000 56.410000 1186.000000 59.590000 ;
      RECT 1169.500000 56.410000 1170.500000 57.590000 ;
      RECT 1169.500000 55.590000 1186.000000 56.410000 ;
      RECT 1169.500000 54.410000 1170.500000 55.590000 ;
      RECT 0.000000 54.410000 1156.500000 57.590000 ;
      RECT 0.000000 53.590000 1170.500000 54.410000 ;
      RECT 1183.500000 52.410000 1186.000000 55.590000 ;
      RECT 1169.500000 52.410000 1170.500000 53.590000 ;
      RECT 1169.500000 51.590000 1186.000000 52.410000 ;
      RECT 1169.500000 50.410000 1170.500000 51.590000 ;
      RECT 0.000000 50.410000 1156.500000 53.590000 ;
      RECT 0.000000 49.590000 1170.500000 50.410000 ;
      RECT 1183.500000 48.410000 1186.000000 51.590000 ;
      RECT 1169.500000 48.410000 1170.500000 49.590000 ;
      RECT 1169.500000 47.590000 1186.000000 48.410000 ;
      RECT 0.000000 47.170000 1156.500000 49.590000 ;
      RECT 1183.500000 47.165000 1186.000000 47.590000 ;
      RECT 1169.500000 46.410000 1170.500000 47.590000 ;
      RECT 2.020000 46.410000 1156.500000 47.170000 ;
      RECT 2.020000 45.590000 1170.500000 46.410000 ;
      RECT 1183.500000 44.410000 1183.980000 47.165000 ;
      RECT 1169.500000 44.410000 1170.500000 45.590000 ;
      RECT 2.020000 44.070000 1156.500000 45.590000 ;
      RECT 1169.500000 44.065000 1183.980000 44.410000 ;
      RECT 1169.500000 43.590000 1186.000000 44.065000 ;
      RECT 1169.500000 42.410000 1170.500000 43.590000 ;
      RECT 0.000000 42.410000 1156.500000 44.070000 ;
      RECT 0.000000 41.590000 1170.500000 42.410000 ;
      RECT 1183.500000 41.485000 1186.000000 43.590000 ;
      RECT 1183.500000 40.410000 1183.980000 41.485000 ;
      RECT 1169.500000 40.410000 1170.500000 41.590000 ;
      RECT 1169.500000 39.590000 1183.980000 40.410000 ;
      RECT 1169.500000 38.410000 1170.500000 39.590000 ;
      RECT 0.000000 38.410000 1156.500000 41.590000 ;
      RECT 1183.500000 38.385000 1183.980000 39.590000 ;
      RECT 0.000000 37.590000 1170.500000 38.410000 ;
      RECT 1183.500000 37.525000 1186.000000 38.385000 ;
      RECT 0.000000 36.575000 1156.500000 37.590000 ;
      RECT 1183.500000 36.410000 1183.980000 37.525000 ;
      RECT 1169.500000 36.410000 1170.500000 37.590000 ;
      RECT 1169.500000 35.590000 1183.980000 36.410000 ;
      RECT 1183.500000 34.425000 1183.980000 35.590000 ;
      RECT 1169.500000 34.410000 1170.500000 35.590000 ;
      RECT 2.020000 34.410000 1156.500000 36.575000 ;
      RECT 2.020000 33.590000 1170.500000 34.410000 ;
      RECT 2.020000 33.475000 1156.500000 33.590000 ;
      RECT 0.000000 32.615000 1156.500000 33.475000 ;
      RECT 1183.500000 32.410000 1186.000000 34.425000 ;
      RECT 1169.500000 32.410000 1170.500000 33.590000 ;
      RECT 1169.500000 31.590000 1186.000000 32.410000 ;
      RECT 1169.500000 30.410000 1170.500000 31.590000 ;
      RECT 2.020000 30.410000 1156.500000 32.615000 ;
      RECT 2.020000 29.590000 1170.500000 30.410000 ;
      RECT 2.020000 29.515000 1156.500000 29.590000 ;
      RECT 1183.500000 28.410000 1186.000000 31.590000 ;
      RECT 1169.500000 28.410000 1170.500000 29.590000 ;
      RECT 1169.500000 27.590000 1186.000000 28.410000 ;
      RECT 0.000000 26.935000 1156.500000 29.515000 ;
      RECT 1183.500000 26.930000 1186.000000 27.590000 ;
      RECT 1169.500000 26.410000 1170.500000 27.590000 ;
      RECT 2.020000 26.410000 1156.500000 26.935000 ;
      RECT 2.020000 25.590000 1170.500000 26.410000 ;
      RECT 1183.500000 24.410000 1183.980000 26.930000 ;
      RECT 1169.500000 24.410000 1170.500000 25.590000 ;
      RECT 2.020000 23.835000 1156.500000 25.590000 ;
      RECT 1169.500000 23.830000 1183.980000 24.410000 ;
      RECT 1169.500000 23.590000 1186.000000 23.830000 ;
      RECT 1169.500000 22.410000 1170.500000 23.590000 ;
      RECT 0.000000 22.410000 1156.500000 23.835000 ;
      RECT 0.000000 21.590000 1170.500000 22.410000 ;
      RECT 1183.500000 20.410000 1186.000000 23.590000 ;
      RECT 1169.500000 20.410000 1170.500000 21.590000 ;
      RECT 1169.500000 19.590000 1186.000000 20.410000 ;
      RECT 1169.500000 18.410000 1170.500000 19.590000 ;
      RECT 0.000000 18.410000 1156.500000 21.590000 ;
      RECT 0.000000 17.590000 1170.500000 18.410000 ;
      RECT 1183.500000 16.410000 1186.000000 19.590000 ;
      RECT 1166.500000 16.410000 1170.500000 17.590000 ;
      RECT 1166.500000 15.590000 1186.000000 16.410000 ;
      RECT 1166.500000 14.410000 1170.500000 15.590000 ;
      RECT 0.000000 14.410000 1158.500000 17.590000 ;
      RECT 0.000000 13.590000 1170.500000 14.410000 ;
      RECT 1183.500000 12.410000 1186.000000 15.590000 ;
      RECT 1166.500000 12.410000 1170.500000 13.590000 ;
      RECT 1166.500000 11.590000 1186.000000 12.410000 ;
      RECT 1166.500000 10.410000 1170.500000 11.590000 ;
      RECT 0.000000 10.410000 1158.500000 13.590000 ;
      RECT 0.000000 9.590000 1170.500000 10.410000 ;
      RECT 1183.500000 8.410000 1186.000000 11.590000 ;
      RECT 1166.500000 8.410000 1170.500000 9.590000 ;
      RECT 1166.500000 7.590000 1186.000000 8.410000 ;
      RECT 1116.500000 7.590000 1158.500000 9.590000 ;
      RECT 1066.500000 7.590000 1108.500000 9.590000 ;
      RECT 1016.500000 7.590000 1058.500000 9.590000 ;
      RECT 966.500000 7.590000 1008.500000 9.590000 ;
      RECT 916.500000 7.590000 958.500000 9.590000 ;
      RECT 866.500000 7.590000 908.500000 9.590000 ;
      RECT 816.500000 7.590000 858.500000 9.590000 ;
      RECT 766.500000 7.590000 808.500000 9.590000 ;
      RECT 716.500000 7.590000 758.500000 9.590000 ;
      RECT 666.500000 7.590000 708.500000 9.590000 ;
      RECT 616.500000 7.590000 658.500000 9.590000 ;
      RECT 566.500000 7.590000 608.500000 9.590000 ;
      RECT 516.500000 7.590000 558.500000 9.590000 ;
      RECT 466.500000 7.590000 508.500000 9.590000 ;
      RECT 416.500000 7.590000 458.500000 9.590000 ;
      RECT 366.500000 7.590000 408.500000 9.590000 ;
      RECT 316.500000 7.590000 358.500000 9.590000 ;
      RECT 266.500000 7.590000 308.500000 9.590000 ;
      RECT 216.500000 7.590000 258.500000 9.590000 ;
      RECT 166.500000 7.590000 208.500000 9.590000 ;
      RECT 116.500000 7.590000 158.500000 9.590000 ;
      RECT 66.500000 7.590000 108.500000 9.590000 ;
      RECT 0.000000 7.590000 58.500000 9.590000 ;
      RECT 1166.500000 6.410000 1170.500000 7.590000 ;
      RECT 1157.500000 6.410000 1158.500000 7.590000 ;
      RECT 1116.500000 6.410000 1149.500000 7.590000 ;
      RECT 1107.500000 6.410000 1108.500000 7.590000 ;
      RECT 1066.500000 6.410000 1099.500000 7.590000 ;
      RECT 1057.500000 6.410000 1058.500000 7.590000 ;
      RECT 1016.500000 6.410000 1049.500000 7.590000 ;
      RECT 1007.500000 6.410000 1008.500000 7.590000 ;
      RECT 966.500000 6.410000 999.500000 7.590000 ;
      RECT 957.500000 6.410000 958.500000 7.590000 ;
      RECT 916.500000 6.410000 949.500000 7.590000 ;
      RECT 907.500000 6.410000 908.500000 7.590000 ;
      RECT 866.500000 6.410000 899.500000 7.590000 ;
      RECT 857.500000 6.410000 858.500000 7.590000 ;
      RECT 816.500000 6.410000 849.500000 7.590000 ;
      RECT 807.500000 6.410000 808.500000 7.590000 ;
      RECT 766.500000 6.410000 799.500000 7.590000 ;
      RECT 757.500000 6.410000 758.500000 7.590000 ;
      RECT 716.500000 6.410000 749.500000 7.590000 ;
      RECT 707.500000 6.410000 708.500000 7.590000 ;
      RECT 666.500000 6.410000 699.500000 7.590000 ;
      RECT 657.500000 6.410000 658.500000 7.590000 ;
      RECT 616.500000 6.410000 649.500000 7.590000 ;
      RECT 607.500000 6.410000 608.500000 7.590000 ;
      RECT 566.500000 6.410000 599.500000 7.590000 ;
      RECT 557.500000 6.410000 558.500000 7.590000 ;
      RECT 516.500000 6.410000 549.500000 7.590000 ;
      RECT 507.500000 6.410000 508.500000 7.590000 ;
      RECT 466.500000 6.410000 499.500000 7.590000 ;
      RECT 457.500000 6.410000 458.500000 7.590000 ;
      RECT 416.500000 6.410000 449.500000 7.590000 ;
      RECT 407.500000 6.410000 408.500000 7.590000 ;
      RECT 366.500000 6.410000 399.500000 7.590000 ;
      RECT 357.500000 6.410000 358.500000 7.590000 ;
      RECT 316.500000 6.410000 349.500000 7.590000 ;
      RECT 307.500000 6.410000 308.500000 7.590000 ;
      RECT 266.500000 6.410000 299.500000 7.590000 ;
      RECT 257.500000 6.410000 258.500000 7.590000 ;
      RECT 216.500000 6.410000 249.500000 7.590000 ;
      RECT 207.500000 6.410000 208.500000 7.590000 ;
      RECT 166.500000 6.410000 199.500000 7.590000 ;
      RECT 157.500000 6.410000 158.500000 7.590000 ;
      RECT 116.500000 6.410000 149.500000 7.590000 ;
      RECT 107.500000 6.410000 108.500000 7.590000 ;
      RECT 66.500000 6.410000 99.500000 7.590000 ;
      RECT 57.500000 6.410000 58.500000 7.590000 ;
      RECT 1157.500000 5.590000 1170.500000 6.410000 ;
      RECT 1107.500000 5.590000 1149.500000 6.410000 ;
      RECT 1057.500000 5.590000 1099.500000 6.410000 ;
      RECT 1007.500000 5.590000 1049.500000 6.410000 ;
      RECT 957.500000 5.590000 999.500000 6.410000 ;
      RECT 907.500000 5.590000 949.500000 6.410000 ;
      RECT 857.500000 5.590000 899.500000 6.410000 ;
      RECT 807.500000 5.590000 849.500000 6.410000 ;
      RECT 757.500000 5.590000 799.500000 6.410000 ;
      RECT 707.500000 5.590000 749.500000 6.410000 ;
      RECT 657.500000 5.590000 699.500000 6.410000 ;
      RECT 607.500000 5.590000 649.500000 6.410000 ;
      RECT 557.500000 5.590000 599.500000 6.410000 ;
      RECT 507.500000 5.590000 549.500000 6.410000 ;
      RECT 457.500000 5.590000 499.500000 6.410000 ;
      RECT 407.500000 5.590000 449.500000 6.410000 ;
      RECT 357.500000 5.590000 399.500000 6.410000 ;
      RECT 307.500000 5.590000 349.500000 6.410000 ;
      RECT 257.500000 5.590000 299.500000 6.410000 ;
      RECT 207.500000 5.590000 249.500000 6.410000 ;
      RECT 157.500000 5.590000 199.500000 6.410000 ;
      RECT 107.500000 5.590000 149.500000 6.410000 ;
      RECT 57.500000 5.590000 99.500000 6.410000 ;
      RECT 1183.500000 4.410000 1186.000000 7.590000 ;
      RECT 1166.500000 4.410000 1170.500000 5.590000 ;
      RECT 1157.500000 4.410000 1158.500000 5.590000 ;
      RECT 1116.500000 4.410000 1149.500000 5.590000 ;
      RECT 1107.500000 4.410000 1108.500000 5.590000 ;
      RECT 1066.500000 4.410000 1099.500000 5.590000 ;
      RECT 1057.500000 4.410000 1058.500000 5.590000 ;
      RECT 1016.500000 4.410000 1049.500000 5.590000 ;
      RECT 1007.500000 4.410000 1008.500000 5.590000 ;
      RECT 966.500000 4.410000 999.500000 5.590000 ;
      RECT 957.500000 4.410000 958.500000 5.590000 ;
      RECT 916.500000 4.410000 949.500000 5.590000 ;
      RECT 907.500000 4.410000 908.500000 5.590000 ;
      RECT 866.500000 4.410000 899.500000 5.590000 ;
      RECT 857.500000 4.410000 858.500000 5.590000 ;
      RECT 816.500000 4.410000 849.500000 5.590000 ;
      RECT 807.500000 4.410000 808.500000 5.590000 ;
      RECT 766.500000 4.410000 799.500000 5.590000 ;
      RECT 757.500000 4.410000 758.500000 5.590000 ;
      RECT 716.500000 4.410000 749.500000 5.590000 ;
      RECT 707.500000 4.410000 708.500000 5.590000 ;
      RECT 666.500000 4.410000 699.500000 5.590000 ;
      RECT 657.500000 4.410000 658.500000 5.590000 ;
      RECT 616.500000 4.410000 649.500000 5.590000 ;
      RECT 607.500000 4.410000 608.500000 5.590000 ;
      RECT 566.500000 4.410000 599.500000 5.590000 ;
      RECT 557.500000 4.410000 558.500000 5.590000 ;
      RECT 516.500000 4.410000 549.500000 5.590000 ;
      RECT 507.500000 4.410000 508.500000 5.590000 ;
      RECT 466.500000 4.410000 499.500000 5.590000 ;
      RECT 457.500000 4.410000 458.500000 5.590000 ;
      RECT 416.500000 4.410000 449.500000 5.590000 ;
      RECT 407.500000 4.410000 408.500000 5.590000 ;
      RECT 366.500000 4.410000 399.500000 5.590000 ;
      RECT 357.500000 4.410000 358.500000 5.590000 ;
      RECT 316.500000 4.410000 349.500000 5.590000 ;
      RECT 307.500000 4.410000 308.500000 5.590000 ;
      RECT 266.500000 4.410000 299.500000 5.590000 ;
      RECT 257.500000 4.410000 258.500000 5.590000 ;
      RECT 216.500000 4.410000 249.500000 5.590000 ;
      RECT 207.500000 4.410000 208.500000 5.590000 ;
      RECT 166.500000 4.410000 199.500000 5.590000 ;
      RECT 157.500000 4.410000 158.500000 5.590000 ;
      RECT 116.500000 4.410000 149.500000 5.590000 ;
      RECT 107.500000 4.410000 108.500000 5.590000 ;
      RECT 66.500000 4.410000 99.500000 5.590000 ;
      RECT 57.500000 4.410000 58.500000 5.590000 ;
      RECT 15.500000 4.410000 49.500000 7.590000 ;
      RECT 0.000000 4.410000 2.500000 7.590000 ;
      RECT 1116.500000 3.590000 1158.500000 4.410000 ;
      RECT 1066.500000 3.590000 1108.500000 4.410000 ;
      RECT 1016.500000 3.590000 1058.500000 4.410000 ;
      RECT 966.500000 3.590000 1008.500000 4.410000 ;
      RECT 916.500000 3.590000 958.500000 4.410000 ;
      RECT 866.500000 3.590000 908.500000 4.410000 ;
      RECT 816.500000 3.590000 858.500000 4.410000 ;
      RECT 766.500000 3.590000 808.500000 4.410000 ;
      RECT 716.500000 3.590000 758.500000 4.410000 ;
      RECT 666.500000 3.590000 708.500000 4.410000 ;
      RECT 616.500000 3.590000 658.500000 4.410000 ;
      RECT 566.500000 3.590000 608.500000 4.410000 ;
      RECT 516.500000 3.590000 558.500000 4.410000 ;
      RECT 466.500000 3.590000 508.500000 4.410000 ;
      RECT 416.500000 3.590000 458.500000 4.410000 ;
      RECT 366.500000 3.590000 408.500000 4.410000 ;
      RECT 316.500000 3.590000 358.500000 4.410000 ;
      RECT 266.500000 3.590000 308.500000 4.410000 ;
      RECT 216.500000 3.590000 258.500000 4.410000 ;
      RECT 166.500000 3.590000 208.500000 4.410000 ;
      RECT 116.500000 3.590000 158.500000 4.410000 ;
      RECT 66.500000 3.590000 108.500000 4.410000 ;
      RECT 0.000000 3.590000 58.500000 4.410000 ;
      RECT 1166.500000 2.410000 1186.000000 4.410000 ;
      RECT 1157.500000 2.410000 1158.500000 3.590000 ;
      RECT 1116.500000 2.410000 1149.500000 3.590000 ;
      RECT 1107.500000 2.410000 1108.500000 3.590000 ;
      RECT 1066.500000 2.410000 1099.500000 3.590000 ;
      RECT 1057.500000 2.410000 1058.500000 3.590000 ;
      RECT 1016.500000 2.410000 1049.500000 3.590000 ;
      RECT 1007.500000 2.410000 1008.500000 3.590000 ;
      RECT 966.500000 2.410000 999.500000 3.590000 ;
      RECT 957.500000 2.410000 958.500000 3.590000 ;
      RECT 916.500000 2.410000 949.500000 3.590000 ;
      RECT 907.500000 2.410000 908.500000 3.590000 ;
      RECT 866.500000 2.410000 899.500000 3.590000 ;
      RECT 857.500000 2.410000 858.500000 3.590000 ;
      RECT 816.500000 2.410000 849.500000 3.590000 ;
      RECT 807.500000 2.410000 808.500000 3.590000 ;
      RECT 766.500000 2.410000 799.500000 3.590000 ;
      RECT 757.500000 2.410000 758.500000 3.590000 ;
      RECT 716.500000 2.410000 749.500000 3.590000 ;
      RECT 707.500000 2.410000 708.500000 3.590000 ;
      RECT 666.500000 2.410000 699.500000 3.590000 ;
      RECT 657.500000 2.410000 658.500000 3.590000 ;
      RECT 616.500000 2.410000 649.500000 3.590000 ;
      RECT 607.500000 2.410000 608.500000 3.590000 ;
      RECT 566.500000 2.410000 599.500000 3.590000 ;
      RECT 557.500000 2.410000 558.500000 3.590000 ;
      RECT 516.500000 2.410000 549.500000 3.590000 ;
      RECT 507.500000 2.410000 508.500000 3.590000 ;
      RECT 466.500000 2.410000 499.500000 3.590000 ;
      RECT 457.500000 2.410000 458.500000 3.590000 ;
      RECT 416.500000 2.410000 449.500000 3.590000 ;
      RECT 407.500000 2.410000 408.500000 3.590000 ;
      RECT 366.500000 2.410000 399.500000 3.590000 ;
      RECT 357.500000 2.410000 358.500000 3.590000 ;
      RECT 316.500000 2.410000 349.500000 3.590000 ;
      RECT 307.500000 2.410000 308.500000 3.590000 ;
      RECT 266.500000 2.410000 299.500000 3.590000 ;
      RECT 257.500000 2.410000 258.500000 3.590000 ;
      RECT 216.500000 2.410000 249.500000 3.590000 ;
      RECT 207.500000 2.410000 208.500000 3.590000 ;
      RECT 166.500000 2.410000 199.500000 3.590000 ;
      RECT 157.500000 2.410000 158.500000 3.590000 ;
      RECT 116.500000 2.410000 149.500000 3.590000 ;
      RECT 107.500000 2.410000 108.500000 3.590000 ;
      RECT 66.500000 2.410000 99.500000 3.590000 ;
      RECT 57.500000 2.410000 58.500000 3.590000 ;
      RECT 857.500000 2.020000 899.500000 2.410000 ;
      RECT 807.500000 2.020000 849.500000 2.410000 ;
      RECT 757.500000 2.020000 799.500000 2.410000 ;
      RECT 707.500000 2.020000 749.500000 2.410000 ;
      RECT 607.500000 2.020000 649.500000 2.410000 ;
      RECT 557.500000 2.020000 599.500000 2.410000 ;
      RECT 507.500000 2.020000 549.500000 2.410000 ;
      RECT 457.500000 2.020000 499.500000 2.410000 ;
      RECT 357.500000 2.020000 399.500000 2.410000 ;
      RECT 257.500000 2.020000 299.500000 2.410000 ;
      RECT 107.500000 2.020000 149.500000 2.410000 ;
      RECT 1157.500000 0.410000 1186.000000 2.410000 ;
      RECT 1107.500000 0.410000 1149.500000 2.410000 ;
      RECT 1057.500000 0.410000 1099.500000 2.410000 ;
      RECT 1007.500000 0.410000 1049.500000 2.410000 ;
      RECT 957.500000 0.410000 999.500000 2.410000 ;
      RECT 907.500000 0.410000 949.500000 2.410000 ;
      RECT 899.485000 0.410000 899.500000 2.020000 ;
      RECT 857.500000 0.410000 881.830000 2.020000 ;
      RECT 819.365000 0.410000 849.500000 2.020000 ;
      RECT 799.130000 0.410000 799.500000 2.020000 ;
      RECT 757.500000 0.410000 796.030000 2.020000 ;
      RECT 733.565000 0.410000 749.500000 2.020000 ;
      RECT 707.500000 0.410000 710.230000 2.020000 ;
      RECT 657.500000 0.410000 699.500000 2.410000 ;
      RECT 647.765000 0.410000 649.500000 2.020000 ;
      RECT 607.500000 0.410000 624.430000 2.020000 ;
      RECT 561.965000 0.410000 599.500000 2.020000 ;
      RECT 557.500000 0.410000 558.865000 2.020000 ;
      RECT 507.500000 0.410000 538.630000 2.020000 ;
      RECT 476.165000 0.410000 499.500000 2.020000 ;
      RECT 457.500000 0.410000 463.425000 2.020000 ;
      RECT 407.500000 0.410000 449.500000 2.410000 ;
      RECT 390.365000 0.410000 399.500000 2.020000 ;
      RECT 357.500000 0.410000 367.030000 2.020000 ;
      RECT 307.500000 0.410000 349.500000 2.410000 ;
      RECT 298.885000 0.410000 299.500000 2.020000 ;
      RECT 257.500000 0.410000 281.230000 2.020000 ;
      RECT 207.500000 0.410000 249.500000 2.410000 ;
      RECT 157.500000 0.410000 199.500000 2.410000 ;
      RECT 132.965000 0.410000 149.500000 2.020000 ;
      RECT 107.500000 0.410000 109.630000 2.020000 ;
      RECT 57.500000 0.410000 99.500000 2.410000 ;
      RECT 0.000000 0.410000 49.500000 3.590000 ;
      RECT 905.165000 0.000000 1186.000000 0.410000 ;
      RECT 899.485000 0.000000 902.065000 0.410000 ;
      RECT 895.525000 0.000000 896.385000 2.020000 ;
      RECT 884.930000 0.000000 892.425000 2.020000 ;
      RECT 819.365000 0.000000 881.830000 0.410000 ;
      RECT 813.685000 0.000000 816.265000 2.020000 ;
      RECT 809.725000 0.000000 810.585000 2.020000 ;
      RECT 799.130000 0.000000 806.625000 0.410000 ;
      RECT 733.565000 0.000000 796.030000 0.410000 ;
      RECT 727.885000 0.000000 730.465000 2.020000 ;
      RECT 723.925000 0.000000 724.785000 2.020000 ;
      RECT 713.330000 0.000000 720.825000 2.020000 ;
      RECT 647.765000 0.000000 710.230000 0.410000 ;
      RECT 642.085000 0.000000 644.665000 2.020000 ;
      RECT 638.125000 0.000000 638.985000 2.020000 ;
      RECT 627.530000 0.000000 635.025000 2.020000 ;
      RECT 561.965000 0.000000 624.430000 0.410000 ;
      RECT 556.285000 0.000000 558.865000 0.410000 ;
      RECT 552.325000 0.000000 553.185000 0.410000 ;
      RECT 541.730000 0.000000 549.225000 2.020000 ;
      RECT 476.165000 0.000000 538.630000 0.410000 ;
      RECT 470.485000 0.000000 473.065000 2.020000 ;
      RECT 466.525000 0.000000 467.385000 2.020000 ;
      RECT 455.930000 0.000000 463.425000 0.410000 ;
      RECT 390.365000 0.000000 452.830000 0.410000 ;
      RECT 384.685000 0.000000 387.265000 2.020000 ;
      RECT 380.725000 0.000000 381.585000 2.020000 ;
      RECT 370.130000 0.000000 377.625000 2.020000 ;
      RECT 304.565000 0.000000 367.030000 0.410000 ;
      RECT 298.885000 0.000000 301.465000 0.410000 ;
      RECT 294.925000 0.000000 295.785000 2.020000 ;
      RECT 284.330000 0.000000 291.825000 2.020000 ;
      RECT 132.965000 0.000000 281.230000 0.410000 ;
      RECT 127.285000 0.000000 129.865000 2.020000 ;
      RECT 123.325000 0.000000 124.185000 2.020000 ;
      RECT 112.730000 0.000000 120.225000 2.020000 ;
      RECT 0.000000 0.000000 109.630000 0.410000 ;
    LAYER M3 ;
      RECT 1139.000000 685.590000 1186.000000 686.000000 ;
      RECT 0.000000 685.590000 670.000000 686.000000 ;
      RECT 1139.000000 683.590000 1158.500000 685.590000 ;
      RECT 616.500000 683.590000 658.500000 685.590000 ;
      RECT 566.500000 683.590000 608.500000 685.590000 ;
      RECT 516.500000 683.590000 558.500000 685.590000 ;
      RECT 466.500000 683.590000 508.500000 685.590000 ;
      RECT 416.500000 683.590000 458.500000 685.590000 ;
      RECT 366.500000 683.590000 408.500000 685.590000 ;
      RECT 316.500000 683.590000 358.500000 685.590000 ;
      RECT 0.000000 683.590000 308.500000 685.590000 ;
      RECT 1166.500000 682.410000 1186.000000 685.590000 ;
      RECT 1157.500000 682.410000 1158.500000 683.590000 ;
      RECT 666.500000 682.410000 670.000000 685.590000 ;
      RECT 657.500000 682.410000 658.500000 683.590000 ;
      RECT 616.500000 682.410000 649.500000 683.590000 ;
      RECT 607.500000 682.410000 608.500000 683.590000 ;
      RECT 566.500000 682.410000 599.500000 683.590000 ;
      RECT 557.500000 682.410000 558.500000 683.590000 ;
      RECT 516.500000 682.410000 549.500000 683.590000 ;
      RECT 507.500000 682.410000 508.500000 683.590000 ;
      RECT 466.500000 682.410000 499.500000 683.590000 ;
      RECT 457.500000 682.410000 458.500000 683.590000 ;
      RECT 416.500000 682.410000 449.500000 683.590000 ;
      RECT 407.500000 682.410000 408.500000 683.590000 ;
      RECT 366.500000 682.410000 373.500000 683.590000 ;
      RECT 357.500000 682.410000 358.500000 683.590000 ;
      RECT 316.500000 682.410000 349.500000 683.590000 ;
      RECT 307.500000 682.410000 308.500000 683.590000 ;
      RECT 1157.500000 681.590000 1186.000000 682.410000 ;
      RECT 657.500000 681.590000 670.000000 682.410000 ;
      RECT 607.500000 681.590000 649.500000 682.410000 ;
      RECT 557.500000 681.590000 599.500000 682.410000 ;
      RECT 507.500000 681.590000 549.500000 682.410000 ;
      RECT 457.500000 681.590000 499.500000 682.410000 ;
      RECT 407.500000 681.590000 449.500000 682.410000 ;
      RECT 357.500000 681.590000 373.500000 682.410000 ;
      RECT 307.500000 681.590000 349.500000 682.410000 ;
      RECT 1157.500000 680.410000 1158.500000 681.590000 ;
      RECT 1139.000000 680.410000 1149.500000 683.590000 ;
      RECT 657.500000 680.410000 658.500000 681.590000 ;
      RECT 616.500000 680.410000 649.500000 681.590000 ;
      RECT 607.500000 680.410000 608.500000 681.590000 ;
      RECT 566.500000 680.410000 599.500000 681.590000 ;
      RECT 557.500000 680.410000 558.500000 681.590000 ;
      RECT 516.500000 680.410000 549.500000 681.590000 ;
      RECT 507.500000 680.410000 508.500000 681.590000 ;
      RECT 466.500000 680.410000 499.500000 681.590000 ;
      RECT 457.500000 680.410000 458.500000 681.590000 ;
      RECT 416.500000 680.410000 449.500000 681.590000 ;
      RECT 407.500000 680.410000 408.500000 681.590000 ;
      RECT 386.500000 680.410000 399.500000 683.590000 ;
      RECT 366.500000 680.410000 373.500000 681.590000 ;
      RECT 357.500000 680.410000 358.500000 681.590000 ;
      RECT 316.500000 680.410000 349.500000 681.590000 ;
      RECT 307.500000 680.410000 308.500000 681.590000 ;
      RECT 0.000000 680.410000 299.500000 683.590000 ;
      RECT 1139.000000 679.590000 1158.500000 680.410000 ;
      RECT 616.500000 679.590000 658.500000 680.410000 ;
      RECT 566.500000 679.590000 608.500000 680.410000 ;
      RECT 516.500000 679.590000 558.500000 680.410000 ;
      RECT 466.500000 679.590000 508.500000 680.410000 ;
      RECT 416.500000 679.590000 458.500000 680.410000 ;
      RECT 366.500000 679.590000 408.500000 680.410000 ;
      RECT 316.500000 679.590000 358.500000 680.410000 ;
      RECT 0.000000 679.590000 308.500000 680.410000 ;
      RECT 1166.500000 678.410000 1186.000000 681.590000 ;
      RECT 1157.500000 678.410000 1158.500000 679.590000 ;
      RECT 666.500000 678.410000 670.000000 681.590000 ;
      RECT 657.500000 678.410000 658.500000 679.590000 ;
      RECT 616.500000 678.410000 649.500000 679.590000 ;
      RECT 607.500000 678.410000 608.500000 679.590000 ;
      RECT 566.500000 678.410000 599.500000 679.590000 ;
      RECT 557.500000 678.410000 558.500000 679.590000 ;
      RECT 516.500000 678.410000 549.500000 679.590000 ;
      RECT 507.500000 678.410000 508.500000 679.590000 ;
      RECT 466.500000 678.410000 499.500000 679.590000 ;
      RECT 457.500000 678.410000 458.500000 679.590000 ;
      RECT 416.500000 678.410000 449.500000 679.590000 ;
      RECT 407.500000 678.410000 408.500000 679.590000 ;
      RECT 366.500000 678.410000 373.500000 679.590000 ;
      RECT 357.500000 678.410000 358.500000 679.590000 ;
      RECT 316.500000 678.410000 349.500000 679.590000 ;
      RECT 307.500000 678.410000 308.500000 679.590000 ;
      RECT 1157.500000 677.590000 1186.000000 678.410000 ;
      RECT 657.500000 677.590000 670.000000 678.410000 ;
      RECT 607.500000 677.590000 649.500000 678.410000 ;
      RECT 557.500000 677.590000 599.500000 678.410000 ;
      RECT 507.500000 677.590000 549.500000 678.410000 ;
      RECT 457.500000 677.590000 499.500000 678.410000 ;
      RECT 407.500000 677.590000 449.500000 678.410000 ;
      RECT 357.500000 677.590000 373.500000 678.410000 ;
      RECT 1157.500000 676.410000 1158.500000 677.590000 ;
      RECT 1139.000000 676.410000 1149.500000 679.590000 ;
      RECT 657.500000 676.410000 658.500000 677.590000 ;
      RECT 616.500000 676.410000 649.500000 677.590000 ;
      RECT 607.500000 676.410000 608.500000 677.590000 ;
      RECT 566.500000 676.410000 599.500000 677.590000 ;
      RECT 557.500000 676.410000 558.500000 677.590000 ;
      RECT 516.500000 676.410000 549.500000 677.590000 ;
      RECT 507.500000 676.410000 508.500000 677.590000 ;
      RECT 466.500000 676.410000 499.500000 677.590000 ;
      RECT 457.500000 676.410000 458.500000 677.590000 ;
      RECT 416.500000 676.410000 449.500000 677.590000 ;
      RECT 407.500000 676.410000 408.500000 677.590000 ;
      RECT 386.500000 676.410000 399.500000 679.590000 ;
      RECT 366.500000 676.410000 373.500000 677.590000 ;
      RECT 357.500000 676.410000 358.500000 677.590000 ;
      RECT 307.500000 676.410000 349.500000 678.410000 ;
      RECT 0.000000 676.410000 299.500000 679.590000 ;
      RECT 1139.000000 675.590000 1158.500000 676.410000 ;
      RECT 616.500000 675.590000 658.500000 676.410000 ;
      RECT 566.500000 675.590000 608.500000 676.410000 ;
      RECT 516.500000 675.590000 558.500000 676.410000 ;
      RECT 466.500000 675.590000 508.500000 676.410000 ;
      RECT 416.500000 675.590000 458.500000 676.410000 ;
      RECT 366.500000 675.590000 408.500000 676.410000 ;
      RECT 0.000000 675.590000 358.500000 676.410000 ;
      RECT 1166.500000 674.410000 1186.000000 677.590000 ;
      RECT 1157.500000 674.410000 1158.500000 675.590000 ;
      RECT 666.500000 674.410000 670.000000 677.590000 ;
      RECT 657.500000 674.410000 658.500000 675.590000 ;
      RECT 616.500000 674.410000 649.500000 675.590000 ;
      RECT 607.500000 674.410000 608.500000 675.590000 ;
      RECT 566.500000 674.410000 599.500000 675.590000 ;
      RECT 557.500000 674.410000 558.500000 675.590000 ;
      RECT 516.500000 674.410000 549.500000 675.590000 ;
      RECT 507.500000 674.410000 508.500000 675.590000 ;
      RECT 466.500000 674.410000 499.500000 675.590000 ;
      RECT 457.500000 674.410000 458.500000 675.590000 ;
      RECT 416.500000 674.410000 449.500000 675.590000 ;
      RECT 407.500000 674.410000 408.500000 675.590000 ;
      RECT 366.500000 674.410000 373.500000 675.590000 ;
      RECT 357.500000 674.410000 358.500000 675.590000 ;
      RECT 1157.500000 673.590000 1186.000000 674.410000 ;
      RECT 657.500000 673.590000 670.000000 674.410000 ;
      RECT 607.500000 673.590000 649.500000 674.410000 ;
      RECT 557.500000 673.590000 599.500000 674.410000 ;
      RECT 507.500000 673.590000 549.500000 674.410000 ;
      RECT 457.500000 673.590000 499.500000 674.410000 ;
      RECT 407.500000 673.590000 449.500000 674.410000 ;
      RECT 357.500000 673.590000 373.500000 674.410000 ;
      RECT 1157.500000 672.410000 1158.500000 673.590000 ;
      RECT 1139.000000 672.410000 1149.500000 675.590000 ;
      RECT 657.500000 672.410000 658.500000 673.590000 ;
      RECT 616.500000 672.410000 649.500000 673.590000 ;
      RECT 607.500000 672.410000 608.500000 673.590000 ;
      RECT 566.500000 672.410000 599.500000 673.590000 ;
      RECT 557.500000 672.410000 558.500000 673.590000 ;
      RECT 516.500000 672.410000 549.500000 673.590000 ;
      RECT 507.500000 672.410000 508.500000 673.590000 ;
      RECT 466.500000 672.410000 499.500000 673.590000 ;
      RECT 457.500000 672.410000 458.500000 673.590000 ;
      RECT 416.500000 672.410000 449.500000 673.590000 ;
      RECT 407.500000 672.410000 408.500000 673.590000 ;
      RECT 386.500000 672.410000 399.500000 675.590000 ;
      RECT 366.500000 672.410000 373.500000 673.590000 ;
      RECT 357.500000 672.410000 358.500000 673.590000 ;
      RECT 0.000000 672.410000 349.500000 675.590000 ;
      RECT 1139.000000 671.590000 1158.500000 672.410000 ;
      RECT 616.500000 671.590000 658.500000 672.410000 ;
      RECT 566.500000 671.590000 608.500000 672.410000 ;
      RECT 516.500000 671.590000 558.500000 672.410000 ;
      RECT 466.500000 671.590000 508.500000 672.410000 ;
      RECT 416.500000 671.590000 458.500000 672.410000 ;
      RECT 366.500000 671.590000 408.500000 672.410000 ;
      RECT 0.000000 671.590000 358.500000 672.410000 ;
      RECT 1166.500000 670.410000 1186.000000 673.590000 ;
      RECT 1157.500000 670.410000 1158.500000 671.590000 ;
      RECT 666.500000 670.410000 670.000000 673.590000 ;
      RECT 657.500000 670.410000 658.500000 671.590000 ;
      RECT 616.500000 670.410000 649.500000 671.590000 ;
      RECT 607.500000 670.410000 608.500000 671.590000 ;
      RECT 566.500000 670.410000 599.500000 671.590000 ;
      RECT 557.500000 670.410000 558.500000 671.590000 ;
      RECT 516.500000 670.410000 549.500000 671.590000 ;
      RECT 507.500000 670.410000 508.500000 671.590000 ;
      RECT 466.500000 670.410000 499.500000 671.590000 ;
      RECT 457.500000 670.410000 458.500000 671.590000 ;
      RECT 416.500000 670.410000 449.500000 671.590000 ;
      RECT 407.500000 670.410000 408.500000 671.590000 ;
      RECT 366.500000 670.410000 373.500000 671.590000 ;
      RECT 357.500000 670.410000 358.500000 671.590000 ;
      RECT 1157.500000 669.590000 1186.000000 670.410000 ;
      RECT 657.500000 669.590000 670.000000 670.410000 ;
      RECT 607.500000 669.590000 649.500000 670.410000 ;
      RECT 557.500000 669.590000 599.500000 670.410000 ;
      RECT 507.500000 669.590000 549.500000 670.410000 ;
      RECT 457.500000 669.590000 499.500000 670.410000 ;
      RECT 407.500000 669.590000 449.500000 670.410000 ;
      RECT 357.500000 669.590000 373.500000 670.410000 ;
      RECT 1157.500000 668.410000 1158.500000 669.590000 ;
      RECT 1139.000000 668.410000 1149.500000 671.590000 ;
      RECT 657.500000 668.410000 658.500000 669.590000 ;
      RECT 616.500000 668.410000 649.500000 669.590000 ;
      RECT 607.500000 668.410000 608.500000 669.590000 ;
      RECT 566.500000 668.410000 599.500000 669.590000 ;
      RECT 557.500000 668.410000 558.500000 669.590000 ;
      RECT 516.500000 668.410000 549.500000 669.590000 ;
      RECT 507.500000 668.410000 508.500000 669.590000 ;
      RECT 466.500000 668.410000 499.500000 669.590000 ;
      RECT 457.500000 668.410000 458.500000 669.590000 ;
      RECT 416.500000 668.410000 449.500000 669.590000 ;
      RECT 407.500000 668.410000 408.500000 669.590000 ;
      RECT 386.500000 668.410000 399.500000 671.590000 ;
      RECT 372.500000 668.410000 373.500000 669.590000 ;
      RECT 357.500000 668.410000 358.500000 669.590000 ;
      RECT 0.000000 668.410000 349.500000 671.590000 ;
      RECT 1139.000000 667.590000 1158.500000 668.410000 ;
      RECT 616.500000 667.590000 658.500000 668.410000 ;
      RECT 566.500000 667.590000 608.500000 668.410000 ;
      RECT 516.500000 667.590000 558.500000 668.410000 ;
      RECT 466.500000 667.590000 508.500000 668.410000 ;
      RECT 416.500000 667.590000 458.500000 668.410000 ;
      RECT 372.500000 667.590000 408.500000 668.410000 ;
      RECT 0.000000 667.590000 358.500000 668.410000 ;
      RECT 1166.500000 666.410000 1186.000000 669.590000 ;
      RECT 1157.500000 666.410000 1158.500000 667.590000 ;
      RECT 666.500000 666.410000 670.000000 669.590000 ;
      RECT 657.500000 666.410000 658.500000 667.590000 ;
      RECT 616.500000 666.410000 649.500000 667.590000 ;
      RECT 607.500000 666.410000 608.500000 667.590000 ;
      RECT 566.500000 666.410000 599.500000 667.590000 ;
      RECT 557.500000 666.410000 558.500000 667.590000 ;
      RECT 516.500000 666.410000 549.500000 667.590000 ;
      RECT 507.500000 666.410000 508.500000 667.590000 ;
      RECT 466.500000 666.410000 499.500000 667.590000 ;
      RECT 457.500000 666.410000 458.500000 667.590000 ;
      RECT 416.500000 666.410000 449.500000 667.590000 ;
      RECT 407.500000 666.410000 408.500000 667.590000 ;
      RECT 372.500000 666.410000 373.500000 667.590000 ;
      RECT 357.500000 666.410000 358.500000 667.590000 ;
      RECT 1157.500000 665.590000 1186.000000 666.410000 ;
      RECT 657.500000 665.590000 670.000000 666.410000 ;
      RECT 607.500000 665.590000 649.500000 666.410000 ;
      RECT 557.500000 665.590000 599.500000 666.410000 ;
      RECT 507.500000 665.590000 549.500000 666.410000 ;
      RECT 457.500000 665.590000 499.500000 666.410000 ;
      RECT 407.500000 665.590000 449.500000 666.410000 ;
      RECT 357.500000 665.590000 373.500000 666.410000 ;
      RECT 1157.500000 664.410000 1158.500000 665.590000 ;
      RECT 1139.000000 664.410000 1149.500000 667.590000 ;
      RECT 657.500000 664.410000 658.500000 665.590000 ;
      RECT 616.500000 664.410000 649.500000 665.590000 ;
      RECT 607.500000 664.410000 608.500000 665.590000 ;
      RECT 566.500000 664.410000 599.500000 665.590000 ;
      RECT 557.500000 664.410000 558.500000 665.590000 ;
      RECT 516.500000 664.410000 549.500000 665.590000 ;
      RECT 507.500000 664.410000 508.500000 665.590000 ;
      RECT 466.500000 664.410000 499.500000 665.590000 ;
      RECT 457.500000 664.410000 458.500000 665.590000 ;
      RECT 416.500000 664.410000 449.500000 665.590000 ;
      RECT 407.500000 664.410000 408.500000 665.590000 ;
      RECT 386.500000 664.410000 399.500000 667.590000 ;
      RECT 372.500000 664.410000 373.500000 665.590000 ;
      RECT 357.500000 664.410000 358.500000 665.590000 ;
      RECT 0.000000 664.410000 349.500000 667.590000 ;
      RECT 1139.000000 663.590000 1158.500000 664.410000 ;
      RECT 616.500000 663.590000 658.500000 664.410000 ;
      RECT 566.500000 663.590000 608.500000 664.410000 ;
      RECT 516.500000 663.590000 558.500000 664.410000 ;
      RECT 466.500000 663.590000 508.500000 664.410000 ;
      RECT 416.500000 663.590000 458.500000 664.410000 ;
      RECT 372.500000 663.590000 408.500000 664.410000 ;
      RECT 0.000000 663.590000 358.500000 664.410000 ;
      RECT 1166.500000 662.410000 1186.000000 665.590000 ;
      RECT 1157.500000 662.410000 1158.500000 663.590000 ;
      RECT 666.500000 662.410000 670.000000 665.590000 ;
      RECT 657.500000 662.410000 658.500000 663.590000 ;
      RECT 616.500000 662.410000 649.500000 663.590000 ;
      RECT 607.500000 662.410000 608.500000 663.590000 ;
      RECT 566.500000 662.410000 599.500000 663.590000 ;
      RECT 557.500000 662.410000 558.500000 663.590000 ;
      RECT 516.500000 662.410000 549.500000 663.590000 ;
      RECT 507.500000 662.410000 508.500000 663.590000 ;
      RECT 466.500000 662.410000 499.500000 663.590000 ;
      RECT 457.500000 662.410000 458.500000 663.590000 ;
      RECT 416.500000 662.410000 449.500000 663.590000 ;
      RECT 407.500000 662.410000 408.500000 663.590000 ;
      RECT 372.500000 662.410000 373.500000 663.590000 ;
      RECT 357.500000 662.410000 358.500000 663.590000 ;
      RECT 1157.500000 661.590000 1186.000000 662.410000 ;
      RECT 657.500000 661.590000 670.000000 662.410000 ;
      RECT 607.500000 661.590000 649.500000 662.410000 ;
      RECT 557.500000 661.590000 599.500000 662.410000 ;
      RECT 507.500000 661.590000 549.500000 662.410000 ;
      RECT 457.500000 661.590000 499.500000 662.410000 ;
      RECT 407.500000 661.590000 449.500000 662.410000 ;
      RECT 357.500000 661.590000 373.500000 662.410000 ;
      RECT 1157.500000 660.410000 1158.500000 661.590000 ;
      RECT 1139.000000 660.410000 1149.500000 663.590000 ;
      RECT 657.500000 660.410000 658.500000 661.590000 ;
      RECT 616.500000 660.410000 649.500000 661.590000 ;
      RECT 607.500000 660.410000 608.500000 661.590000 ;
      RECT 566.500000 660.410000 599.500000 661.590000 ;
      RECT 557.500000 660.410000 558.500000 661.590000 ;
      RECT 516.500000 660.410000 549.500000 661.590000 ;
      RECT 507.500000 660.410000 508.500000 661.590000 ;
      RECT 466.500000 660.410000 499.500000 661.590000 ;
      RECT 457.500000 660.410000 458.500000 661.590000 ;
      RECT 416.500000 660.410000 449.500000 661.590000 ;
      RECT 407.500000 660.410000 408.500000 661.590000 ;
      RECT 386.500000 660.410000 399.500000 663.590000 ;
      RECT 372.500000 660.410000 373.500000 661.590000 ;
      RECT 357.500000 660.410000 358.500000 661.590000 ;
      RECT 0.000000 660.410000 349.500000 663.590000 ;
      RECT 1139.000000 659.590000 1158.500000 660.410000 ;
      RECT 616.500000 659.590000 658.500000 660.410000 ;
      RECT 566.500000 659.590000 608.500000 660.410000 ;
      RECT 516.500000 659.590000 558.500000 660.410000 ;
      RECT 466.500000 659.590000 508.500000 660.410000 ;
      RECT 416.500000 659.590000 458.500000 660.410000 ;
      RECT 372.500000 659.590000 408.500000 660.410000 ;
      RECT 0.000000 659.590000 358.500000 660.410000 ;
      RECT 1166.500000 658.410000 1186.000000 661.590000 ;
      RECT 1157.500000 658.410000 1158.500000 659.590000 ;
      RECT 666.500000 658.410000 670.000000 661.590000 ;
      RECT 657.500000 658.410000 658.500000 659.590000 ;
      RECT 616.500000 658.410000 649.500000 659.590000 ;
      RECT 607.500000 658.410000 608.500000 659.590000 ;
      RECT 566.500000 658.410000 599.500000 659.590000 ;
      RECT 557.500000 658.410000 558.500000 659.590000 ;
      RECT 516.500000 658.410000 549.500000 659.590000 ;
      RECT 507.500000 658.410000 508.500000 659.590000 ;
      RECT 466.500000 658.410000 499.500000 659.590000 ;
      RECT 457.500000 658.410000 458.500000 659.590000 ;
      RECT 416.500000 658.410000 449.500000 659.590000 ;
      RECT 407.500000 658.410000 408.500000 659.590000 ;
      RECT 372.500000 658.410000 373.500000 659.590000 ;
      RECT 357.500000 658.410000 358.500000 659.590000 ;
      RECT 1157.500000 657.590000 1186.000000 658.410000 ;
      RECT 357.500000 657.590000 373.500000 658.410000 ;
      RECT 1157.500000 656.410000 1158.500000 657.590000 ;
      RECT 1139.000000 656.410000 1149.500000 659.590000 ;
      RECT 657.500000 656.410000 670.000000 658.410000 ;
      RECT 607.500000 656.410000 649.500000 658.410000 ;
      RECT 557.500000 656.410000 599.500000 658.410000 ;
      RECT 507.500000 656.410000 549.500000 658.410000 ;
      RECT 457.500000 656.410000 499.500000 658.410000 ;
      RECT 407.500000 656.410000 449.500000 658.410000 ;
      RECT 386.500000 656.410000 399.500000 659.590000 ;
      RECT 372.500000 656.410000 373.500000 657.590000 ;
      RECT 357.500000 656.410000 358.500000 657.590000 ;
      RECT 0.000000 656.410000 349.500000 659.590000 ;
      RECT 372.500000 656.000000 670.000000 656.410000 ;
      RECT 1139.000000 655.590000 1158.500000 656.410000 ;
      RECT 372.500000 655.590000 389.000000 656.000000 ;
      RECT 0.000000 655.590000 358.500000 656.410000 ;
      RECT 1166.500000 654.410000 1186.000000 657.590000 ;
      RECT 1157.500000 654.410000 1158.500000 655.590000 ;
      RECT 372.500000 654.410000 373.500000 655.590000 ;
      RECT 357.500000 654.410000 358.500000 655.590000 ;
      RECT 1157.500000 653.590000 1186.000000 654.410000 ;
      RECT 357.500000 653.590000 373.500000 654.410000 ;
      RECT 1157.500000 652.410000 1158.500000 653.590000 ;
      RECT 1139.000000 652.410000 1149.500000 655.590000 ;
      RECT 386.500000 652.410000 389.000000 655.590000 ;
      RECT 372.500000 652.410000 373.500000 653.590000 ;
      RECT 357.500000 652.410000 358.500000 653.590000 ;
      RECT 0.000000 652.410000 349.500000 655.590000 ;
      RECT 1139.000000 651.590000 1158.500000 652.410000 ;
      RECT 372.500000 651.590000 389.000000 652.410000 ;
      RECT 0.000000 651.590000 358.500000 652.410000 ;
      RECT 1166.500000 650.410000 1186.000000 653.590000 ;
      RECT 1157.500000 650.410000 1158.500000 651.590000 ;
      RECT 372.500000 650.410000 373.500000 651.590000 ;
      RECT 357.500000 650.410000 358.500000 651.590000 ;
      RECT 1157.500000 649.590000 1186.000000 650.410000 ;
      RECT 357.500000 649.590000 373.500000 650.410000 ;
      RECT 1157.500000 648.410000 1158.500000 649.590000 ;
      RECT 1139.000000 648.410000 1149.500000 651.590000 ;
      RECT 386.500000 648.410000 389.000000 651.590000 ;
      RECT 372.500000 648.410000 373.500000 649.590000 ;
      RECT 357.500000 648.410000 358.500000 649.590000 ;
      RECT 0.000000 648.410000 349.500000 651.590000 ;
      RECT 1139.000000 647.590000 1158.500000 648.410000 ;
      RECT 372.500000 647.590000 389.000000 648.410000 ;
      RECT 0.000000 647.590000 358.500000 648.410000 ;
      RECT 1166.500000 646.410000 1186.000000 649.590000 ;
      RECT 1157.500000 646.410000 1158.500000 647.590000 ;
      RECT 372.500000 646.410000 373.500000 647.590000 ;
      RECT 357.500000 646.410000 358.500000 647.590000 ;
      RECT 1157.500000 645.590000 1186.000000 646.410000 ;
      RECT 357.500000 645.590000 373.500000 646.410000 ;
      RECT 1157.500000 644.410000 1158.500000 645.590000 ;
      RECT 1139.000000 644.410000 1149.500000 647.590000 ;
      RECT 386.500000 644.410000 389.000000 647.590000 ;
      RECT 372.500000 644.410000 373.500000 645.590000 ;
      RECT 357.500000 644.410000 358.500000 645.590000 ;
      RECT 0.000000 644.410000 349.500000 647.590000 ;
      RECT 1139.000000 643.590000 1158.500000 644.410000 ;
      RECT 372.500000 643.590000 389.000000 644.410000 ;
      RECT 0.000000 643.590000 358.500000 644.410000 ;
      RECT 1166.500000 642.410000 1186.000000 645.590000 ;
      RECT 1157.500000 642.410000 1158.500000 643.590000 ;
      RECT 372.500000 642.410000 373.500000 643.590000 ;
      RECT 357.500000 642.410000 358.500000 643.590000 ;
      RECT 1157.500000 641.590000 1186.000000 642.410000 ;
      RECT 357.500000 641.590000 373.500000 642.410000 ;
      RECT 1157.500000 640.410000 1158.500000 641.590000 ;
      RECT 1139.000000 640.410000 1149.500000 643.590000 ;
      RECT 386.500000 640.410000 389.000000 643.590000 ;
      RECT 372.500000 640.410000 373.500000 641.590000 ;
      RECT 357.500000 640.410000 358.500000 641.590000 ;
      RECT 0.000000 640.410000 349.500000 643.590000 ;
      RECT 1139.000000 639.590000 1158.500000 640.410000 ;
      RECT 372.500000 639.590000 389.000000 640.410000 ;
      RECT 0.000000 639.590000 358.500000 640.410000 ;
      RECT 1166.500000 638.410000 1186.000000 641.590000 ;
      RECT 1157.500000 638.410000 1158.500000 639.590000 ;
      RECT 372.500000 638.410000 373.500000 639.590000 ;
      RECT 357.500000 638.410000 358.500000 639.590000 ;
      RECT 1157.500000 637.590000 1186.000000 638.410000 ;
      RECT 357.500000 637.590000 373.500000 638.410000 ;
      RECT 1157.500000 636.410000 1158.500000 637.590000 ;
      RECT 1139.000000 636.410000 1149.500000 639.590000 ;
      RECT 386.500000 636.410000 389.000000 639.590000 ;
      RECT 372.500000 636.410000 373.500000 637.590000 ;
      RECT 357.500000 636.410000 358.500000 637.590000 ;
      RECT 0.000000 636.410000 349.500000 639.590000 ;
      RECT 1139.000000 635.590000 1158.500000 636.410000 ;
      RECT 372.500000 635.590000 389.000000 636.410000 ;
      RECT 0.000000 635.590000 358.500000 636.410000 ;
      RECT 1166.500000 634.410000 1186.000000 637.590000 ;
      RECT 1157.500000 634.410000 1158.500000 635.590000 ;
      RECT 372.500000 634.410000 373.500000 635.590000 ;
      RECT 357.500000 634.410000 358.500000 635.590000 ;
      RECT 1157.500000 633.590000 1186.000000 634.410000 ;
      RECT 357.500000 633.590000 373.500000 634.410000 ;
      RECT 1157.500000 632.410000 1158.500000 633.590000 ;
      RECT 1139.000000 632.410000 1149.500000 635.590000 ;
      RECT 386.500000 632.410000 389.000000 635.590000 ;
      RECT 372.500000 632.410000 373.500000 633.590000 ;
      RECT 357.500000 632.410000 358.500000 633.590000 ;
      RECT 0.000000 632.410000 349.500000 635.590000 ;
      RECT 1139.000000 631.590000 1158.500000 632.410000 ;
      RECT 372.500000 631.590000 389.000000 632.410000 ;
      RECT 0.000000 631.590000 358.500000 632.410000 ;
      RECT 1166.500000 630.410000 1186.000000 633.590000 ;
      RECT 1157.500000 630.410000 1158.500000 631.590000 ;
      RECT 372.500000 630.410000 373.500000 631.590000 ;
      RECT 357.500000 630.410000 358.500000 631.590000 ;
      RECT 1157.500000 629.590000 1186.000000 630.410000 ;
      RECT 357.500000 629.590000 373.500000 630.410000 ;
      RECT 1157.500000 628.410000 1158.500000 629.590000 ;
      RECT 1139.000000 628.410000 1149.500000 631.590000 ;
      RECT 386.500000 628.410000 389.000000 631.590000 ;
      RECT 372.500000 628.410000 373.500000 629.590000 ;
      RECT 357.500000 628.410000 358.500000 629.590000 ;
      RECT 0.000000 628.410000 349.500000 631.590000 ;
      RECT 1139.000000 627.590000 1158.500000 628.410000 ;
      RECT 372.500000 627.590000 389.000000 628.410000 ;
      RECT 0.000000 627.590000 358.500000 628.410000 ;
      RECT 1166.500000 626.410000 1186.000000 629.590000 ;
      RECT 1157.500000 626.410000 1158.500000 627.590000 ;
      RECT 372.500000 626.410000 373.500000 627.590000 ;
      RECT 357.500000 626.410000 358.500000 627.590000 ;
      RECT 1157.500000 625.590000 1186.000000 626.410000 ;
      RECT 357.500000 625.590000 373.500000 626.410000 ;
      RECT 1157.500000 624.410000 1158.500000 625.590000 ;
      RECT 1139.000000 624.410000 1149.500000 627.590000 ;
      RECT 386.500000 624.410000 389.000000 627.590000 ;
      RECT 372.500000 624.410000 373.500000 625.590000 ;
      RECT 357.500000 624.410000 358.500000 625.590000 ;
      RECT 0.000000 624.410000 349.500000 627.590000 ;
      RECT 1139.000000 623.590000 1158.500000 624.410000 ;
      RECT 372.500000 623.590000 389.000000 624.410000 ;
      RECT 0.000000 623.590000 358.500000 624.410000 ;
      RECT 1166.500000 622.410000 1186.000000 625.590000 ;
      RECT 1157.500000 622.410000 1158.500000 623.590000 ;
      RECT 372.500000 622.410000 373.500000 623.590000 ;
      RECT 357.500000 622.410000 358.500000 623.590000 ;
      RECT 1157.500000 621.590000 1186.000000 622.410000 ;
      RECT 357.500000 621.590000 373.500000 622.410000 ;
      RECT 1157.500000 620.410000 1158.500000 621.590000 ;
      RECT 1139.000000 620.410000 1149.500000 623.590000 ;
      RECT 386.500000 620.410000 389.000000 623.590000 ;
      RECT 372.500000 620.410000 373.500000 621.590000 ;
      RECT 357.500000 620.410000 358.500000 621.590000 ;
      RECT 0.000000 620.410000 349.500000 623.590000 ;
      RECT 1139.000000 619.590000 1158.500000 620.410000 ;
      RECT 372.500000 619.590000 389.000000 620.410000 ;
      RECT 0.000000 619.590000 358.500000 620.410000 ;
      RECT 1166.500000 618.410000 1186.000000 621.590000 ;
      RECT 1157.500000 618.410000 1158.500000 619.590000 ;
      RECT 372.500000 618.410000 373.500000 619.590000 ;
      RECT 357.500000 618.410000 358.500000 619.590000 ;
      RECT 1157.500000 617.590000 1186.000000 618.410000 ;
      RECT 357.500000 617.590000 373.500000 618.410000 ;
      RECT 1157.500000 616.410000 1158.500000 617.590000 ;
      RECT 1139.000000 616.410000 1149.500000 619.590000 ;
      RECT 386.500000 616.410000 389.000000 619.590000 ;
      RECT 372.500000 616.410000 373.500000 617.590000 ;
      RECT 357.500000 616.410000 358.500000 617.590000 ;
      RECT 0.000000 616.410000 349.500000 619.590000 ;
      RECT 1139.000000 615.590000 1158.500000 616.410000 ;
      RECT 372.500000 615.590000 389.000000 616.410000 ;
      RECT 0.000000 615.590000 358.500000 616.410000 ;
      RECT 1166.500000 614.410000 1186.000000 617.590000 ;
      RECT 1157.500000 614.410000 1158.500000 615.590000 ;
      RECT 372.500000 614.410000 373.500000 615.590000 ;
      RECT 357.500000 614.410000 358.500000 615.590000 ;
      RECT 1157.500000 613.590000 1186.000000 614.410000 ;
      RECT 357.500000 613.590000 373.500000 614.410000 ;
      RECT 1157.500000 612.410000 1158.500000 613.590000 ;
      RECT 1139.000000 612.410000 1149.500000 615.590000 ;
      RECT 386.500000 612.410000 389.000000 615.590000 ;
      RECT 372.500000 612.410000 373.500000 613.590000 ;
      RECT 357.500000 612.410000 358.500000 613.590000 ;
      RECT 0.000000 612.410000 349.500000 615.590000 ;
      RECT 1139.000000 611.590000 1158.500000 612.410000 ;
      RECT 372.500000 611.590000 389.000000 612.410000 ;
      RECT 0.000000 611.590000 358.500000 612.410000 ;
      RECT 1166.500000 610.410000 1186.000000 613.590000 ;
      RECT 1157.500000 610.410000 1158.500000 611.590000 ;
      RECT 372.500000 610.410000 373.500000 611.590000 ;
      RECT 357.500000 610.410000 358.500000 611.590000 ;
      RECT 1157.500000 609.590000 1186.000000 610.410000 ;
      RECT 357.500000 609.590000 373.500000 610.410000 ;
      RECT 1157.500000 608.410000 1158.500000 609.590000 ;
      RECT 1139.000000 608.410000 1149.500000 611.590000 ;
      RECT 386.500000 608.410000 389.000000 611.590000 ;
      RECT 372.500000 608.410000 373.500000 609.590000 ;
      RECT 357.500000 608.410000 358.500000 609.590000 ;
      RECT 0.000000 608.410000 349.500000 611.590000 ;
      RECT 1139.000000 607.590000 1158.500000 608.410000 ;
      RECT 372.500000 607.590000 389.000000 608.410000 ;
      RECT 0.000000 607.590000 358.500000 608.410000 ;
      RECT 1166.500000 606.410000 1186.000000 609.590000 ;
      RECT 1157.500000 606.410000 1158.500000 607.590000 ;
      RECT 372.500000 606.410000 373.500000 607.590000 ;
      RECT 357.500000 606.410000 358.500000 607.590000 ;
      RECT 1157.500000 605.590000 1186.000000 606.410000 ;
      RECT 357.500000 605.590000 373.500000 606.410000 ;
      RECT 1157.500000 604.410000 1158.500000 605.590000 ;
      RECT 1139.000000 604.410000 1149.500000 607.590000 ;
      RECT 386.500000 604.410000 389.000000 607.590000 ;
      RECT 372.500000 604.410000 373.500000 605.590000 ;
      RECT 357.500000 604.410000 358.500000 605.590000 ;
      RECT 0.000000 604.410000 349.500000 607.590000 ;
      RECT 1139.000000 603.590000 1158.500000 604.410000 ;
      RECT 372.500000 603.590000 389.000000 604.410000 ;
      RECT 0.000000 603.590000 358.500000 604.410000 ;
      RECT 1166.500000 602.410000 1186.000000 605.590000 ;
      RECT 1157.500000 602.410000 1158.500000 603.590000 ;
      RECT 372.500000 602.410000 373.500000 603.590000 ;
      RECT 357.500000 602.410000 358.500000 603.590000 ;
      RECT 1157.500000 601.590000 1186.000000 602.410000 ;
      RECT 357.500000 601.590000 373.500000 602.410000 ;
      RECT 1157.500000 600.410000 1158.500000 601.590000 ;
      RECT 1139.000000 600.410000 1149.500000 603.590000 ;
      RECT 386.500000 600.410000 389.000000 603.590000 ;
      RECT 372.500000 600.410000 373.500000 601.590000 ;
      RECT 357.500000 600.410000 358.500000 601.590000 ;
      RECT 0.000000 600.410000 349.500000 603.590000 ;
      RECT 1139.000000 599.590000 1158.500000 600.410000 ;
      RECT 372.500000 599.590000 389.000000 600.410000 ;
      RECT 0.000000 599.590000 358.500000 600.410000 ;
      RECT 1166.500000 598.410000 1186.000000 601.590000 ;
      RECT 1157.500000 598.410000 1158.500000 599.590000 ;
      RECT 372.500000 598.410000 373.500000 599.590000 ;
      RECT 357.500000 598.410000 358.500000 599.590000 ;
      RECT 1157.500000 597.590000 1186.000000 598.410000 ;
      RECT 357.500000 597.590000 373.500000 598.410000 ;
      RECT 1157.500000 596.410000 1158.500000 597.590000 ;
      RECT 1139.000000 596.410000 1149.500000 599.590000 ;
      RECT 386.500000 596.410000 389.000000 599.590000 ;
      RECT 372.500000 596.410000 373.500000 597.590000 ;
      RECT 357.500000 596.410000 358.500000 597.590000 ;
      RECT 0.000000 596.410000 349.500000 599.590000 ;
      RECT 1139.000000 595.590000 1158.500000 596.410000 ;
      RECT 372.500000 595.590000 389.000000 596.410000 ;
      RECT 0.000000 595.590000 358.500000 596.410000 ;
      RECT 1166.500000 594.410000 1186.000000 597.590000 ;
      RECT 1157.500000 594.410000 1158.500000 595.590000 ;
      RECT 372.500000 594.410000 373.500000 595.590000 ;
      RECT 357.500000 594.410000 358.500000 595.590000 ;
      RECT 1157.500000 593.590000 1186.000000 594.410000 ;
      RECT 357.500000 593.590000 373.500000 594.410000 ;
      RECT 1157.500000 592.410000 1158.500000 593.590000 ;
      RECT 1139.000000 592.410000 1149.500000 595.590000 ;
      RECT 386.500000 592.410000 389.000000 595.590000 ;
      RECT 372.500000 592.410000 373.500000 593.590000 ;
      RECT 357.500000 592.410000 358.500000 593.590000 ;
      RECT 0.000000 592.410000 349.500000 595.590000 ;
      RECT 1139.000000 591.590000 1158.500000 592.410000 ;
      RECT 372.500000 591.590000 389.000000 592.410000 ;
      RECT 0.000000 591.590000 358.500000 592.410000 ;
      RECT 1166.500000 590.410000 1186.000000 593.590000 ;
      RECT 1157.500000 590.410000 1158.500000 591.590000 ;
      RECT 372.500000 590.410000 373.500000 591.590000 ;
      RECT 357.500000 590.410000 358.500000 591.590000 ;
      RECT 1157.500000 589.590000 1186.000000 590.410000 ;
      RECT 357.500000 589.590000 373.500000 590.410000 ;
      RECT 1157.500000 588.410000 1158.500000 589.590000 ;
      RECT 1139.000000 588.410000 1149.500000 591.590000 ;
      RECT 386.500000 588.410000 389.000000 591.590000 ;
      RECT 372.500000 588.410000 373.500000 589.590000 ;
      RECT 357.500000 588.410000 358.500000 589.590000 ;
      RECT 0.000000 588.410000 349.500000 591.590000 ;
      RECT 1139.000000 587.590000 1158.500000 588.410000 ;
      RECT 372.500000 587.590000 389.000000 588.410000 ;
      RECT 0.000000 587.590000 358.500000 588.410000 ;
      RECT 1166.500000 586.410000 1186.000000 589.590000 ;
      RECT 1157.500000 586.410000 1158.500000 587.590000 ;
      RECT 372.500000 586.410000 373.500000 587.590000 ;
      RECT 357.500000 586.410000 358.500000 587.590000 ;
      RECT 1157.500000 585.590000 1186.000000 586.410000 ;
      RECT 357.500000 585.590000 373.500000 586.410000 ;
      RECT 1157.500000 584.410000 1158.500000 585.590000 ;
      RECT 1139.000000 584.410000 1149.500000 587.590000 ;
      RECT 386.500000 584.410000 389.000000 587.590000 ;
      RECT 372.500000 584.410000 373.500000 585.590000 ;
      RECT 357.500000 584.410000 358.500000 585.590000 ;
      RECT 0.000000 584.410000 349.500000 587.590000 ;
      RECT 1139.000000 583.590000 1158.500000 584.410000 ;
      RECT 372.500000 583.590000 389.000000 584.410000 ;
      RECT 0.000000 583.590000 358.500000 584.410000 ;
      RECT 1166.500000 582.410000 1186.000000 585.590000 ;
      RECT 1157.500000 582.410000 1158.500000 583.590000 ;
      RECT 372.500000 582.410000 373.500000 583.590000 ;
      RECT 357.500000 582.410000 358.500000 583.590000 ;
      RECT 1157.500000 581.590000 1186.000000 582.410000 ;
      RECT 357.500000 581.590000 373.500000 582.410000 ;
      RECT 1157.500000 580.410000 1158.500000 581.590000 ;
      RECT 1139.000000 580.410000 1149.500000 583.590000 ;
      RECT 386.500000 580.410000 389.000000 583.590000 ;
      RECT 372.500000 580.410000 373.500000 581.590000 ;
      RECT 357.500000 580.410000 358.500000 581.590000 ;
      RECT 0.000000 580.410000 349.500000 583.590000 ;
      RECT 1139.000000 579.590000 1158.500000 580.410000 ;
      RECT 372.500000 579.590000 389.000000 580.410000 ;
      RECT 0.000000 579.590000 358.500000 580.410000 ;
      RECT 1166.500000 578.410000 1186.000000 581.590000 ;
      RECT 1157.500000 578.410000 1158.500000 579.590000 ;
      RECT 372.500000 578.410000 373.500000 579.590000 ;
      RECT 357.500000 578.410000 358.500000 579.590000 ;
      RECT 1157.500000 577.590000 1186.000000 578.410000 ;
      RECT 357.500000 577.590000 373.500000 578.410000 ;
      RECT 1157.500000 576.410000 1158.500000 577.590000 ;
      RECT 1139.000000 576.410000 1149.500000 579.590000 ;
      RECT 386.500000 576.410000 389.000000 579.590000 ;
      RECT 372.500000 576.410000 373.500000 577.590000 ;
      RECT 357.500000 576.410000 358.500000 577.590000 ;
      RECT 0.000000 576.410000 349.500000 579.590000 ;
      RECT 1139.000000 575.590000 1158.500000 576.410000 ;
      RECT 372.500000 575.590000 389.000000 576.410000 ;
      RECT 0.000000 575.590000 358.500000 576.410000 ;
      RECT 1166.500000 574.410000 1186.000000 577.590000 ;
      RECT 1157.500000 574.410000 1158.500000 575.590000 ;
      RECT 372.500000 574.410000 373.500000 575.590000 ;
      RECT 357.500000 574.410000 358.500000 575.590000 ;
      RECT 1157.500000 573.590000 1186.000000 574.410000 ;
      RECT 357.500000 573.590000 373.500000 574.410000 ;
      RECT 1157.500000 572.410000 1158.500000 573.590000 ;
      RECT 1139.000000 572.410000 1149.500000 575.590000 ;
      RECT 386.500000 572.410000 389.000000 575.590000 ;
      RECT 372.500000 572.410000 373.500000 573.590000 ;
      RECT 357.500000 572.410000 358.500000 573.590000 ;
      RECT 0.000000 572.410000 349.500000 575.590000 ;
      RECT 1139.000000 571.590000 1158.500000 572.410000 ;
      RECT 372.500000 571.590000 389.000000 572.410000 ;
      RECT 0.000000 571.590000 358.500000 572.410000 ;
      RECT 1166.500000 570.410000 1186.000000 573.590000 ;
      RECT 1157.500000 570.410000 1158.500000 571.590000 ;
      RECT 372.500000 570.410000 373.500000 571.590000 ;
      RECT 357.500000 570.410000 358.500000 571.590000 ;
      RECT 1157.500000 569.590000 1186.000000 570.410000 ;
      RECT 357.500000 569.590000 373.500000 570.410000 ;
      RECT 1157.500000 568.410000 1158.500000 569.590000 ;
      RECT 1139.000000 568.410000 1149.500000 571.590000 ;
      RECT 386.500000 568.410000 389.000000 571.590000 ;
      RECT 372.500000 568.410000 373.500000 569.590000 ;
      RECT 357.500000 568.410000 358.500000 569.590000 ;
      RECT 0.000000 568.410000 349.500000 571.590000 ;
      RECT 1139.000000 567.590000 1158.500000 568.410000 ;
      RECT 372.500000 567.590000 389.000000 568.410000 ;
      RECT 0.000000 567.590000 358.500000 568.410000 ;
      RECT 1166.500000 566.410000 1186.000000 569.590000 ;
      RECT 1157.500000 566.410000 1158.500000 567.590000 ;
      RECT 372.500000 566.410000 373.500000 567.590000 ;
      RECT 357.500000 566.410000 358.500000 567.590000 ;
      RECT 1157.500000 565.590000 1186.000000 566.410000 ;
      RECT 357.500000 565.590000 373.500000 566.410000 ;
      RECT 1157.500000 564.410000 1158.500000 565.590000 ;
      RECT 1139.000000 564.410000 1149.500000 567.590000 ;
      RECT 386.500000 564.410000 389.000000 567.590000 ;
      RECT 372.500000 564.410000 373.500000 565.590000 ;
      RECT 357.500000 564.410000 358.500000 565.590000 ;
      RECT 0.000000 564.410000 349.500000 567.590000 ;
      RECT 1139.000000 563.590000 1158.500000 564.410000 ;
      RECT 372.500000 563.590000 389.000000 564.410000 ;
      RECT 0.000000 563.590000 358.500000 564.410000 ;
      RECT 1166.500000 562.410000 1186.000000 565.590000 ;
      RECT 1157.500000 562.410000 1158.500000 563.590000 ;
      RECT 372.500000 562.410000 373.500000 563.590000 ;
      RECT 357.500000 562.410000 358.500000 563.590000 ;
      RECT 1157.500000 561.590000 1186.000000 562.410000 ;
      RECT 357.500000 561.590000 373.500000 562.410000 ;
      RECT 1157.500000 560.410000 1158.500000 561.590000 ;
      RECT 1139.000000 560.410000 1149.500000 563.590000 ;
      RECT 386.500000 560.410000 389.000000 563.590000 ;
      RECT 372.500000 560.410000 373.500000 561.590000 ;
      RECT 357.500000 560.410000 358.500000 561.590000 ;
      RECT 0.000000 560.410000 349.500000 563.590000 ;
      RECT 1139.000000 559.590000 1158.500000 560.410000 ;
      RECT 372.500000 559.590000 389.000000 560.410000 ;
      RECT 0.000000 559.590000 358.500000 560.410000 ;
      RECT 1166.500000 558.410000 1186.000000 561.590000 ;
      RECT 1157.500000 558.410000 1158.500000 559.590000 ;
      RECT 372.500000 558.410000 373.500000 559.590000 ;
      RECT 357.500000 558.410000 358.500000 559.590000 ;
      RECT 1157.500000 557.590000 1186.000000 558.410000 ;
      RECT 357.500000 557.590000 373.500000 558.410000 ;
      RECT 1157.500000 556.410000 1158.500000 557.590000 ;
      RECT 1139.000000 556.410000 1149.500000 559.590000 ;
      RECT 386.500000 556.410000 389.000000 559.590000 ;
      RECT 372.500000 556.410000 373.500000 557.590000 ;
      RECT 357.500000 556.410000 358.500000 557.590000 ;
      RECT 0.000000 556.410000 349.500000 559.590000 ;
      RECT 1139.000000 555.590000 1158.500000 556.410000 ;
      RECT 372.500000 555.590000 389.000000 556.410000 ;
      RECT 0.000000 555.590000 358.500000 556.410000 ;
      RECT 1166.500000 554.410000 1186.000000 557.590000 ;
      RECT 1157.500000 554.410000 1158.500000 555.590000 ;
      RECT 372.500000 554.410000 373.500000 555.590000 ;
      RECT 357.500000 554.410000 358.500000 555.590000 ;
      RECT 1157.500000 553.590000 1186.000000 554.410000 ;
      RECT 357.500000 553.590000 373.500000 554.410000 ;
      RECT 1157.500000 552.410000 1158.500000 553.590000 ;
      RECT 1139.000000 552.410000 1149.500000 555.590000 ;
      RECT 386.500000 552.410000 389.000000 555.590000 ;
      RECT 372.500000 552.410000 373.500000 553.590000 ;
      RECT 357.500000 552.410000 358.500000 553.590000 ;
      RECT 0.000000 552.410000 349.500000 555.590000 ;
      RECT 1139.000000 551.590000 1158.500000 552.410000 ;
      RECT 372.500000 551.590000 389.000000 552.410000 ;
      RECT 0.000000 551.590000 358.500000 552.410000 ;
      RECT 1166.500000 550.410000 1186.000000 553.590000 ;
      RECT 1157.500000 550.410000 1158.500000 551.590000 ;
      RECT 372.500000 550.410000 373.500000 551.590000 ;
      RECT 357.500000 550.410000 358.500000 551.590000 ;
      RECT 1157.500000 549.590000 1186.000000 550.410000 ;
      RECT 357.500000 549.590000 373.500000 550.410000 ;
      RECT 1157.500000 548.410000 1158.500000 549.590000 ;
      RECT 1139.000000 548.410000 1149.500000 551.590000 ;
      RECT 386.500000 548.410000 389.000000 551.590000 ;
      RECT 372.500000 548.410000 373.500000 549.590000 ;
      RECT 357.500000 548.410000 358.500000 549.590000 ;
      RECT 0.000000 548.410000 349.500000 551.590000 ;
      RECT 1139.000000 547.590000 1158.500000 548.410000 ;
      RECT 372.500000 547.590000 389.000000 548.410000 ;
      RECT 0.000000 547.590000 358.500000 548.410000 ;
      RECT 1166.500000 546.410000 1186.000000 549.590000 ;
      RECT 1157.500000 546.410000 1158.500000 547.590000 ;
      RECT 372.500000 546.410000 373.500000 547.590000 ;
      RECT 357.500000 546.410000 358.500000 547.590000 ;
      RECT 1157.500000 545.590000 1186.000000 546.410000 ;
      RECT 357.500000 545.590000 373.500000 546.410000 ;
      RECT 1157.500000 544.410000 1158.500000 545.590000 ;
      RECT 1139.000000 544.410000 1149.500000 547.590000 ;
      RECT 386.500000 544.410000 389.000000 547.590000 ;
      RECT 372.500000 544.410000 373.500000 545.590000 ;
      RECT 357.500000 544.410000 358.500000 545.590000 ;
      RECT 0.000000 544.410000 349.500000 547.590000 ;
      RECT 1139.000000 543.590000 1158.500000 544.410000 ;
      RECT 372.500000 543.590000 389.000000 544.410000 ;
      RECT 0.000000 543.590000 358.500000 544.410000 ;
      RECT 1166.500000 542.410000 1186.000000 545.590000 ;
      RECT 1157.500000 542.410000 1158.500000 543.590000 ;
      RECT 372.500000 542.410000 373.500000 543.590000 ;
      RECT 357.500000 542.410000 358.500000 543.590000 ;
      RECT 1157.500000 541.590000 1186.000000 542.410000 ;
      RECT 357.500000 541.590000 373.500000 542.410000 ;
      RECT 1157.500000 540.410000 1158.500000 541.590000 ;
      RECT 1139.000000 540.410000 1149.500000 543.590000 ;
      RECT 386.500000 540.410000 389.000000 543.590000 ;
      RECT 372.500000 540.410000 373.500000 541.590000 ;
      RECT 357.500000 540.410000 358.500000 541.590000 ;
      RECT 0.000000 540.410000 349.500000 543.590000 ;
      RECT 1139.000000 539.590000 1158.500000 540.410000 ;
      RECT 372.500000 539.590000 389.000000 540.410000 ;
      RECT 0.000000 539.590000 358.500000 540.410000 ;
      RECT 1166.500000 538.410000 1186.000000 541.590000 ;
      RECT 1157.500000 538.410000 1158.500000 539.590000 ;
      RECT 372.500000 538.410000 373.500000 539.590000 ;
      RECT 357.500000 538.410000 358.500000 539.590000 ;
      RECT 1157.500000 537.590000 1186.000000 538.410000 ;
      RECT 357.500000 537.590000 373.500000 538.410000 ;
      RECT 1157.500000 536.410000 1158.500000 537.590000 ;
      RECT 1139.000000 536.410000 1149.500000 539.590000 ;
      RECT 386.500000 536.410000 389.000000 539.590000 ;
      RECT 372.500000 536.410000 373.500000 537.590000 ;
      RECT 357.500000 536.410000 358.500000 537.590000 ;
      RECT 0.000000 536.410000 349.500000 539.590000 ;
      RECT 1139.000000 535.590000 1158.500000 536.410000 ;
      RECT 372.500000 535.590000 389.000000 536.410000 ;
      RECT 0.000000 535.590000 358.500000 536.410000 ;
      RECT 1166.500000 534.410000 1186.000000 537.590000 ;
      RECT 1157.500000 534.410000 1158.500000 535.590000 ;
      RECT 372.500000 534.410000 373.500000 535.590000 ;
      RECT 357.500000 534.410000 358.500000 535.590000 ;
      RECT 1157.500000 533.590000 1186.000000 534.410000 ;
      RECT 357.500000 533.590000 373.500000 534.410000 ;
      RECT 1157.500000 532.410000 1158.500000 533.590000 ;
      RECT 1139.000000 532.410000 1149.500000 535.590000 ;
      RECT 386.500000 532.410000 389.000000 535.590000 ;
      RECT 372.500000 532.410000 373.500000 533.590000 ;
      RECT 357.500000 532.410000 358.500000 533.590000 ;
      RECT 0.000000 532.410000 349.500000 535.590000 ;
      RECT 1139.000000 531.590000 1158.500000 532.410000 ;
      RECT 372.500000 531.590000 389.000000 532.410000 ;
      RECT 0.000000 531.590000 358.500000 532.410000 ;
      RECT 1166.500000 530.410000 1186.000000 533.590000 ;
      RECT 1157.500000 530.410000 1158.500000 531.590000 ;
      RECT 372.500000 530.410000 373.500000 531.590000 ;
      RECT 357.500000 530.410000 358.500000 531.590000 ;
      RECT 1157.500000 529.590000 1186.000000 530.410000 ;
      RECT 357.500000 529.590000 373.500000 530.410000 ;
      RECT 1157.500000 528.410000 1158.500000 529.590000 ;
      RECT 1139.000000 528.410000 1149.500000 531.590000 ;
      RECT 386.500000 528.410000 389.000000 531.590000 ;
      RECT 372.500000 528.410000 373.500000 529.590000 ;
      RECT 357.500000 528.410000 358.500000 529.590000 ;
      RECT 0.000000 528.410000 349.500000 531.590000 ;
      RECT 1139.000000 527.590000 1158.500000 528.410000 ;
      RECT 372.500000 527.590000 389.000000 528.410000 ;
      RECT 0.000000 527.590000 358.500000 528.410000 ;
      RECT 1166.500000 526.410000 1186.000000 529.590000 ;
      RECT 1157.500000 526.410000 1158.500000 527.590000 ;
      RECT 372.500000 526.410000 373.500000 527.590000 ;
      RECT 357.500000 526.410000 358.500000 527.590000 ;
      RECT 1157.500000 525.590000 1186.000000 526.410000 ;
      RECT 357.500000 525.590000 373.500000 526.410000 ;
      RECT 1157.500000 524.410000 1158.500000 525.590000 ;
      RECT 1139.000000 524.410000 1149.500000 527.590000 ;
      RECT 386.500000 524.410000 389.000000 527.590000 ;
      RECT 372.500000 524.410000 373.500000 525.590000 ;
      RECT 357.500000 524.410000 358.500000 525.590000 ;
      RECT 0.000000 524.410000 349.500000 527.590000 ;
      RECT 1139.000000 523.590000 1158.500000 524.410000 ;
      RECT 372.500000 523.590000 389.000000 524.410000 ;
      RECT 0.000000 523.590000 358.500000 524.410000 ;
      RECT 1166.500000 522.410000 1186.000000 525.590000 ;
      RECT 1157.500000 522.410000 1158.500000 523.590000 ;
      RECT 372.500000 522.410000 373.500000 523.590000 ;
      RECT 357.500000 522.410000 358.500000 523.590000 ;
      RECT 1157.500000 521.590000 1186.000000 522.410000 ;
      RECT 357.500000 521.590000 373.500000 522.410000 ;
      RECT 1157.500000 520.410000 1158.500000 521.590000 ;
      RECT 1139.000000 520.410000 1149.500000 523.590000 ;
      RECT 386.500000 520.410000 389.000000 523.590000 ;
      RECT 372.500000 520.410000 373.500000 521.590000 ;
      RECT 357.500000 520.410000 358.500000 521.590000 ;
      RECT 0.000000 520.410000 349.500000 523.590000 ;
      RECT 1139.000000 519.590000 1158.500000 520.410000 ;
      RECT 372.500000 519.590000 389.000000 520.410000 ;
      RECT 0.000000 519.590000 358.500000 520.410000 ;
      RECT 1166.500000 518.410000 1186.000000 521.590000 ;
      RECT 1157.500000 518.410000 1158.500000 519.590000 ;
      RECT 372.500000 518.410000 373.500000 519.590000 ;
      RECT 357.500000 518.410000 358.500000 519.590000 ;
      RECT 1157.500000 517.590000 1186.000000 518.410000 ;
      RECT 357.500000 517.590000 373.500000 518.410000 ;
      RECT 307.500000 517.590000 349.500000 519.590000 ;
      RECT 0.000000 517.590000 299.500000 519.590000 ;
      RECT 1157.500000 516.410000 1158.500000 517.590000 ;
      RECT 1139.000000 516.410000 1149.500000 519.590000 ;
      RECT 386.500000 516.410000 389.000000 519.590000 ;
      RECT 372.500000 516.410000 373.500000 517.590000 ;
      RECT 357.500000 516.410000 358.500000 517.590000 ;
      RECT 316.500000 516.410000 349.500000 517.590000 ;
      RECT 307.500000 516.410000 308.500000 517.590000 ;
      RECT 266.500000 516.410000 299.500000 517.590000 ;
      RECT 1139.000000 515.590000 1158.500000 516.410000 ;
      RECT 372.500000 515.590000 389.000000 516.410000 ;
      RECT 316.500000 515.590000 358.500000 516.410000 ;
      RECT 266.500000 515.590000 308.500000 516.410000 ;
      RECT 216.500000 515.590000 258.500000 517.590000 ;
      RECT 166.500000 515.590000 208.500000 517.590000 ;
      RECT 116.500000 515.590000 158.500000 517.590000 ;
      RECT 66.500000 515.590000 108.500000 517.590000 ;
      RECT 29.500000 515.590000 58.500000 517.590000 ;
      RECT 0.000000 515.590000 16.500000 517.590000 ;
      RECT 1166.500000 514.410000 1186.000000 517.590000 ;
      RECT 1157.500000 514.410000 1158.500000 515.590000 ;
      RECT 372.500000 514.410000 373.500000 515.590000 ;
      RECT 357.500000 514.410000 358.500000 515.590000 ;
      RECT 316.500000 514.410000 349.500000 515.590000 ;
      RECT 307.500000 514.410000 308.500000 515.590000 ;
      RECT 266.500000 514.410000 299.500000 515.590000 ;
      RECT 257.500000 514.410000 258.500000 515.590000 ;
      RECT 216.500000 514.410000 249.500000 515.590000 ;
      RECT 207.500000 514.410000 208.500000 515.590000 ;
      RECT 166.500000 514.410000 199.500000 515.590000 ;
      RECT 157.500000 514.410000 158.500000 515.590000 ;
      RECT 116.500000 514.410000 149.500000 515.590000 ;
      RECT 107.500000 514.410000 108.500000 515.590000 ;
      RECT 66.500000 514.410000 99.500000 515.590000 ;
      RECT 57.500000 514.410000 58.500000 515.590000 ;
      RECT 29.500000 514.410000 49.500000 515.590000 ;
      RECT 15.500000 514.410000 16.500000 515.590000 ;
      RECT 1157.500000 513.590000 1186.000000 514.410000 ;
      RECT 357.500000 513.590000 373.500000 514.410000 ;
      RECT 307.500000 513.590000 349.500000 514.410000 ;
      RECT 257.500000 513.590000 299.500000 514.410000 ;
      RECT 207.500000 513.590000 249.500000 514.410000 ;
      RECT 157.500000 513.590000 199.500000 514.410000 ;
      RECT 107.500000 513.590000 149.500000 514.410000 ;
      RECT 57.500000 513.590000 99.500000 514.410000 ;
      RECT 15.500000 513.590000 49.500000 514.410000 ;
      RECT 1157.500000 512.410000 1158.500000 513.590000 ;
      RECT 1139.000000 512.410000 1149.500000 515.590000 ;
      RECT 386.500000 512.410000 389.000000 515.590000 ;
      RECT 372.500000 512.410000 373.500000 513.590000 ;
      RECT 357.500000 512.410000 358.500000 513.590000 ;
      RECT 316.500000 512.410000 349.500000 513.590000 ;
      RECT 307.500000 512.410000 308.500000 513.590000 ;
      RECT 266.500000 512.410000 299.500000 513.590000 ;
      RECT 257.500000 512.410000 258.500000 513.590000 ;
      RECT 216.500000 512.410000 249.500000 513.590000 ;
      RECT 207.500000 512.410000 208.500000 513.590000 ;
      RECT 166.500000 512.410000 199.500000 513.590000 ;
      RECT 157.500000 512.410000 158.500000 513.590000 ;
      RECT 116.500000 512.410000 149.500000 513.590000 ;
      RECT 107.500000 512.410000 108.500000 513.590000 ;
      RECT 66.500000 512.410000 99.500000 513.590000 ;
      RECT 57.500000 512.410000 58.500000 513.590000 ;
      RECT 29.500000 512.410000 49.500000 513.590000 ;
      RECT 15.500000 512.410000 16.500000 513.590000 ;
      RECT 0.000000 512.410000 2.500000 515.590000 ;
      RECT 1139.000000 511.590000 1158.500000 512.410000 ;
      RECT 372.500000 511.590000 389.000000 512.410000 ;
      RECT 316.500000 511.590000 358.500000 512.410000 ;
      RECT 266.500000 511.590000 308.500000 512.410000 ;
      RECT 216.500000 511.590000 258.500000 512.410000 ;
      RECT 166.500000 511.590000 208.500000 512.410000 ;
      RECT 116.500000 511.590000 158.500000 512.410000 ;
      RECT 66.500000 511.590000 108.500000 512.410000 ;
      RECT 29.500000 511.590000 58.500000 512.410000 ;
      RECT 0.000000 511.590000 16.500000 512.410000 ;
      RECT 1166.500000 510.410000 1186.000000 513.590000 ;
      RECT 1157.500000 510.410000 1158.500000 511.590000 ;
      RECT 372.500000 510.410000 373.500000 511.590000 ;
      RECT 357.500000 510.410000 358.500000 511.590000 ;
      RECT 316.500000 510.410000 349.500000 511.590000 ;
      RECT 307.500000 510.410000 308.500000 511.590000 ;
      RECT 266.500000 510.410000 299.500000 511.590000 ;
      RECT 257.500000 510.410000 258.500000 511.590000 ;
      RECT 216.500000 510.410000 249.500000 511.590000 ;
      RECT 207.500000 510.410000 208.500000 511.590000 ;
      RECT 166.500000 510.410000 199.500000 511.590000 ;
      RECT 157.500000 510.410000 158.500000 511.590000 ;
      RECT 116.500000 510.410000 149.500000 511.590000 ;
      RECT 107.500000 510.410000 108.500000 511.590000 ;
      RECT 66.500000 510.410000 99.500000 511.590000 ;
      RECT 57.500000 510.410000 58.500000 511.590000 ;
      RECT 29.500000 510.410000 49.500000 511.590000 ;
      RECT 15.500000 510.410000 16.500000 511.590000 ;
      RECT 1157.500000 509.590000 1186.000000 510.410000 ;
      RECT 357.500000 509.590000 373.500000 510.410000 ;
      RECT 307.500000 509.590000 349.500000 510.410000 ;
      RECT 257.500000 509.590000 299.500000 510.410000 ;
      RECT 207.500000 509.590000 249.500000 510.410000 ;
      RECT 157.500000 509.590000 199.500000 510.410000 ;
      RECT 107.500000 509.590000 149.500000 510.410000 ;
      RECT 57.500000 509.590000 99.500000 510.410000 ;
      RECT 15.500000 509.590000 49.500000 510.410000 ;
      RECT 1157.500000 508.410000 1158.500000 509.590000 ;
      RECT 1139.000000 508.410000 1149.500000 511.590000 ;
      RECT 386.500000 508.410000 389.000000 511.590000 ;
      RECT 372.500000 508.410000 373.500000 509.590000 ;
      RECT 357.500000 508.410000 358.500000 509.590000 ;
      RECT 316.500000 508.410000 349.500000 509.590000 ;
      RECT 307.500000 508.410000 308.500000 509.590000 ;
      RECT 266.500000 508.410000 299.500000 509.590000 ;
      RECT 257.500000 508.410000 258.500000 509.590000 ;
      RECT 216.500000 508.410000 249.500000 509.590000 ;
      RECT 207.500000 508.410000 208.500000 509.590000 ;
      RECT 166.500000 508.410000 199.500000 509.590000 ;
      RECT 157.500000 508.410000 158.500000 509.590000 ;
      RECT 116.500000 508.410000 149.500000 509.590000 ;
      RECT 107.500000 508.410000 108.500000 509.590000 ;
      RECT 66.500000 508.410000 99.500000 509.590000 ;
      RECT 57.500000 508.410000 58.500000 509.590000 ;
      RECT 29.500000 508.410000 49.500000 509.590000 ;
      RECT 15.500000 508.410000 16.500000 509.590000 ;
      RECT 0.000000 508.410000 2.500000 511.590000 ;
      RECT 1139.000000 507.590000 1158.500000 508.410000 ;
      RECT 372.500000 507.590000 389.000000 508.410000 ;
      RECT 316.500000 507.590000 358.500000 508.410000 ;
      RECT 266.500000 507.590000 308.500000 508.410000 ;
      RECT 216.500000 507.590000 258.500000 508.410000 ;
      RECT 166.500000 507.590000 208.500000 508.410000 ;
      RECT 116.500000 507.590000 158.500000 508.410000 ;
      RECT 66.500000 507.590000 108.500000 508.410000 ;
      RECT 29.500000 507.590000 58.500000 508.410000 ;
      RECT 0.000000 507.590000 16.500000 508.410000 ;
      RECT 1166.500000 506.410000 1186.000000 509.590000 ;
      RECT 1157.500000 506.410000 1158.500000 507.590000 ;
      RECT 372.500000 506.410000 373.500000 507.590000 ;
      RECT 357.500000 506.410000 358.500000 507.590000 ;
      RECT 316.500000 506.410000 349.500000 507.590000 ;
      RECT 307.500000 506.410000 308.500000 507.590000 ;
      RECT 266.500000 506.410000 299.500000 507.590000 ;
      RECT 257.500000 506.410000 258.500000 507.590000 ;
      RECT 216.500000 506.410000 249.500000 507.590000 ;
      RECT 207.500000 506.410000 208.500000 507.590000 ;
      RECT 166.500000 506.410000 199.500000 507.590000 ;
      RECT 157.500000 506.410000 158.500000 507.590000 ;
      RECT 116.500000 506.410000 149.500000 507.590000 ;
      RECT 107.500000 506.410000 108.500000 507.590000 ;
      RECT 66.500000 506.410000 99.500000 507.590000 ;
      RECT 57.500000 506.410000 58.500000 507.590000 ;
      RECT 29.500000 506.410000 49.500000 507.590000 ;
      RECT 15.500000 506.410000 16.500000 507.590000 ;
      RECT 386.500000 506.000000 389.000000 507.590000 ;
      RECT 1157.500000 505.590000 1186.000000 506.410000 ;
      RECT 386.500000 505.590000 739.000000 506.000000 ;
      RECT 357.500000 505.590000 373.500000 506.410000 ;
      RECT 307.500000 505.590000 349.500000 506.410000 ;
      RECT 257.500000 505.590000 299.500000 506.410000 ;
      RECT 207.500000 505.590000 249.500000 506.410000 ;
      RECT 157.500000 505.590000 199.500000 506.410000 ;
      RECT 107.500000 505.590000 149.500000 506.410000 ;
      RECT 57.500000 505.590000 99.500000 506.410000 ;
      RECT 15.500000 505.590000 49.500000 506.410000 ;
      RECT 1157.500000 504.410000 1158.500000 505.590000 ;
      RECT 1139.000000 504.410000 1149.500000 507.590000 ;
      RECT 386.500000 504.410000 408.500000 505.590000 ;
      RECT 372.500000 504.410000 373.500000 505.590000 ;
      RECT 357.500000 504.410000 358.500000 505.590000 ;
      RECT 316.500000 504.410000 349.500000 505.590000 ;
      RECT 307.500000 504.410000 308.500000 505.590000 ;
      RECT 266.500000 504.410000 299.500000 505.590000 ;
      RECT 257.500000 504.410000 258.500000 505.590000 ;
      RECT 216.500000 504.410000 249.500000 505.590000 ;
      RECT 207.500000 504.410000 208.500000 505.590000 ;
      RECT 166.500000 504.410000 199.500000 505.590000 ;
      RECT 157.500000 504.410000 158.500000 505.590000 ;
      RECT 116.500000 504.410000 149.500000 505.590000 ;
      RECT 107.500000 504.410000 108.500000 505.590000 ;
      RECT 66.500000 504.410000 99.500000 505.590000 ;
      RECT 57.500000 504.410000 58.500000 505.590000 ;
      RECT 29.500000 504.410000 49.500000 505.590000 ;
      RECT 15.500000 504.410000 16.500000 505.590000 ;
      RECT 0.000000 504.410000 2.500000 507.590000 ;
      RECT 1139.000000 503.590000 1158.500000 504.410000 ;
      RECT 716.500000 503.590000 739.000000 505.590000 ;
      RECT 666.500000 503.590000 708.500000 505.590000 ;
      RECT 616.500000 503.590000 658.500000 505.590000 ;
      RECT 566.500000 503.590000 608.500000 505.590000 ;
      RECT 516.500000 503.590000 558.500000 505.590000 ;
      RECT 466.500000 503.590000 508.500000 505.590000 ;
      RECT 416.500000 503.590000 458.500000 505.590000 ;
      RECT 372.500000 503.590000 408.500000 504.410000 ;
      RECT 316.500000 503.590000 358.500000 504.410000 ;
      RECT 266.500000 503.590000 308.500000 504.410000 ;
      RECT 216.500000 503.590000 258.500000 504.410000 ;
      RECT 166.500000 503.590000 208.500000 504.410000 ;
      RECT 116.500000 503.590000 158.500000 504.410000 ;
      RECT 66.500000 503.590000 108.500000 504.410000 ;
      RECT 29.500000 503.590000 58.500000 504.410000 ;
      RECT 0.000000 503.590000 16.500000 504.410000 ;
      RECT 1166.500000 502.410000 1186.000000 505.590000 ;
      RECT 1157.500000 502.410000 1158.500000 503.590000 ;
      RECT 716.500000 502.410000 723.500000 503.590000 ;
      RECT 707.500000 502.410000 708.500000 503.590000 ;
      RECT 666.500000 502.410000 699.500000 503.590000 ;
      RECT 657.500000 502.410000 658.500000 503.590000 ;
      RECT 616.500000 502.410000 649.500000 503.590000 ;
      RECT 607.500000 502.410000 608.500000 503.590000 ;
      RECT 566.500000 502.410000 599.500000 503.590000 ;
      RECT 557.500000 502.410000 558.500000 503.590000 ;
      RECT 516.500000 502.410000 549.500000 503.590000 ;
      RECT 507.500000 502.410000 508.500000 503.590000 ;
      RECT 466.500000 502.410000 499.500000 503.590000 ;
      RECT 457.500000 502.410000 458.500000 503.590000 ;
      RECT 416.500000 502.410000 449.500000 503.590000 ;
      RECT 407.500000 502.410000 408.500000 503.590000 ;
      RECT 372.500000 502.410000 373.500000 503.590000 ;
      RECT 357.500000 502.410000 358.500000 503.590000 ;
      RECT 316.500000 502.410000 349.500000 503.590000 ;
      RECT 307.500000 502.410000 308.500000 503.590000 ;
      RECT 266.500000 502.410000 299.500000 503.590000 ;
      RECT 257.500000 502.410000 258.500000 503.590000 ;
      RECT 216.500000 502.410000 249.500000 503.590000 ;
      RECT 207.500000 502.410000 208.500000 503.590000 ;
      RECT 166.500000 502.410000 199.500000 503.590000 ;
      RECT 157.500000 502.410000 158.500000 503.590000 ;
      RECT 116.500000 502.410000 149.500000 503.590000 ;
      RECT 107.500000 502.410000 108.500000 503.590000 ;
      RECT 66.500000 502.410000 99.500000 503.590000 ;
      RECT 57.500000 502.410000 58.500000 503.590000 ;
      RECT 29.500000 502.410000 49.500000 503.590000 ;
      RECT 15.500000 502.410000 16.500000 503.590000 ;
      RECT 1157.500000 501.590000 1186.000000 502.410000 ;
      RECT 707.500000 501.590000 723.500000 502.410000 ;
      RECT 657.500000 501.590000 699.500000 502.410000 ;
      RECT 607.500000 501.590000 649.500000 502.410000 ;
      RECT 557.500000 501.590000 599.500000 502.410000 ;
      RECT 507.500000 501.590000 549.500000 502.410000 ;
      RECT 457.500000 501.590000 499.500000 502.410000 ;
      RECT 407.500000 501.590000 449.500000 502.410000 ;
      RECT 357.500000 501.590000 373.500000 502.410000 ;
      RECT 307.500000 501.590000 349.500000 502.410000 ;
      RECT 257.500000 501.590000 299.500000 502.410000 ;
      RECT 207.500000 501.590000 249.500000 502.410000 ;
      RECT 157.500000 501.590000 199.500000 502.410000 ;
      RECT 107.500000 501.590000 149.500000 502.410000 ;
      RECT 57.500000 501.590000 99.500000 502.410000 ;
      RECT 15.500000 501.590000 49.500000 502.410000 ;
      RECT 1157.500000 500.410000 1158.500000 501.590000 ;
      RECT 1139.000000 500.410000 1149.500000 503.590000 ;
      RECT 736.500000 500.410000 739.000000 503.590000 ;
      RECT 716.500000 500.410000 723.500000 501.590000 ;
      RECT 707.500000 500.410000 708.500000 501.590000 ;
      RECT 666.500000 500.410000 699.500000 501.590000 ;
      RECT 657.500000 500.410000 658.500000 501.590000 ;
      RECT 616.500000 500.410000 649.500000 501.590000 ;
      RECT 607.500000 500.410000 608.500000 501.590000 ;
      RECT 566.500000 500.410000 599.500000 501.590000 ;
      RECT 557.500000 500.410000 558.500000 501.590000 ;
      RECT 516.500000 500.410000 549.500000 501.590000 ;
      RECT 507.500000 500.410000 508.500000 501.590000 ;
      RECT 466.500000 500.410000 499.500000 501.590000 ;
      RECT 457.500000 500.410000 458.500000 501.590000 ;
      RECT 416.500000 500.410000 449.500000 501.590000 ;
      RECT 407.500000 500.410000 408.500000 501.590000 ;
      RECT 386.500000 500.410000 399.500000 503.590000 ;
      RECT 372.500000 500.410000 373.500000 501.590000 ;
      RECT 357.500000 500.410000 358.500000 501.590000 ;
      RECT 316.500000 500.410000 349.500000 501.590000 ;
      RECT 307.500000 500.410000 308.500000 501.590000 ;
      RECT 266.500000 500.410000 299.500000 501.590000 ;
      RECT 257.500000 500.410000 258.500000 501.590000 ;
      RECT 216.500000 500.410000 249.500000 501.590000 ;
      RECT 207.500000 500.410000 208.500000 501.590000 ;
      RECT 166.500000 500.410000 199.500000 501.590000 ;
      RECT 157.500000 500.410000 158.500000 501.590000 ;
      RECT 116.500000 500.410000 149.500000 501.590000 ;
      RECT 107.500000 500.410000 108.500000 501.590000 ;
      RECT 66.500000 500.410000 99.500000 501.590000 ;
      RECT 57.500000 500.410000 58.500000 501.590000 ;
      RECT 29.500000 500.410000 49.500000 501.590000 ;
      RECT 15.500000 500.410000 16.500000 501.590000 ;
      RECT 0.000000 500.410000 2.500000 503.590000 ;
      RECT 1139.000000 499.590000 1158.500000 500.410000 ;
      RECT 716.500000 499.590000 739.000000 500.410000 ;
      RECT 666.500000 499.590000 708.500000 500.410000 ;
      RECT 616.500000 499.590000 658.500000 500.410000 ;
      RECT 566.500000 499.590000 608.500000 500.410000 ;
      RECT 516.500000 499.590000 558.500000 500.410000 ;
      RECT 466.500000 499.590000 508.500000 500.410000 ;
      RECT 416.500000 499.590000 458.500000 500.410000 ;
      RECT 372.500000 499.590000 408.500000 500.410000 ;
      RECT 316.500000 499.590000 358.500000 500.410000 ;
      RECT 266.500000 499.590000 308.500000 500.410000 ;
      RECT 216.500000 499.590000 258.500000 500.410000 ;
      RECT 166.500000 499.590000 208.500000 500.410000 ;
      RECT 116.500000 499.590000 158.500000 500.410000 ;
      RECT 66.500000 499.590000 108.500000 500.410000 ;
      RECT 29.500000 499.590000 58.500000 500.410000 ;
      RECT 0.000000 499.590000 16.500000 500.410000 ;
      RECT 1166.500000 498.410000 1186.000000 501.590000 ;
      RECT 1157.500000 498.410000 1158.500000 499.590000 ;
      RECT 716.500000 498.410000 723.500000 499.590000 ;
      RECT 707.500000 498.410000 708.500000 499.590000 ;
      RECT 666.500000 498.410000 699.500000 499.590000 ;
      RECT 657.500000 498.410000 658.500000 499.590000 ;
      RECT 616.500000 498.410000 649.500000 499.590000 ;
      RECT 607.500000 498.410000 608.500000 499.590000 ;
      RECT 566.500000 498.410000 599.500000 499.590000 ;
      RECT 557.500000 498.410000 558.500000 499.590000 ;
      RECT 516.500000 498.410000 549.500000 499.590000 ;
      RECT 507.500000 498.410000 508.500000 499.590000 ;
      RECT 466.500000 498.410000 499.500000 499.590000 ;
      RECT 457.500000 498.410000 458.500000 499.590000 ;
      RECT 416.500000 498.410000 449.500000 499.590000 ;
      RECT 407.500000 498.410000 408.500000 499.590000 ;
      RECT 372.500000 498.410000 373.500000 499.590000 ;
      RECT 357.500000 498.410000 358.500000 499.590000 ;
      RECT 316.500000 498.410000 349.500000 499.590000 ;
      RECT 307.500000 498.410000 308.500000 499.590000 ;
      RECT 266.500000 498.410000 299.500000 499.590000 ;
      RECT 257.500000 498.410000 258.500000 499.590000 ;
      RECT 216.500000 498.410000 249.500000 499.590000 ;
      RECT 207.500000 498.410000 208.500000 499.590000 ;
      RECT 166.500000 498.410000 199.500000 499.590000 ;
      RECT 157.500000 498.410000 158.500000 499.590000 ;
      RECT 116.500000 498.410000 149.500000 499.590000 ;
      RECT 107.500000 498.410000 108.500000 499.590000 ;
      RECT 66.500000 498.410000 99.500000 499.590000 ;
      RECT 57.500000 498.410000 58.500000 499.590000 ;
      RECT 29.500000 498.410000 49.500000 499.590000 ;
      RECT 15.500000 498.410000 16.500000 499.590000 ;
      RECT 1157.500000 497.590000 1186.000000 498.410000 ;
      RECT 707.500000 497.590000 723.500000 498.410000 ;
      RECT 657.500000 497.590000 699.500000 498.410000 ;
      RECT 607.500000 497.590000 649.500000 498.410000 ;
      RECT 557.500000 497.590000 599.500000 498.410000 ;
      RECT 507.500000 497.590000 549.500000 498.410000 ;
      RECT 457.500000 497.590000 499.500000 498.410000 ;
      RECT 407.500000 497.590000 449.500000 498.410000 ;
      RECT 357.500000 497.590000 373.500000 498.410000 ;
      RECT 307.500000 497.590000 349.500000 498.410000 ;
      RECT 257.500000 497.590000 299.500000 498.410000 ;
      RECT 207.500000 497.590000 249.500000 498.410000 ;
      RECT 157.500000 497.590000 199.500000 498.410000 ;
      RECT 107.500000 497.590000 149.500000 498.410000 ;
      RECT 57.500000 497.590000 99.500000 498.410000 ;
      RECT 15.500000 497.590000 49.500000 498.410000 ;
      RECT 1157.500000 496.410000 1158.500000 497.590000 ;
      RECT 1139.000000 496.410000 1149.500000 499.590000 ;
      RECT 736.500000 496.410000 739.000000 499.590000 ;
      RECT 716.500000 496.410000 723.500000 497.590000 ;
      RECT 707.500000 496.410000 708.500000 497.590000 ;
      RECT 666.500000 496.410000 699.500000 497.590000 ;
      RECT 657.500000 496.410000 658.500000 497.590000 ;
      RECT 616.500000 496.410000 649.500000 497.590000 ;
      RECT 607.500000 496.410000 608.500000 497.590000 ;
      RECT 566.500000 496.410000 599.500000 497.590000 ;
      RECT 557.500000 496.410000 558.500000 497.590000 ;
      RECT 516.500000 496.410000 549.500000 497.590000 ;
      RECT 507.500000 496.410000 508.500000 497.590000 ;
      RECT 466.500000 496.410000 499.500000 497.590000 ;
      RECT 457.500000 496.410000 458.500000 497.590000 ;
      RECT 416.500000 496.410000 449.500000 497.590000 ;
      RECT 407.500000 496.410000 408.500000 497.590000 ;
      RECT 386.500000 496.410000 399.500000 499.590000 ;
      RECT 372.500000 496.410000 373.500000 497.590000 ;
      RECT 357.500000 496.410000 358.500000 497.590000 ;
      RECT 316.500000 496.410000 349.500000 497.590000 ;
      RECT 307.500000 496.410000 308.500000 497.590000 ;
      RECT 266.500000 496.410000 299.500000 497.590000 ;
      RECT 257.500000 496.410000 258.500000 497.590000 ;
      RECT 216.500000 496.410000 249.500000 497.590000 ;
      RECT 207.500000 496.410000 208.500000 497.590000 ;
      RECT 166.500000 496.410000 199.500000 497.590000 ;
      RECT 157.500000 496.410000 158.500000 497.590000 ;
      RECT 116.500000 496.410000 149.500000 497.590000 ;
      RECT 107.500000 496.410000 108.500000 497.590000 ;
      RECT 66.500000 496.410000 99.500000 497.590000 ;
      RECT 57.500000 496.410000 58.500000 497.590000 ;
      RECT 29.500000 496.410000 49.500000 497.590000 ;
      RECT 15.500000 496.410000 16.500000 497.590000 ;
      RECT 0.000000 496.410000 2.500000 499.590000 ;
      RECT 1139.000000 495.590000 1158.500000 496.410000 ;
      RECT 716.500000 495.590000 739.000000 496.410000 ;
      RECT 666.500000 495.590000 708.500000 496.410000 ;
      RECT 616.500000 495.590000 658.500000 496.410000 ;
      RECT 566.500000 495.590000 608.500000 496.410000 ;
      RECT 516.500000 495.590000 558.500000 496.410000 ;
      RECT 466.500000 495.590000 508.500000 496.410000 ;
      RECT 416.500000 495.590000 458.500000 496.410000 ;
      RECT 372.500000 495.590000 408.500000 496.410000 ;
      RECT 316.500000 495.590000 358.500000 496.410000 ;
      RECT 266.500000 495.590000 308.500000 496.410000 ;
      RECT 216.500000 495.590000 258.500000 496.410000 ;
      RECT 166.500000 495.590000 208.500000 496.410000 ;
      RECT 116.500000 495.590000 158.500000 496.410000 ;
      RECT 66.500000 495.590000 108.500000 496.410000 ;
      RECT 29.500000 495.590000 58.500000 496.410000 ;
      RECT 0.000000 495.590000 16.500000 496.410000 ;
      RECT 1166.500000 494.410000 1186.000000 497.590000 ;
      RECT 1157.500000 494.410000 1158.500000 495.590000 ;
      RECT 716.500000 494.410000 723.500000 495.590000 ;
      RECT 707.500000 494.410000 708.500000 495.590000 ;
      RECT 666.500000 494.410000 699.500000 495.590000 ;
      RECT 657.500000 494.410000 658.500000 495.590000 ;
      RECT 616.500000 494.410000 649.500000 495.590000 ;
      RECT 607.500000 494.410000 608.500000 495.590000 ;
      RECT 566.500000 494.410000 599.500000 495.590000 ;
      RECT 557.500000 494.410000 558.500000 495.590000 ;
      RECT 516.500000 494.410000 549.500000 495.590000 ;
      RECT 507.500000 494.410000 508.500000 495.590000 ;
      RECT 466.500000 494.410000 499.500000 495.590000 ;
      RECT 457.500000 494.410000 458.500000 495.590000 ;
      RECT 416.500000 494.410000 449.500000 495.590000 ;
      RECT 407.500000 494.410000 408.500000 495.590000 ;
      RECT 372.500000 494.410000 373.500000 495.590000 ;
      RECT 357.500000 494.410000 358.500000 495.590000 ;
      RECT 316.500000 494.410000 349.500000 495.590000 ;
      RECT 307.500000 494.410000 308.500000 495.590000 ;
      RECT 266.500000 494.410000 299.500000 495.590000 ;
      RECT 257.500000 494.410000 258.500000 495.590000 ;
      RECT 216.500000 494.410000 249.500000 495.590000 ;
      RECT 207.500000 494.410000 208.500000 495.590000 ;
      RECT 166.500000 494.410000 199.500000 495.590000 ;
      RECT 157.500000 494.410000 158.500000 495.590000 ;
      RECT 116.500000 494.410000 149.500000 495.590000 ;
      RECT 107.500000 494.410000 108.500000 495.590000 ;
      RECT 66.500000 494.410000 99.500000 495.590000 ;
      RECT 57.500000 494.410000 58.500000 495.590000 ;
      RECT 29.500000 494.410000 49.500000 495.590000 ;
      RECT 15.500000 494.410000 16.500000 495.590000 ;
      RECT 1157.500000 493.590000 1186.000000 494.410000 ;
      RECT 707.500000 493.590000 723.500000 494.410000 ;
      RECT 657.500000 493.590000 699.500000 494.410000 ;
      RECT 607.500000 493.590000 649.500000 494.410000 ;
      RECT 557.500000 493.590000 599.500000 494.410000 ;
      RECT 507.500000 493.590000 549.500000 494.410000 ;
      RECT 457.500000 493.590000 499.500000 494.410000 ;
      RECT 407.500000 493.590000 449.500000 494.410000 ;
      RECT 357.500000 493.590000 373.500000 494.410000 ;
      RECT 307.500000 493.590000 349.500000 494.410000 ;
      RECT 257.500000 493.590000 299.500000 494.410000 ;
      RECT 207.500000 493.590000 249.500000 494.410000 ;
      RECT 157.500000 493.590000 199.500000 494.410000 ;
      RECT 107.500000 493.590000 149.500000 494.410000 ;
      RECT 57.500000 493.590000 99.500000 494.410000 ;
      RECT 15.500000 493.590000 49.500000 494.410000 ;
      RECT 1157.500000 492.410000 1158.500000 493.590000 ;
      RECT 1139.000000 492.410000 1149.500000 495.590000 ;
      RECT 736.500000 492.410000 739.000000 495.590000 ;
      RECT 716.500000 492.410000 723.500000 493.590000 ;
      RECT 707.500000 492.410000 708.500000 493.590000 ;
      RECT 666.500000 492.410000 699.500000 493.590000 ;
      RECT 657.500000 492.410000 658.500000 493.590000 ;
      RECT 616.500000 492.410000 649.500000 493.590000 ;
      RECT 607.500000 492.410000 608.500000 493.590000 ;
      RECT 566.500000 492.410000 599.500000 493.590000 ;
      RECT 557.500000 492.410000 558.500000 493.590000 ;
      RECT 516.500000 492.410000 549.500000 493.590000 ;
      RECT 507.500000 492.410000 508.500000 493.590000 ;
      RECT 466.500000 492.410000 499.500000 493.590000 ;
      RECT 457.500000 492.410000 458.500000 493.590000 ;
      RECT 416.500000 492.410000 449.500000 493.590000 ;
      RECT 407.500000 492.410000 408.500000 493.590000 ;
      RECT 386.500000 492.410000 399.500000 495.590000 ;
      RECT 372.500000 492.410000 373.500000 493.590000 ;
      RECT 357.500000 492.410000 358.500000 493.590000 ;
      RECT 316.500000 492.410000 349.500000 493.590000 ;
      RECT 307.500000 492.410000 308.500000 493.590000 ;
      RECT 266.500000 492.410000 299.500000 493.590000 ;
      RECT 257.500000 492.410000 258.500000 493.590000 ;
      RECT 216.500000 492.410000 249.500000 493.590000 ;
      RECT 207.500000 492.410000 208.500000 493.590000 ;
      RECT 166.500000 492.410000 199.500000 493.590000 ;
      RECT 157.500000 492.410000 158.500000 493.590000 ;
      RECT 116.500000 492.410000 149.500000 493.590000 ;
      RECT 107.500000 492.410000 108.500000 493.590000 ;
      RECT 66.500000 492.410000 99.500000 493.590000 ;
      RECT 57.500000 492.410000 58.500000 493.590000 ;
      RECT 29.500000 492.410000 49.500000 493.590000 ;
      RECT 15.500000 492.410000 16.500000 493.590000 ;
      RECT 0.000000 492.410000 2.500000 495.590000 ;
      RECT 1139.000000 491.590000 1158.500000 492.410000 ;
      RECT 716.500000 491.590000 739.000000 492.410000 ;
      RECT 666.500000 491.590000 708.500000 492.410000 ;
      RECT 616.500000 491.590000 658.500000 492.410000 ;
      RECT 566.500000 491.590000 608.500000 492.410000 ;
      RECT 516.500000 491.590000 558.500000 492.410000 ;
      RECT 466.500000 491.590000 508.500000 492.410000 ;
      RECT 416.500000 491.590000 458.500000 492.410000 ;
      RECT 372.500000 491.590000 408.500000 492.410000 ;
      RECT 316.500000 491.590000 358.500000 492.410000 ;
      RECT 266.500000 491.590000 308.500000 492.410000 ;
      RECT 216.500000 491.590000 258.500000 492.410000 ;
      RECT 166.500000 491.590000 208.500000 492.410000 ;
      RECT 116.500000 491.590000 158.500000 492.410000 ;
      RECT 66.500000 491.590000 108.500000 492.410000 ;
      RECT 29.500000 491.590000 58.500000 492.410000 ;
      RECT 0.000000 491.590000 16.500000 492.410000 ;
      RECT 1166.500000 490.410000 1186.000000 493.590000 ;
      RECT 1157.500000 490.410000 1158.500000 491.590000 ;
      RECT 716.500000 490.410000 723.500000 491.590000 ;
      RECT 707.500000 490.410000 708.500000 491.590000 ;
      RECT 666.500000 490.410000 699.500000 491.590000 ;
      RECT 657.500000 490.410000 658.500000 491.590000 ;
      RECT 616.500000 490.410000 649.500000 491.590000 ;
      RECT 607.500000 490.410000 608.500000 491.590000 ;
      RECT 566.500000 490.410000 599.500000 491.590000 ;
      RECT 557.500000 490.410000 558.500000 491.590000 ;
      RECT 516.500000 490.410000 549.500000 491.590000 ;
      RECT 507.500000 490.410000 508.500000 491.590000 ;
      RECT 466.500000 490.410000 499.500000 491.590000 ;
      RECT 457.500000 490.410000 458.500000 491.590000 ;
      RECT 416.500000 490.410000 449.500000 491.590000 ;
      RECT 407.500000 490.410000 408.500000 491.590000 ;
      RECT 372.500000 490.410000 399.500000 491.590000 ;
      RECT 357.500000 490.410000 358.500000 491.590000 ;
      RECT 316.500000 490.410000 349.500000 491.590000 ;
      RECT 307.500000 490.410000 308.500000 491.590000 ;
      RECT 266.500000 490.410000 299.500000 491.590000 ;
      RECT 257.500000 490.410000 258.500000 491.590000 ;
      RECT 216.500000 490.410000 249.500000 491.590000 ;
      RECT 207.500000 490.410000 208.500000 491.590000 ;
      RECT 166.500000 490.410000 199.500000 491.590000 ;
      RECT 157.500000 490.410000 158.500000 491.590000 ;
      RECT 116.500000 490.410000 149.500000 491.590000 ;
      RECT 107.500000 490.410000 108.500000 491.590000 ;
      RECT 66.500000 490.410000 99.500000 491.590000 ;
      RECT 57.500000 490.410000 58.500000 491.590000 ;
      RECT 29.500000 490.410000 49.500000 491.590000 ;
      RECT 15.500000 490.410000 16.500000 491.590000 ;
      RECT 1157.500000 489.590000 1186.000000 490.410000 ;
      RECT 707.500000 489.590000 723.500000 490.410000 ;
      RECT 657.500000 489.590000 699.500000 490.410000 ;
      RECT 607.500000 489.590000 649.500000 490.410000 ;
      RECT 557.500000 489.590000 599.500000 490.410000 ;
      RECT 507.500000 489.590000 549.500000 490.410000 ;
      RECT 457.500000 489.590000 499.500000 490.410000 ;
      RECT 407.500000 489.590000 449.500000 490.410000 ;
      RECT 357.500000 489.590000 399.500000 490.410000 ;
      RECT 307.500000 489.590000 349.500000 490.410000 ;
      RECT 257.500000 489.590000 299.500000 490.410000 ;
      RECT 207.500000 489.590000 249.500000 490.410000 ;
      RECT 157.500000 489.590000 199.500000 490.410000 ;
      RECT 107.500000 489.590000 149.500000 490.410000 ;
      RECT 57.500000 489.590000 99.500000 490.410000 ;
      RECT 15.500000 489.590000 49.500000 490.410000 ;
      RECT 1157.500000 488.410000 1158.500000 489.590000 ;
      RECT 1139.000000 488.410000 1149.500000 491.590000 ;
      RECT 736.500000 488.410000 739.000000 491.590000 ;
      RECT 722.500000 488.410000 723.500000 489.590000 ;
      RECT 707.500000 488.410000 708.500000 489.590000 ;
      RECT 666.500000 488.410000 699.500000 489.590000 ;
      RECT 657.500000 488.410000 658.500000 489.590000 ;
      RECT 616.500000 488.410000 649.500000 489.590000 ;
      RECT 607.500000 488.410000 608.500000 489.590000 ;
      RECT 566.500000 488.410000 599.500000 489.590000 ;
      RECT 557.500000 488.410000 558.500000 489.590000 ;
      RECT 516.500000 488.410000 549.500000 489.590000 ;
      RECT 507.500000 488.410000 508.500000 489.590000 ;
      RECT 466.500000 488.410000 499.500000 489.590000 ;
      RECT 457.500000 488.410000 458.500000 489.590000 ;
      RECT 416.500000 488.410000 449.500000 489.590000 ;
      RECT 407.500000 488.410000 408.500000 489.590000 ;
      RECT 372.500000 488.410000 399.500000 489.590000 ;
      RECT 357.500000 488.410000 359.500000 489.590000 ;
      RECT 316.500000 488.410000 349.500000 489.590000 ;
      RECT 307.500000 488.410000 308.500000 489.590000 ;
      RECT 266.500000 488.410000 299.500000 489.590000 ;
      RECT 257.500000 488.410000 258.500000 489.590000 ;
      RECT 216.500000 488.410000 249.500000 489.590000 ;
      RECT 207.500000 488.410000 208.500000 489.590000 ;
      RECT 166.500000 488.410000 199.500000 489.590000 ;
      RECT 157.500000 488.410000 158.500000 489.590000 ;
      RECT 116.500000 488.410000 149.500000 489.590000 ;
      RECT 107.500000 488.410000 108.500000 489.590000 ;
      RECT 66.500000 488.410000 99.500000 489.590000 ;
      RECT 57.500000 488.410000 58.500000 489.590000 ;
      RECT 29.500000 488.410000 49.500000 489.590000 ;
      RECT 15.500000 488.410000 16.500000 489.590000 ;
      RECT 0.000000 488.410000 2.500000 491.590000 ;
      RECT 1139.000000 487.590000 1158.500000 488.410000 ;
      RECT 722.500000 487.590000 739.000000 488.410000 ;
      RECT 666.500000 487.590000 708.500000 488.410000 ;
      RECT 616.500000 487.590000 658.500000 488.410000 ;
      RECT 566.500000 487.590000 608.500000 488.410000 ;
      RECT 516.500000 487.590000 558.500000 488.410000 ;
      RECT 466.500000 487.590000 508.500000 488.410000 ;
      RECT 416.500000 487.590000 458.500000 488.410000 ;
      RECT 372.500000 487.590000 408.500000 488.410000 ;
      RECT 316.500000 487.590000 359.500000 488.410000 ;
      RECT 266.500000 487.590000 308.500000 488.410000 ;
      RECT 216.500000 487.590000 258.500000 488.410000 ;
      RECT 166.500000 487.590000 208.500000 488.410000 ;
      RECT 116.500000 487.590000 158.500000 488.410000 ;
      RECT 66.500000 487.590000 108.500000 488.410000 ;
      RECT 29.500000 487.590000 58.500000 488.410000 ;
      RECT 0.000000 487.590000 16.500000 488.410000 ;
      RECT 1166.500000 486.410000 1186.000000 489.590000 ;
      RECT 1157.500000 486.410000 1158.500000 487.590000 ;
      RECT 722.500000 486.410000 723.500000 487.590000 ;
      RECT 707.500000 486.410000 708.500000 487.590000 ;
      RECT 666.500000 486.410000 699.500000 487.590000 ;
      RECT 657.500000 486.410000 658.500000 487.590000 ;
      RECT 616.500000 486.410000 649.500000 487.590000 ;
      RECT 607.500000 486.410000 608.500000 487.590000 ;
      RECT 566.500000 486.410000 599.500000 487.590000 ;
      RECT 557.500000 486.410000 558.500000 487.590000 ;
      RECT 516.500000 486.410000 549.500000 487.590000 ;
      RECT 507.500000 486.410000 508.500000 487.590000 ;
      RECT 466.500000 486.410000 499.500000 487.590000 ;
      RECT 457.500000 486.410000 458.500000 487.590000 ;
      RECT 416.500000 486.410000 449.500000 487.590000 ;
      RECT 407.500000 486.410000 408.500000 487.590000 ;
      RECT 372.500000 486.410000 399.500000 487.590000 ;
      RECT 357.500000 486.410000 359.500000 487.590000 ;
      RECT 316.500000 486.410000 349.500000 487.590000 ;
      RECT 307.500000 486.410000 308.500000 487.590000 ;
      RECT 266.500000 486.410000 299.500000 487.590000 ;
      RECT 257.500000 486.410000 258.500000 487.590000 ;
      RECT 216.500000 486.410000 249.500000 487.590000 ;
      RECT 207.500000 486.410000 208.500000 487.590000 ;
      RECT 166.500000 486.410000 199.500000 487.590000 ;
      RECT 157.500000 486.410000 158.500000 487.590000 ;
      RECT 116.500000 486.410000 149.500000 487.590000 ;
      RECT 107.500000 486.410000 108.500000 487.590000 ;
      RECT 66.500000 486.410000 99.500000 487.590000 ;
      RECT 57.500000 486.410000 58.500000 487.590000 ;
      RECT 29.500000 486.410000 49.500000 487.590000 ;
      RECT 15.500000 486.410000 16.500000 487.590000 ;
      RECT 1157.500000 485.590000 1186.000000 486.410000 ;
      RECT 707.500000 485.590000 723.500000 486.410000 ;
      RECT 657.500000 485.590000 699.500000 486.410000 ;
      RECT 607.500000 485.590000 649.500000 486.410000 ;
      RECT 557.500000 485.590000 599.500000 486.410000 ;
      RECT 507.500000 485.590000 549.500000 486.410000 ;
      RECT 457.500000 485.590000 499.500000 486.410000 ;
      RECT 407.500000 485.590000 449.500000 486.410000 ;
      RECT 357.500000 485.590000 399.500000 486.410000 ;
      RECT 307.500000 485.590000 349.500000 486.410000 ;
      RECT 257.500000 485.590000 299.500000 486.410000 ;
      RECT 207.500000 485.590000 249.500000 486.410000 ;
      RECT 157.500000 485.590000 199.500000 486.410000 ;
      RECT 107.500000 485.590000 149.500000 486.410000 ;
      RECT 57.500000 485.590000 99.500000 486.410000 ;
      RECT 15.500000 485.590000 49.500000 486.410000 ;
      RECT 1157.500000 484.410000 1158.500000 485.590000 ;
      RECT 1139.000000 484.410000 1149.500000 487.590000 ;
      RECT 736.500000 484.410000 739.000000 487.590000 ;
      RECT 722.500000 484.410000 723.500000 485.590000 ;
      RECT 707.500000 484.410000 708.500000 485.590000 ;
      RECT 666.500000 484.410000 699.500000 485.590000 ;
      RECT 657.500000 484.410000 658.500000 485.590000 ;
      RECT 616.500000 484.410000 649.500000 485.590000 ;
      RECT 607.500000 484.410000 608.500000 485.590000 ;
      RECT 566.500000 484.410000 599.500000 485.590000 ;
      RECT 557.500000 484.410000 558.500000 485.590000 ;
      RECT 516.500000 484.410000 549.500000 485.590000 ;
      RECT 507.500000 484.410000 508.500000 485.590000 ;
      RECT 466.500000 484.410000 499.500000 485.590000 ;
      RECT 457.500000 484.410000 458.500000 485.590000 ;
      RECT 416.500000 484.410000 449.500000 485.590000 ;
      RECT 407.500000 484.410000 408.500000 485.590000 ;
      RECT 372.500000 484.410000 399.500000 485.590000 ;
      RECT 357.500000 484.410000 359.500000 485.590000 ;
      RECT 316.500000 484.410000 349.500000 485.590000 ;
      RECT 307.500000 484.410000 308.500000 485.590000 ;
      RECT 266.500000 484.410000 299.500000 485.590000 ;
      RECT 257.500000 484.410000 258.500000 485.590000 ;
      RECT 216.500000 484.410000 249.500000 485.590000 ;
      RECT 207.500000 484.410000 208.500000 485.590000 ;
      RECT 166.500000 484.410000 199.500000 485.590000 ;
      RECT 157.500000 484.410000 158.500000 485.590000 ;
      RECT 116.500000 484.410000 149.500000 485.590000 ;
      RECT 107.500000 484.410000 108.500000 485.590000 ;
      RECT 66.500000 484.410000 99.500000 485.590000 ;
      RECT 57.500000 484.410000 58.500000 485.590000 ;
      RECT 29.500000 484.410000 49.500000 485.590000 ;
      RECT 15.500000 484.410000 16.500000 485.590000 ;
      RECT 0.000000 484.410000 2.500000 487.590000 ;
      RECT 1139.000000 483.590000 1158.500000 484.410000 ;
      RECT 722.500000 483.590000 739.000000 484.410000 ;
      RECT 666.500000 483.590000 708.500000 484.410000 ;
      RECT 616.500000 483.590000 658.500000 484.410000 ;
      RECT 566.500000 483.590000 608.500000 484.410000 ;
      RECT 516.500000 483.590000 558.500000 484.410000 ;
      RECT 466.500000 483.590000 508.500000 484.410000 ;
      RECT 416.500000 483.590000 458.500000 484.410000 ;
      RECT 372.500000 483.590000 408.500000 484.410000 ;
      RECT 316.500000 483.590000 359.500000 484.410000 ;
      RECT 266.500000 483.590000 308.500000 484.410000 ;
      RECT 216.500000 483.590000 258.500000 484.410000 ;
      RECT 166.500000 483.590000 208.500000 484.410000 ;
      RECT 116.500000 483.590000 158.500000 484.410000 ;
      RECT 66.500000 483.590000 108.500000 484.410000 ;
      RECT 29.500000 483.590000 58.500000 484.410000 ;
      RECT 0.000000 483.590000 16.500000 484.410000 ;
      RECT 1166.500000 482.410000 1186.000000 485.590000 ;
      RECT 1157.500000 482.410000 1158.500000 483.590000 ;
      RECT 722.500000 482.410000 723.500000 483.590000 ;
      RECT 707.500000 482.410000 708.500000 483.590000 ;
      RECT 666.500000 482.410000 699.500000 483.590000 ;
      RECT 657.500000 482.410000 658.500000 483.590000 ;
      RECT 616.500000 482.410000 649.500000 483.590000 ;
      RECT 607.500000 482.410000 608.500000 483.590000 ;
      RECT 566.500000 482.410000 599.500000 483.590000 ;
      RECT 557.500000 482.410000 558.500000 483.590000 ;
      RECT 516.500000 482.410000 549.500000 483.590000 ;
      RECT 507.500000 482.410000 508.500000 483.590000 ;
      RECT 466.500000 482.410000 499.500000 483.590000 ;
      RECT 457.500000 482.410000 458.500000 483.590000 ;
      RECT 416.500000 482.410000 449.500000 483.590000 ;
      RECT 407.500000 482.410000 408.500000 483.590000 ;
      RECT 372.500000 482.410000 399.500000 483.590000 ;
      RECT 357.500000 482.410000 359.500000 483.590000 ;
      RECT 316.500000 482.410000 349.500000 483.590000 ;
      RECT 307.500000 482.410000 308.500000 483.590000 ;
      RECT 266.500000 482.410000 299.500000 483.590000 ;
      RECT 257.500000 482.410000 258.500000 483.590000 ;
      RECT 216.500000 482.410000 249.500000 483.590000 ;
      RECT 207.500000 482.410000 208.500000 483.590000 ;
      RECT 166.500000 482.410000 199.500000 483.590000 ;
      RECT 157.500000 482.410000 158.500000 483.590000 ;
      RECT 116.500000 482.410000 149.500000 483.590000 ;
      RECT 107.500000 482.410000 108.500000 483.590000 ;
      RECT 66.500000 482.410000 99.500000 483.590000 ;
      RECT 57.500000 482.410000 58.500000 483.590000 ;
      RECT 29.500000 482.410000 49.500000 483.590000 ;
      RECT 15.500000 482.410000 16.500000 483.590000 ;
      RECT 1157.500000 481.590000 1186.000000 482.410000 ;
      RECT 707.500000 481.590000 723.500000 482.410000 ;
      RECT 657.500000 481.590000 699.500000 482.410000 ;
      RECT 607.500000 481.590000 649.500000 482.410000 ;
      RECT 557.500000 481.590000 599.500000 482.410000 ;
      RECT 507.500000 481.590000 549.500000 482.410000 ;
      RECT 457.500000 481.590000 499.500000 482.410000 ;
      RECT 407.500000 481.590000 449.500000 482.410000 ;
      RECT 357.500000 481.590000 399.500000 482.410000 ;
      RECT 307.500000 481.590000 349.500000 482.410000 ;
      RECT 257.500000 481.590000 299.500000 482.410000 ;
      RECT 207.500000 481.590000 249.500000 482.410000 ;
      RECT 157.500000 481.590000 199.500000 482.410000 ;
      RECT 107.500000 481.590000 149.500000 482.410000 ;
      RECT 57.500000 481.590000 99.500000 482.410000 ;
      RECT 15.500000 481.590000 49.500000 482.410000 ;
      RECT 1157.500000 480.410000 1158.500000 481.590000 ;
      RECT 1139.000000 480.410000 1149.500000 483.590000 ;
      RECT 736.500000 480.410000 739.000000 483.590000 ;
      RECT 722.500000 480.410000 723.500000 481.590000 ;
      RECT 707.500000 480.410000 708.500000 481.590000 ;
      RECT 666.500000 480.410000 699.500000 481.590000 ;
      RECT 657.500000 480.410000 658.500000 481.590000 ;
      RECT 616.500000 480.410000 649.500000 481.590000 ;
      RECT 607.500000 480.410000 608.500000 481.590000 ;
      RECT 566.500000 480.410000 599.500000 481.590000 ;
      RECT 557.500000 480.410000 558.500000 481.590000 ;
      RECT 516.500000 480.410000 549.500000 481.590000 ;
      RECT 507.500000 480.410000 508.500000 481.590000 ;
      RECT 466.500000 480.410000 499.500000 481.590000 ;
      RECT 457.500000 480.410000 458.500000 481.590000 ;
      RECT 416.500000 480.410000 449.500000 481.590000 ;
      RECT 407.500000 480.410000 408.500000 481.590000 ;
      RECT 372.500000 480.410000 399.500000 481.590000 ;
      RECT 357.500000 480.410000 359.500000 481.590000 ;
      RECT 316.500000 480.410000 349.500000 481.590000 ;
      RECT 307.500000 480.410000 308.500000 481.590000 ;
      RECT 266.500000 480.410000 299.500000 481.590000 ;
      RECT 257.500000 480.410000 258.500000 481.590000 ;
      RECT 216.500000 480.410000 249.500000 481.590000 ;
      RECT 207.500000 480.410000 208.500000 481.590000 ;
      RECT 166.500000 480.410000 199.500000 481.590000 ;
      RECT 157.500000 480.410000 158.500000 481.590000 ;
      RECT 116.500000 480.410000 149.500000 481.590000 ;
      RECT 107.500000 480.410000 108.500000 481.590000 ;
      RECT 66.500000 480.410000 99.500000 481.590000 ;
      RECT 57.500000 480.410000 58.500000 481.590000 ;
      RECT 29.500000 480.410000 49.500000 481.590000 ;
      RECT 15.500000 480.410000 16.500000 481.590000 ;
      RECT 0.000000 480.410000 2.500000 483.590000 ;
      RECT 1139.000000 479.590000 1158.500000 480.410000 ;
      RECT 722.500000 479.590000 739.000000 480.410000 ;
      RECT 666.500000 479.590000 708.500000 480.410000 ;
      RECT 616.500000 479.590000 658.500000 480.410000 ;
      RECT 566.500000 479.590000 608.500000 480.410000 ;
      RECT 516.500000 479.590000 558.500000 480.410000 ;
      RECT 466.500000 479.590000 508.500000 480.410000 ;
      RECT 416.500000 479.590000 458.500000 480.410000 ;
      RECT 372.500000 479.590000 408.500000 480.410000 ;
      RECT 316.500000 479.590000 359.500000 480.410000 ;
      RECT 266.500000 479.590000 308.500000 480.410000 ;
      RECT 216.500000 479.590000 258.500000 480.410000 ;
      RECT 166.500000 479.590000 208.500000 480.410000 ;
      RECT 116.500000 479.590000 158.500000 480.410000 ;
      RECT 66.500000 479.590000 108.500000 480.410000 ;
      RECT 29.500000 479.590000 58.500000 480.410000 ;
      RECT 0.000000 479.590000 16.500000 480.410000 ;
      RECT 1166.500000 478.410000 1186.000000 481.590000 ;
      RECT 1157.500000 478.410000 1158.500000 479.590000 ;
      RECT 722.500000 478.410000 723.500000 479.590000 ;
      RECT 707.500000 478.410000 708.500000 479.590000 ;
      RECT 666.500000 478.410000 699.500000 479.590000 ;
      RECT 657.500000 478.410000 658.500000 479.590000 ;
      RECT 616.500000 478.410000 649.500000 479.590000 ;
      RECT 607.500000 478.410000 608.500000 479.590000 ;
      RECT 566.500000 478.410000 599.500000 479.590000 ;
      RECT 557.500000 478.410000 558.500000 479.590000 ;
      RECT 516.500000 478.410000 549.500000 479.590000 ;
      RECT 507.500000 478.410000 508.500000 479.590000 ;
      RECT 466.500000 478.410000 499.500000 479.590000 ;
      RECT 457.500000 478.410000 458.500000 479.590000 ;
      RECT 416.500000 478.410000 449.500000 479.590000 ;
      RECT 407.500000 478.410000 408.500000 479.590000 ;
      RECT 372.500000 478.410000 399.500000 479.590000 ;
      RECT 357.500000 478.410000 359.500000 479.590000 ;
      RECT 316.500000 478.410000 349.500000 479.590000 ;
      RECT 307.500000 478.410000 308.500000 479.590000 ;
      RECT 266.500000 478.410000 299.500000 479.590000 ;
      RECT 257.500000 478.410000 258.500000 479.590000 ;
      RECT 216.500000 478.410000 249.500000 479.590000 ;
      RECT 207.500000 478.410000 208.500000 479.590000 ;
      RECT 166.500000 478.410000 199.500000 479.590000 ;
      RECT 157.500000 478.410000 158.500000 479.590000 ;
      RECT 116.500000 478.410000 149.500000 479.590000 ;
      RECT 107.500000 478.410000 108.500000 479.590000 ;
      RECT 66.500000 478.410000 99.500000 479.590000 ;
      RECT 57.500000 478.410000 58.500000 479.590000 ;
      RECT 29.500000 478.410000 49.500000 479.590000 ;
      RECT 15.500000 478.410000 16.500000 479.590000 ;
      RECT 1157.500000 477.590000 1186.000000 478.410000 ;
      RECT 707.500000 477.590000 723.500000 478.410000 ;
      RECT 657.500000 477.590000 699.500000 478.410000 ;
      RECT 607.500000 477.590000 649.500000 478.410000 ;
      RECT 557.500000 477.590000 599.500000 478.410000 ;
      RECT 507.500000 477.590000 549.500000 478.410000 ;
      RECT 457.500000 477.590000 499.500000 478.410000 ;
      RECT 407.500000 477.590000 449.500000 478.410000 ;
      RECT 357.500000 477.590000 399.500000 478.410000 ;
      RECT 307.500000 477.590000 349.500000 478.410000 ;
      RECT 257.500000 477.590000 299.500000 478.410000 ;
      RECT 207.500000 477.590000 249.500000 478.410000 ;
      RECT 157.500000 477.590000 199.500000 478.410000 ;
      RECT 107.500000 477.590000 149.500000 478.410000 ;
      RECT 57.500000 477.590000 99.500000 478.410000 ;
      RECT 15.500000 477.590000 49.500000 478.410000 ;
      RECT 1157.500000 476.410000 1158.500000 477.590000 ;
      RECT 1139.000000 476.410000 1149.500000 479.590000 ;
      RECT 736.500000 476.410000 739.000000 479.590000 ;
      RECT 722.500000 476.410000 723.500000 477.590000 ;
      RECT 707.500000 476.410000 708.500000 477.590000 ;
      RECT 666.500000 476.410000 699.500000 477.590000 ;
      RECT 657.500000 476.410000 658.500000 477.590000 ;
      RECT 616.500000 476.410000 649.500000 477.590000 ;
      RECT 607.500000 476.410000 608.500000 477.590000 ;
      RECT 566.500000 476.410000 599.500000 477.590000 ;
      RECT 557.500000 476.410000 558.500000 477.590000 ;
      RECT 516.500000 476.410000 549.500000 477.590000 ;
      RECT 507.500000 476.410000 508.500000 477.590000 ;
      RECT 466.500000 476.410000 499.500000 477.590000 ;
      RECT 457.500000 476.410000 458.500000 477.590000 ;
      RECT 416.500000 476.410000 449.500000 477.590000 ;
      RECT 407.500000 476.410000 408.500000 477.590000 ;
      RECT 370.000000 476.410000 399.500000 477.590000 ;
      RECT 357.500000 476.410000 362.000000 477.590000 ;
      RECT 316.500000 476.410000 349.500000 477.590000 ;
      RECT 307.500000 476.410000 308.500000 477.590000 ;
      RECT 266.500000 476.410000 299.500000 477.590000 ;
      RECT 257.500000 476.410000 258.500000 477.590000 ;
      RECT 216.500000 476.410000 249.500000 477.590000 ;
      RECT 207.500000 476.410000 208.500000 477.590000 ;
      RECT 166.500000 476.410000 199.500000 477.590000 ;
      RECT 157.500000 476.410000 158.500000 477.590000 ;
      RECT 116.500000 476.410000 149.500000 477.590000 ;
      RECT 107.500000 476.410000 108.500000 477.590000 ;
      RECT 66.500000 476.410000 99.500000 477.590000 ;
      RECT 57.500000 476.410000 58.500000 477.590000 ;
      RECT 29.500000 476.410000 49.500000 477.590000 ;
      RECT 15.500000 476.410000 16.500000 477.590000 ;
      RECT 0.000000 476.410000 2.500000 479.590000 ;
      RECT 1139.000000 475.590000 1158.500000 476.410000 ;
      RECT 722.500000 475.590000 739.000000 476.410000 ;
      RECT 666.500000 475.590000 708.500000 476.410000 ;
      RECT 616.500000 475.590000 658.500000 476.410000 ;
      RECT 566.500000 475.590000 608.500000 476.410000 ;
      RECT 516.500000 475.590000 558.500000 476.410000 ;
      RECT 466.500000 475.590000 508.500000 476.410000 ;
      RECT 416.500000 475.590000 458.500000 476.410000 ;
      RECT 370.000000 475.590000 408.500000 476.410000 ;
      RECT 316.500000 475.590000 362.000000 476.410000 ;
      RECT 266.500000 475.590000 308.500000 476.410000 ;
      RECT 216.500000 475.590000 258.500000 476.410000 ;
      RECT 166.500000 475.590000 208.500000 476.410000 ;
      RECT 116.500000 475.590000 158.500000 476.410000 ;
      RECT 66.500000 475.590000 108.500000 476.410000 ;
      RECT 29.500000 475.590000 58.500000 476.410000 ;
      RECT 0.000000 475.590000 16.500000 476.410000 ;
      RECT 1166.500000 474.410000 1186.000000 477.590000 ;
      RECT 1157.500000 474.410000 1158.500000 475.590000 ;
      RECT 722.500000 474.410000 723.500000 475.590000 ;
      RECT 707.500000 474.410000 708.500000 475.590000 ;
      RECT 666.500000 474.410000 699.500000 475.590000 ;
      RECT 657.500000 474.410000 658.500000 475.590000 ;
      RECT 616.500000 474.410000 649.500000 475.590000 ;
      RECT 607.500000 474.410000 608.500000 475.590000 ;
      RECT 566.500000 474.410000 599.500000 475.590000 ;
      RECT 557.500000 474.410000 558.500000 475.590000 ;
      RECT 516.500000 474.410000 549.500000 475.590000 ;
      RECT 507.500000 474.410000 508.500000 475.590000 ;
      RECT 466.500000 474.410000 499.500000 475.590000 ;
      RECT 457.500000 474.410000 458.500000 475.590000 ;
      RECT 416.500000 474.410000 449.500000 475.590000 ;
      RECT 407.500000 474.410000 408.500000 475.590000 ;
      RECT 370.000000 474.410000 399.500000 475.590000 ;
      RECT 357.500000 474.410000 362.000000 475.590000 ;
      RECT 316.500000 474.410000 349.500000 475.590000 ;
      RECT 307.500000 474.410000 308.500000 475.590000 ;
      RECT 266.500000 474.410000 299.500000 475.590000 ;
      RECT 257.500000 474.410000 258.500000 475.590000 ;
      RECT 216.500000 474.410000 249.500000 475.590000 ;
      RECT 207.500000 474.410000 208.500000 475.590000 ;
      RECT 166.500000 474.410000 199.500000 475.590000 ;
      RECT 157.500000 474.410000 158.500000 475.590000 ;
      RECT 116.500000 474.410000 149.500000 475.590000 ;
      RECT 107.500000 474.410000 108.500000 475.590000 ;
      RECT 66.500000 474.410000 99.500000 475.590000 ;
      RECT 57.500000 474.410000 58.500000 475.590000 ;
      RECT 29.500000 474.410000 49.500000 475.590000 ;
      RECT 15.500000 474.410000 16.500000 475.590000 ;
      RECT 1157.500000 473.590000 1186.000000 474.410000 ;
      RECT 707.500000 473.590000 723.500000 474.410000 ;
      RECT 657.500000 473.590000 699.500000 474.410000 ;
      RECT 607.500000 473.590000 649.500000 474.410000 ;
      RECT 557.500000 473.590000 599.500000 474.410000 ;
      RECT 507.500000 473.590000 549.500000 474.410000 ;
      RECT 457.500000 473.590000 499.500000 474.410000 ;
      RECT 407.500000 473.590000 449.500000 474.410000 ;
      RECT 357.500000 473.590000 399.500000 474.410000 ;
      RECT 307.500000 473.590000 349.500000 474.410000 ;
      RECT 257.500000 473.590000 299.500000 474.410000 ;
      RECT 207.500000 473.590000 249.500000 474.410000 ;
      RECT 157.500000 473.590000 199.500000 474.410000 ;
      RECT 107.500000 473.590000 149.500000 474.410000 ;
      RECT 57.500000 473.590000 99.500000 474.410000 ;
      RECT 15.500000 473.590000 49.500000 474.410000 ;
      RECT 1157.500000 472.410000 1158.500000 473.590000 ;
      RECT 1139.000000 472.410000 1149.500000 475.590000 ;
      RECT 736.500000 472.410000 739.000000 475.590000 ;
      RECT 722.500000 472.410000 723.500000 473.590000 ;
      RECT 707.500000 472.410000 708.500000 473.590000 ;
      RECT 666.500000 472.410000 699.500000 473.590000 ;
      RECT 657.500000 472.410000 658.500000 473.590000 ;
      RECT 616.500000 472.410000 649.500000 473.590000 ;
      RECT 607.500000 472.410000 608.500000 473.590000 ;
      RECT 566.500000 472.410000 599.500000 473.590000 ;
      RECT 557.500000 472.410000 558.500000 473.590000 ;
      RECT 516.500000 472.410000 549.500000 473.590000 ;
      RECT 507.500000 472.410000 508.500000 473.590000 ;
      RECT 466.500000 472.410000 499.500000 473.590000 ;
      RECT 457.500000 472.410000 458.500000 473.590000 ;
      RECT 416.500000 472.410000 449.500000 473.590000 ;
      RECT 407.500000 472.410000 408.500000 473.590000 ;
      RECT 370.000000 472.410000 399.500000 473.590000 ;
      RECT 357.500000 472.410000 358.500000 473.590000 ;
      RECT 316.500000 472.410000 349.500000 473.590000 ;
      RECT 307.500000 472.410000 308.500000 473.590000 ;
      RECT 266.500000 472.410000 299.500000 473.590000 ;
      RECT 257.500000 472.410000 258.500000 473.590000 ;
      RECT 216.500000 472.410000 249.500000 473.590000 ;
      RECT 207.500000 472.410000 208.500000 473.590000 ;
      RECT 166.500000 472.410000 199.500000 473.590000 ;
      RECT 157.500000 472.410000 158.500000 473.590000 ;
      RECT 116.500000 472.410000 149.500000 473.590000 ;
      RECT 107.500000 472.410000 108.500000 473.590000 ;
      RECT 66.500000 472.410000 99.500000 473.590000 ;
      RECT 57.500000 472.410000 58.500000 473.590000 ;
      RECT 29.500000 472.410000 49.500000 473.590000 ;
      RECT 15.500000 472.410000 16.500000 473.590000 ;
      RECT 0.000000 472.410000 2.500000 475.590000 ;
      RECT 1139.000000 471.590000 1158.500000 472.410000 ;
      RECT 722.500000 471.590000 739.000000 472.410000 ;
      RECT 666.500000 471.590000 708.500000 472.410000 ;
      RECT 616.500000 471.590000 658.500000 472.410000 ;
      RECT 566.500000 471.590000 608.500000 472.410000 ;
      RECT 516.500000 471.590000 558.500000 472.410000 ;
      RECT 466.500000 471.590000 508.500000 472.410000 ;
      RECT 416.500000 471.590000 458.500000 472.410000 ;
      RECT 370.000000 471.590000 408.500000 472.410000 ;
      RECT 316.500000 471.590000 358.500000 472.410000 ;
      RECT 266.500000 471.590000 308.500000 472.410000 ;
      RECT 216.500000 471.590000 258.500000 472.410000 ;
      RECT 166.500000 471.590000 208.500000 472.410000 ;
      RECT 116.500000 471.590000 158.500000 472.410000 ;
      RECT 66.500000 471.590000 108.500000 472.410000 ;
      RECT 29.500000 471.590000 58.500000 472.410000 ;
      RECT 0.000000 471.590000 16.500000 472.410000 ;
      RECT 1166.500000 470.410000 1186.000000 473.590000 ;
      RECT 1157.500000 470.410000 1158.500000 471.590000 ;
      RECT 722.500000 470.410000 723.500000 471.590000 ;
      RECT 707.500000 470.410000 708.500000 471.590000 ;
      RECT 666.500000 470.410000 699.500000 471.590000 ;
      RECT 657.500000 470.410000 658.500000 471.590000 ;
      RECT 616.500000 470.410000 649.500000 471.590000 ;
      RECT 607.500000 470.410000 608.500000 471.590000 ;
      RECT 566.500000 470.410000 599.500000 471.590000 ;
      RECT 557.500000 470.410000 558.500000 471.590000 ;
      RECT 516.500000 470.410000 549.500000 471.590000 ;
      RECT 507.500000 470.410000 508.500000 471.590000 ;
      RECT 466.500000 470.410000 499.500000 471.590000 ;
      RECT 457.500000 470.410000 458.500000 471.590000 ;
      RECT 416.500000 470.410000 449.500000 471.590000 ;
      RECT 407.500000 470.410000 408.500000 471.590000 ;
      RECT 370.000000 470.410000 399.500000 471.590000 ;
      RECT 357.500000 470.410000 358.500000 471.590000 ;
      RECT 316.500000 470.410000 349.500000 471.590000 ;
      RECT 307.500000 470.410000 308.500000 471.590000 ;
      RECT 266.500000 470.410000 299.500000 471.590000 ;
      RECT 257.500000 470.410000 258.500000 471.590000 ;
      RECT 216.500000 470.410000 249.500000 471.590000 ;
      RECT 207.500000 470.410000 208.500000 471.590000 ;
      RECT 166.500000 470.410000 199.500000 471.590000 ;
      RECT 157.500000 470.410000 158.500000 471.590000 ;
      RECT 116.500000 470.410000 149.500000 471.590000 ;
      RECT 107.500000 470.410000 108.500000 471.590000 ;
      RECT 66.500000 470.410000 99.500000 471.590000 ;
      RECT 57.500000 470.410000 58.500000 471.590000 ;
      RECT 29.500000 470.410000 49.500000 471.590000 ;
      RECT 15.500000 470.410000 16.500000 471.590000 ;
      RECT 1157.500000 469.590000 1186.000000 470.410000 ;
      RECT 707.500000 469.590000 723.500000 470.410000 ;
      RECT 657.500000 469.590000 699.500000 470.410000 ;
      RECT 607.500000 469.590000 649.500000 470.410000 ;
      RECT 557.500000 469.590000 599.500000 470.410000 ;
      RECT 507.500000 469.590000 549.500000 470.410000 ;
      RECT 457.500000 469.590000 499.500000 470.410000 ;
      RECT 407.500000 469.590000 449.500000 470.410000 ;
      RECT 357.500000 469.590000 399.500000 470.410000 ;
      RECT 307.500000 469.590000 349.500000 470.410000 ;
      RECT 257.500000 469.590000 299.500000 470.410000 ;
      RECT 207.500000 469.590000 249.500000 470.410000 ;
      RECT 157.500000 469.590000 199.500000 470.410000 ;
      RECT 107.500000 469.590000 149.500000 470.410000 ;
      RECT 57.500000 469.590000 99.500000 470.410000 ;
      RECT 15.500000 469.590000 49.500000 470.410000 ;
      RECT 1157.500000 468.410000 1158.500000 469.590000 ;
      RECT 1139.000000 468.410000 1149.500000 471.590000 ;
      RECT 736.500000 468.410000 739.000000 471.590000 ;
      RECT 722.500000 468.410000 723.500000 469.590000 ;
      RECT 707.500000 468.410000 708.500000 469.590000 ;
      RECT 666.500000 468.410000 699.500000 469.590000 ;
      RECT 657.500000 468.410000 658.500000 469.590000 ;
      RECT 616.500000 468.410000 649.500000 469.590000 ;
      RECT 607.500000 468.410000 608.500000 469.590000 ;
      RECT 566.500000 468.410000 599.500000 469.590000 ;
      RECT 557.500000 468.410000 558.500000 469.590000 ;
      RECT 516.500000 468.410000 549.500000 469.590000 ;
      RECT 507.500000 468.410000 508.500000 469.590000 ;
      RECT 466.500000 468.410000 499.500000 469.590000 ;
      RECT 457.500000 468.410000 458.500000 469.590000 ;
      RECT 416.500000 468.410000 449.500000 469.590000 ;
      RECT 407.500000 468.410000 408.500000 469.590000 ;
      RECT 366.500000 468.410000 399.500000 469.590000 ;
      RECT 357.500000 468.410000 358.500000 469.590000 ;
      RECT 316.500000 468.410000 349.500000 469.590000 ;
      RECT 307.500000 468.410000 308.500000 469.590000 ;
      RECT 266.500000 468.410000 299.500000 469.590000 ;
      RECT 257.500000 468.410000 258.500000 469.590000 ;
      RECT 216.500000 468.410000 249.500000 469.590000 ;
      RECT 207.500000 468.410000 208.500000 469.590000 ;
      RECT 166.500000 468.410000 199.500000 469.590000 ;
      RECT 157.500000 468.410000 158.500000 469.590000 ;
      RECT 116.500000 468.410000 149.500000 469.590000 ;
      RECT 107.500000 468.410000 108.500000 469.590000 ;
      RECT 66.500000 468.410000 99.500000 469.590000 ;
      RECT 57.500000 468.410000 58.500000 469.590000 ;
      RECT 29.500000 468.410000 49.500000 469.590000 ;
      RECT 15.500000 468.410000 16.500000 469.590000 ;
      RECT 0.000000 468.410000 2.500000 471.590000 ;
      RECT 1139.000000 467.590000 1158.500000 468.410000 ;
      RECT 722.500000 467.590000 739.000000 468.410000 ;
      RECT 666.500000 467.590000 708.500000 468.410000 ;
      RECT 616.500000 467.590000 658.500000 468.410000 ;
      RECT 566.500000 467.590000 608.500000 468.410000 ;
      RECT 516.500000 467.590000 558.500000 468.410000 ;
      RECT 466.500000 467.590000 508.500000 468.410000 ;
      RECT 416.500000 467.590000 458.500000 468.410000 ;
      RECT 366.500000 467.590000 408.500000 468.410000 ;
      RECT 316.500000 467.590000 358.500000 468.410000 ;
      RECT 266.500000 467.590000 308.500000 468.410000 ;
      RECT 216.500000 467.590000 258.500000 468.410000 ;
      RECT 166.500000 467.590000 208.500000 468.410000 ;
      RECT 116.500000 467.590000 158.500000 468.410000 ;
      RECT 66.500000 467.590000 108.500000 468.410000 ;
      RECT 29.500000 467.590000 58.500000 468.410000 ;
      RECT 0.000000 467.590000 16.500000 468.410000 ;
      RECT 1166.500000 466.410000 1186.000000 469.590000 ;
      RECT 1157.500000 466.410000 1158.500000 467.590000 ;
      RECT 722.500000 466.410000 723.500000 467.590000 ;
      RECT 707.500000 466.410000 708.500000 467.590000 ;
      RECT 666.500000 466.410000 699.500000 467.590000 ;
      RECT 657.500000 466.410000 658.500000 467.590000 ;
      RECT 616.500000 466.410000 649.500000 467.590000 ;
      RECT 607.500000 466.410000 608.500000 467.590000 ;
      RECT 566.500000 466.410000 599.500000 467.590000 ;
      RECT 557.500000 466.410000 558.500000 467.590000 ;
      RECT 516.500000 466.410000 549.500000 467.590000 ;
      RECT 507.500000 466.410000 508.500000 467.590000 ;
      RECT 466.500000 466.410000 499.500000 467.590000 ;
      RECT 457.500000 466.410000 458.500000 467.590000 ;
      RECT 416.500000 466.410000 449.500000 467.590000 ;
      RECT 407.500000 466.410000 408.500000 467.590000 ;
      RECT 366.500000 466.410000 399.500000 467.590000 ;
      RECT 357.500000 466.410000 358.500000 467.590000 ;
      RECT 316.500000 466.410000 349.500000 467.590000 ;
      RECT 307.500000 466.410000 308.500000 467.590000 ;
      RECT 266.500000 466.410000 299.500000 467.590000 ;
      RECT 257.500000 466.410000 258.500000 467.590000 ;
      RECT 216.500000 466.410000 249.500000 467.590000 ;
      RECT 207.500000 466.410000 208.500000 467.590000 ;
      RECT 166.500000 466.410000 199.500000 467.590000 ;
      RECT 157.500000 466.410000 158.500000 467.590000 ;
      RECT 116.500000 466.410000 149.500000 467.590000 ;
      RECT 107.500000 466.410000 108.500000 467.590000 ;
      RECT 66.500000 466.410000 99.500000 467.590000 ;
      RECT 57.500000 466.410000 58.500000 467.590000 ;
      RECT 29.500000 466.410000 49.500000 467.590000 ;
      RECT 15.500000 466.410000 16.500000 467.590000 ;
      RECT 1157.500000 465.590000 1186.000000 466.410000 ;
      RECT 707.500000 465.590000 723.500000 466.410000 ;
      RECT 657.500000 465.590000 699.500000 466.410000 ;
      RECT 607.500000 465.590000 649.500000 466.410000 ;
      RECT 557.500000 465.590000 599.500000 466.410000 ;
      RECT 507.500000 465.590000 549.500000 466.410000 ;
      RECT 457.500000 465.590000 499.500000 466.410000 ;
      RECT 407.500000 465.590000 449.500000 466.410000 ;
      RECT 357.500000 465.590000 399.500000 466.410000 ;
      RECT 307.500000 465.590000 349.500000 466.410000 ;
      RECT 257.500000 465.590000 299.500000 466.410000 ;
      RECT 207.500000 465.590000 249.500000 466.410000 ;
      RECT 157.500000 465.590000 199.500000 466.410000 ;
      RECT 107.500000 465.590000 149.500000 466.410000 ;
      RECT 57.500000 465.590000 99.500000 466.410000 ;
      RECT 15.500000 465.590000 49.500000 466.410000 ;
      RECT 1157.500000 464.410000 1158.500000 465.590000 ;
      RECT 1139.000000 464.410000 1149.500000 467.590000 ;
      RECT 736.500000 464.410000 739.000000 467.590000 ;
      RECT 722.500000 464.410000 723.500000 465.590000 ;
      RECT 707.500000 464.410000 708.500000 465.590000 ;
      RECT 666.500000 464.410000 699.500000 465.590000 ;
      RECT 657.500000 464.410000 658.500000 465.590000 ;
      RECT 616.500000 464.410000 649.500000 465.590000 ;
      RECT 607.500000 464.410000 608.500000 465.590000 ;
      RECT 566.500000 464.410000 599.500000 465.590000 ;
      RECT 557.500000 464.410000 558.500000 465.590000 ;
      RECT 516.500000 464.410000 549.500000 465.590000 ;
      RECT 507.500000 464.410000 508.500000 465.590000 ;
      RECT 466.500000 464.410000 499.500000 465.590000 ;
      RECT 457.500000 464.410000 458.500000 465.590000 ;
      RECT 416.500000 464.410000 449.500000 465.590000 ;
      RECT 407.500000 464.410000 408.500000 465.590000 ;
      RECT 366.500000 464.410000 399.500000 465.590000 ;
      RECT 357.500000 464.410000 358.500000 465.590000 ;
      RECT 316.500000 464.410000 349.500000 465.590000 ;
      RECT 307.500000 464.410000 308.500000 465.590000 ;
      RECT 266.500000 464.410000 299.500000 465.590000 ;
      RECT 257.500000 464.410000 258.500000 465.590000 ;
      RECT 216.500000 464.410000 249.500000 465.590000 ;
      RECT 207.500000 464.410000 208.500000 465.590000 ;
      RECT 166.500000 464.410000 199.500000 465.590000 ;
      RECT 157.500000 464.410000 158.500000 465.590000 ;
      RECT 116.500000 464.410000 149.500000 465.590000 ;
      RECT 107.500000 464.410000 108.500000 465.590000 ;
      RECT 66.500000 464.410000 99.500000 465.590000 ;
      RECT 57.500000 464.410000 58.500000 465.590000 ;
      RECT 29.500000 464.410000 49.500000 465.590000 ;
      RECT 15.500000 464.410000 16.500000 465.590000 ;
      RECT 0.000000 464.410000 2.500000 467.590000 ;
      RECT 1139.000000 463.590000 1158.500000 464.410000 ;
      RECT 722.500000 463.590000 739.000000 464.410000 ;
      RECT 666.500000 463.590000 708.500000 464.410000 ;
      RECT 616.500000 463.590000 658.500000 464.410000 ;
      RECT 566.500000 463.590000 608.500000 464.410000 ;
      RECT 516.500000 463.590000 558.500000 464.410000 ;
      RECT 466.500000 463.590000 508.500000 464.410000 ;
      RECT 416.500000 463.590000 458.500000 464.410000 ;
      RECT 366.500000 463.590000 408.500000 464.410000 ;
      RECT 316.500000 463.590000 358.500000 464.410000 ;
      RECT 266.500000 463.590000 308.500000 464.410000 ;
      RECT 216.500000 463.590000 258.500000 464.410000 ;
      RECT 166.500000 463.590000 208.500000 464.410000 ;
      RECT 116.500000 463.590000 158.500000 464.410000 ;
      RECT 66.500000 463.590000 108.500000 464.410000 ;
      RECT 29.500000 463.590000 58.500000 464.410000 ;
      RECT 0.000000 463.590000 16.500000 464.410000 ;
      RECT 1166.500000 462.410000 1186.000000 465.590000 ;
      RECT 1157.500000 462.410000 1158.500000 463.590000 ;
      RECT 722.500000 462.410000 723.500000 463.590000 ;
      RECT 707.500000 462.410000 708.500000 463.590000 ;
      RECT 666.500000 462.410000 699.500000 463.590000 ;
      RECT 657.500000 462.410000 658.500000 463.590000 ;
      RECT 616.500000 462.410000 649.500000 463.590000 ;
      RECT 607.500000 462.410000 608.500000 463.590000 ;
      RECT 566.500000 462.410000 599.500000 463.590000 ;
      RECT 557.500000 462.410000 558.500000 463.590000 ;
      RECT 516.500000 462.410000 549.500000 463.590000 ;
      RECT 507.500000 462.410000 508.500000 463.590000 ;
      RECT 466.500000 462.410000 499.500000 463.590000 ;
      RECT 457.500000 462.410000 458.500000 463.590000 ;
      RECT 416.500000 462.410000 449.500000 463.590000 ;
      RECT 407.500000 462.410000 408.500000 463.590000 ;
      RECT 366.500000 462.410000 399.500000 463.590000 ;
      RECT 357.500000 462.410000 358.500000 463.590000 ;
      RECT 316.500000 462.410000 349.500000 463.590000 ;
      RECT 307.500000 462.410000 308.500000 463.590000 ;
      RECT 266.500000 462.410000 299.500000 463.590000 ;
      RECT 257.500000 462.410000 258.500000 463.590000 ;
      RECT 216.500000 462.410000 249.500000 463.590000 ;
      RECT 207.500000 462.410000 208.500000 463.590000 ;
      RECT 166.500000 462.410000 199.500000 463.590000 ;
      RECT 157.500000 462.410000 158.500000 463.590000 ;
      RECT 116.500000 462.410000 149.500000 463.590000 ;
      RECT 107.500000 462.410000 108.500000 463.590000 ;
      RECT 66.500000 462.410000 99.500000 463.590000 ;
      RECT 57.500000 462.410000 58.500000 463.590000 ;
      RECT 29.500000 462.410000 49.500000 463.590000 ;
      RECT 15.500000 462.410000 16.500000 463.590000 ;
      RECT 1157.500000 461.590000 1186.000000 462.410000 ;
      RECT 707.500000 461.590000 723.500000 462.410000 ;
      RECT 657.500000 461.590000 699.500000 462.410000 ;
      RECT 607.500000 461.590000 649.500000 462.410000 ;
      RECT 557.500000 461.590000 599.500000 462.410000 ;
      RECT 507.500000 461.590000 549.500000 462.410000 ;
      RECT 457.500000 461.590000 499.500000 462.410000 ;
      RECT 407.500000 461.590000 449.500000 462.410000 ;
      RECT 357.500000 461.590000 399.500000 462.410000 ;
      RECT 307.500000 461.590000 349.500000 462.410000 ;
      RECT 207.500000 461.590000 249.500000 462.410000 ;
      RECT 107.500000 461.590000 149.500000 462.410000 ;
      RECT 57.500000 461.590000 99.500000 462.410000 ;
      RECT 15.500000 461.590000 49.500000 462.410000 ;
      RECT 1157.500000 460.410000 1158.500000 461.590000 ;
      RECT 1139.000000 460.410000 1149.500000 463.590000 ;
      RECT 736.500000 460.410000 739.000000 463.590000 ;
      RECT 722.500000 460.410000 723.500000 461.590000 ;
      RECT 707.500000 460.410000 708.500000 461.590000 ;
      RECT 666.500000 460.410000 699.500000 461.590000 ;
      RECT 657.500000 460.410000 658.500000 461.590000 ;
      RECT 616.500000 460.410000 649.500000 461.590000 ;
      RECT 607.500000 460.410000 608.500000 461.590000 ;
      RECT 566.500000 460.410000 599.500000 461.590000 ;
      RECT 557.500000 460.410000 558.500000 461.590000 ;
      RECT 516.500000 460.410000 549.500000 461.590000 ;
      RECT 507.500000 460.410000 508.500000 461.590000 ;
      RECT 466.500000 460.410000 499.500000 461.590000 ;
      RECT 457.500000 460.410000 458.500000 461.590000 ;
      RECT 416.500000 460.410000 449.500000 461.590000 ;
      RECT 407.500000 460.410000 408.500000 461.590000 ;
      RECT 366.500000 460.410000 399.500000 461.590000 ;
      RECT 357.500000 460.410000 358.500000 461.590000 ;
      RECT 316.500000 460.410000 349.500000 461.590000 ;
      RECT 307.500000 460.410000 308.500000 461.590000 ;
      RECT 257.500000 460.410000 299.500000 462.410000 ;
      RECT 216.500000 460.410000 249.500000 461.590000 ;
      RECT 207.500000 460.410000 208.500000 461.590000 ;
      RECT 157.500000 460.410000 199.500000 462.410000 ;
      RECT 116.500000 460.410000 149.500000 461.590000 ;
      RECT 107.500000 460.410000 108.500000 461.590000 ;
      RECT 66.500000 460.410000 99.500000 461.590000 ;
      RECT 57.500000 460.410000 58.500000 461.590000 ;
      RECT 29.500000 460.410000 49.500000 461.590000 ;
      RECT 15.500000 460.410000 16.500000 461.590000 ;
      RECT 0.000000 460.410000 2.500000 463.590000 ;
      RECT 1139.000000 459.590000 1158.500000 460.410000 ;
      RECT 722.500000 459.590000 739.000000 460.410000 ;
      RECT 666.500000 459.590000 708.500000 460.410000 ;
      RECT 616.500000 459.590000 658.500000 460.410000 ;
      RECT 566.500000 459.590000 608.500000 460.410000 ;
      RECT 516.500000 459.590000 558.500000 460.410000 ;
      RECT 466.500000 459.590000 508.500000 460.410000 ;
      RECT 416.500000 459.590000 458.500000 460.410000 ;
      RECT 366.500000 459.590000 408.500000 460.410000 ;
      RECT 316.500000 459.590000 358.500000 460.410000 ;
      RECT 216.500000 459.590000 308.500000 460.410000 ;
      RECT 116.500000 459.590000 208.500000 460.410000 ;
      RECT 66.500000 459.590000 108.500000 460.410000 ;
      RECT 29.500000 459.590000 58.500000 460.410000 ;
      RECT 0.000000 459.590000 16.500000 460.410000 ;
      RECT 1166.500000 458.410000 1186.000000 461.590000 ;
      RECT 1157.500000 458.410000 1158.500000 459.590000 ;
      RECT 722.500000 458.410000 723.500000 459.590000 ;
      RECT 707.500000 458.410000 708.500000 459.590000 ;
      RECT 666.500000 458.410000 699.500000 459.590000 ;
      RECT 657.500000 458.410000 658.500000 459.590000 ;
      RECT 616.500000 458.410000 649.500000 459.590000 ;
      RECT 607.500000 458.410000 608.500000 459.590000 ;
      RECT 566.500000 458.410000 599.500000 459.590000 ;
      RECT 557.500000 458.410000 558.500000 459.590000 ;
      RECT 516.500000 458.410000 549.500000 459.590000 ;
      RECT 507.500000 458.410000 508.500000 459.590000 ;
      RECT 466.500000 458.410000 499.500000 459.590000 ;
      RECT 457.500000 458.410000 458.500000 459.590000 ;
      RECT 416.500000 458.410000 449.500000 459.590000 ;
      RECT 407.500000 458.410000 408.500000 459.590000 ;
      RECT 366.500000 458.410000 399.500000 459.590000 ;
      RECT 357.500000 458.410000 358.500000 459.590000 ;
      RECT 316.500000 458.410000 349.500000 459.590000 ;
      RECT 307.500000 458.410000 308.500000 459.590000 ;
      RECT 216.500000 458.410000 249.500000 459.590000 ;
      RECT 207.500000 458.410000 208.500000 459.590000 ;
      RECT 116.500000 458.410000 149.500000 459.590000 ;
      RECT 107.500000 458.410000 108.500000 459.590000 ;
      RECT 66.500000 458.410000 99.500000 459.590000 ;
      RECT 57.500000 458.410000 58.500000 459.590000 ;
      RECT 29.500000 458.410000 49.500000 459.590000 ;
      RECT 15.500000 458.410000 16.500000 459.590000 ;
      RECT 1157.500000 457.590000 1186.000000 458.410000 ;
      RECT 707.500000 457.590000 723.500000 458.410000 ;
      RECT 657.500000 457.590000 699.500000 458.410000 ;
      RECT 607.500000 457.590000 649.500000 458.410000 ;
      RECT 557.500000 457.590000 599.500000 458.410000 ;
      RECT 507.500000 457.590000 549.500000 458.410000 ;
      RECT 457.500000 457.590000 499.500000 458.410000 ;
      RECT 407.500000 457.590000 449.500000 458.410000 ;
      RECT 357.500000 457.590000 399.500000 458.410000 ;
      RECT 307.500000 457.590000 349.500000 458.410000 ;
      RECT 207.500000 457.590000 249.500000 458.410000 ;
      RECT 107.500000 457.590000 149.500000 458.410000 ;
      RECT 57.500000 457.590000 99.500000 458.410000 ;
      RECT 15.500000 457.590000 49.500000 458.410000 ;
      RECT 1157.500000 456.410000 1158.500000 457.590000 ;
      RECT 1139.000000 456.410000 1149.500000 459.590000 ;
      RECT 736.500000 456.410000 739.000000 459.590000 ;
      RECT 722.500000 456.410000 723.500000 457.590000 ;
      RECT 707.500000 456.410000 708.500000 457.590000 ;
      RECT 666.500000 456.410000 699.500000 457.590000 ;
      RECT 657.500000 456.410000 658.500000 457.590000 ;
      RECT 616.500000 456.410000 649.500000 457.590000 ;
      RECT 607.500000 456.410000 608.500000 457.590000 ;
      RECT 566.500000 456.410000 599.500000 457.590000 ;
      RECT 557.500000 456.410000 558.500000 457.590000 ;
      RECT 516.500000 456.410000 549.500000 457.590000 ;
      RECT 507.500000 456.410000 508.500000 457.590000 ;
      RECT 466.500000 456.410000 499.500000 457.590000 ;
      RECT 457.500000 456.410000 458.500000 457.590000 ;
      RECT 416.500000 456.410000 449.500000 457.590000 ;
      RECT 407.500000 456.410000 408.500000 457.590000 ;
      RECT 366.500000 456.410000 399.500000 457.590000 ;
      RECT 357.500000 456.410000 358.500000 457.590000 ;
      RECT 316.500000 456.410000 349.500000 457.590000 ;
      RECT 307.500000 456.410000 308.500000 457.590000 ;
      RECT 257.500000 456.410000 299.500000 459.590000 ;
      RECT 216.500000 456.410000 249.500000 457.590000 ;
      RECT 207.500000 456.410000 208.500000 457.590000 ;
      RECT 157.500000 456.410000 199.500000 459.590000 ;
      RECT 116.500000 456.410000 149.500000 457.590000 ;
      RECT 107.500000 456.410000 108.500000 457.590000 ;
      RECT 66.500000 456.410000 99.500000 457.590000 ;
      RECT 57.500000 456.410000 58.500000 457.590000 ;
      RECT 29.500000 456.410000 49.500000 457.590000 ;
      RECT 15.500000 456.410000 16.500000 457.590000 ;
      RECT 0.000000 456.410000 2.500000 459.590000 ;
      RECT 1139.000000 455.590000 1158.500000 456.410000 ;
      RECT 722.500000 455.590000 739.000000 456.410000 ;
      RECT 666.500000 455.590000 708.500000 456.410000 ;
      RECT 616.500000 455.590000 658.500000 456.410000 ;
      RECT 566.500000 455.590000 608.500000 456.410000 ;
      RECT 516.500000 455.590000 558.500000 456.410000 ;
      RECT 466.500000 455.590000 508.500000 456.410000 ;
      RECT 416.500000 455.590000 458.500000 456.410000 ;
      RECT 366.500000 455.590000 408.500000 456.410000 ;
      RECT 316.500000 455.590000 358.500000 456.410000 ;
      RECT 216.500000 455.590000 308.500000 456.410000 ;
      RECT 116.500000 455.590000 208.500000 456.410000 ;
      RECT 66.500000 455.590000 108.500000 456.410000 ;
      RECT 29.500000 455.590000 58.500000 456.410000 ;
      RECT 0.000000 455.590000 16.500000 456.410000 ;
      RECT 1166.500000 454.410000 1186.000000 457.590000 ;
      RECT 1157.500000 454.410000 1158.500000 455.590000 ;
      RECT 722.500000 454.410000 723.500000 455.590000 ;
      RECT 707.500000 454.410000 708.500000 455.590000 ;
      RECT 666.500000 454.410000 699.500000 455.590000 ;
      RECT 657.500000 454.410000 658.500000 455.590000 ;
      RECT 616.500000 454.410000 649.500000 455.590000 ;
      RECT 607.500000 454.410000 608.500000 455.590000 ;
      RECT 566.500000 454.410000 599.500000 455.590000 ;
      RECT 557.500000 454.410000 558.500000 455.590000 ;
      RECT 516.500000 454.410000 549.500000 455.590000 ;
      RECT 507.500000 454.410000 508.500000 455.590000 ;
      RECT 466.500000 454.410000 499.500000 455.590000 ;
      RECT 457.500000 454.410000 458.500000 455.590000 ;
      RECT 416.500000 454.410000 449.500000 455.590000 ;
      RECT 407.500000 454.410000 408.500000 455.590000 ;
      RECT 366.500000 454.410000 399.500000 455.590000 ;
      RECT 357.500000 454.410000 358.500000 455.590000 ;
      RECT 316.500000 454.410000 349.500000 455.590000 ;
      RECT 307.500000 454.410000 308.500000 455.590000 ;
      RECT 216.500000 454.410000 249.500000 455.590000 ;
      RECT 207.500000 454.410000 208.500000 455.590000 ;
      RECT 116.500000 454.410000 149.500000 455.590000 ;
      RECT 107.500000 454.410000 108.500000 455.590000 ;
      RECT 66.500000 454.410000 99.500000 455.590000 ;
      RECT 57.500000 454.410000 58.500000 455.590000 ;
      RECT 29.500000 454.410000 49.500000 455.590000 ;
      RECT 15.500000 454.410000 16.500000 455.590000 ;
      RECT 1157.500000 453.590000 1186.000000 454.410000 ;
      RECT 707.500000 453.590000 723.500000 454.410000 ;
      RECT 657.500000 453.590000 699.500000 454.410000 ;
      RECT 607.500000 453.590000 649.500000 454.410000 ;
      RECT 557.500000 453.590000 599.500000 454.410000 ;
      RECT 507.500000 453.590000 549.500000 454.410000 ;
      RECT 457.500000 453.590000 499.500000 454.410000 ;
      RECT 407.500000 453.590000 449.500000 454.410000 ;
      RECT 357.500000 453.590000 399.500000 454.410000 ;
      RECT 307.500000 453.590000 349.500000 454.410000 ;
      RECT 207.500000 453.590000 249.500000 454.410000 ;
      RECT 107.500000 453.590000 149.500000 454.410000 ;
      RECT 57.500000 453.590000 99.500000 454.410000 ;
      RECT 15.500000 453.590000 49.500000 454.410000 ;
      RECT 1157.500000 452.410000 1158.500000 453.590000 ;
      RECT 1139.000000 452.410000 1149.500000 455.590000 ;
      RECT 736.500000 452.410000 739.000000 455.590000 ;
      RECT 722.500000 452.410000 723.500000 453.590000 ;
      RECT 707.500000 452.410000 708.500000 453.590000 ;
      RECT 666.500000 452.410000 699.500000 453.590000 ;
      RECT 657.500000 452.410000 658.500000 453.590000 ;
      RECT 616.500000 452.410000 649.500000 453.590000 ;
      RECT 607.500000 452.410000 608.500000 453.590000 ;
      RECT 566.500000 452.410000 599.500000 453.590000 ;
      RECT 557.500000 452.410000 558.500000 453.590000 ;
      RECT 516.500000 452.410000 549.500000 453.590000 ;
      RECT 507.500000 452.410000 508.500000 453.590000 ;
      RECT 466.500000 452.410000 499.500000 453.590000 ;
      RECT 457.500000 452.410000 458.500000 453.590000 ;
      RECT 416.500000 452.410000 449.500000 453.590000 ;
      RECT 407.500000 452.410000 408.500000 453.590000 ;
      RECT 366.500000 452.410000 399.500000 453.590000 ;
      RECT 357.500000 452.410000 358.500000 453.590000 ;
      RECT 316.500000 452.410000 349.500000 453.590000 ;
      RECT 307.500000 452.410000 308.500000 453.590000 ;
      RECT 257.500000 452.410000 299.500000 455.590000 ;
      RECT 216.500000 452.410000 249.500000 453.590000 ;
      RECT 207.500000 452.410000 208.500000 453.590000 ;
      RECT 157.500000 452.410000 199.500000 455.590000 ;
      RECT 116.500000 452.410000 149.500000 453.590000 ;
      RECT 107.500000 452.410000 108.500000 453.590000 ;
      RECT 66.500000 452.410000 99.500000 453.590000 ;
      RECT 57.500000 452.410000 58.500000 453.590000 ;
      RECT 29.500000 452.410000 49.500000 453.590000 ;
      RECT 15.500000 452.410000 16.500000 453.590000 ;
      RECT 0.000000 452.410000 2.500000 455.590000 ;
      RECT 1139.000000 451.590000 1158.500000 452.410000 ;
      RECT 722.500000 451.590000 739.000000 452.410000 ;
      RECT 666.500000 451.590000 708.500000 452.410000 ;
      RECT 616.500000 451.590000 658.500000 452.410000 ;
      RECT 566.500000 451.590000 608.500000 452.410000 ;
      RECT 516.500000 451.590000 558.500000 452.410000 ;
      RECT 466.500000 451.590000 508.500000 452.410000 ;
      RECT 416.500000 451.590000 458.500000 452.410000 ;
      RECT 366.500000 451.590000 408.500000 452.410000 ;
      RECT 316.500000 451.590000 358.500000 452.410000 ;
      RECT 216.500000 451.590000 308.500000 452.410000 ;
      RECT 116.500000 451.590000 208.500000 452.410000 ;
      RECT 66.500000 451.590000 108.500000 452.410000 ;
      RECT 29.500000 451.590000 58.500000 452.410000 ;
      RECT 0.000000 451.590000 16.500000 452.410000 ;
      RECT 1166.500000 450.410000 1186.000000 453.590000 ;
      RECT 1157.500000 450.410000 1158.500000 451.590000 ;
      RECT 722.500000 450.410000 723.500000 451.590000 ;
      RECT 707.500000 450.410000 708.500000 451.590000 ;
      RECT 666.500000 450.410000 699.500000 451.590000 ;
      RECT 657.500000 450.410000 658.500000 451.590000 ;
      RECT 616.500000 450.410000 649.500000 451.590000 ;
      RECT 607.500000 450.410000 608.500000 451.590000 ;
      RECT 566.500000 450.410000 599.500000 451.590000 ;
      RECT 557.500000 450.410000 558.500000 451.590000 ;
      RECT 516.500000 450.410000 549.500000 451.590000 ;
      RECT 507.500000 450.410000 508.500000 451.590000 ;
      RECT 466.500000 450.410000 499.500000 451.590000 ;
      RECT 457.500000 450.410000 458.500000 451.590000 ;
      RECT 416.500000 450.410000 449.500000 451.590000 ;
      RECT 407.500000 450.410000 408.500000 451.590000 ;
      RECT 366.500000 450.410000 399.500000 451.590000 ;
      RECT 357.500000 450.410000 358.500000 451.590000 ;
      RECT 316.500000 450.410000 349.500000 451.590000 ;
      RECT 307.500000 450.410000 308.500000 451.590000 ;
      RECT 216.500000 450.410000 299.500000 451.590000 ;
      RECT 207.500000 450.410000 208.500000 451.590000 ;
      RECT 116.500000 450.410000 199.500000 451.590000 ;
      RECT 107.500000 450.410000 108.500000 451.590000 ;
      RECT 66.500000 450.410000 99.500000 451.590000 ;
      RECT 57.500000 450.410000 58.500000 451.590000 ;
      RECT 29.500000 450.410000 49.500000 451.590000 ;
      RECT 15.500000 450.410000 16.500000 451.590000 ;
      RECT 1157.500000 449.590000 1186.000000 450.410000 ;
      RECT 707.500000 449.590000 723.500000 450.410000 ;
      RECT 657.500000 449.590000 699.500000 450.410000 ;
      RECT 607.500000 449.590000 649.500000 450.410000 ;
      RECT 557.500000 449.590000 599.500000 450.410000 ;
      RECT 507.500000 449.590000 549.500000 450.410000 ;
      RECT 457.500000 449.590000 499.500000 450.410000 ;
      RECT 407.500000 449.590000 449.500000 450.410000 ;
      RECT 357.500000 449.590000 399.500000 450.410000 ;
      RECT 307.500000 449.590000 349.500000 450.410000 ;
      RECT 207.500000 449.590000 299.500000 450.410000 ;
      RECT 107.500000 449.590000 199.500000 450.410000 ;
      RECT 57.500000 449.590000 99.500000 450.410000 ;
      RECT 15.500000 449.590000 49.500000 450.410000 ;
      RECT 1157.500000 448.410000 1158.500000 449.590000 ;
      RECT 1139.000000 448.410000 1149.500000 451.590000 ;
      RECT 736.500000 448.410000 739.000000 451.590000 ;
      RECT 722.500000 448.410000 723.500000 449.590000 ;
      RECT 707.500000 448.410000 708.500000 449.590000 ;
      RECT 666.500000 448.410000 699.500000 449.590000 ;
      RECT 657.500000 448.410000 658.500000 449.590000 ;
      RECT 616.500000 448.410000 649.500000 449.590000 ;
      RECT 607.500000 448.410000 608.500000 449.590000 ;
      RECT 566.500000 448.410000 599.500000 449.590000 ;
      RECT 557.500000 448.410000 558.500000 449.590000 ;
      RECT 516.500000 448.410000 549.500000 449.590000 ;
      RECT 507.500000 448.410000 508.500000 449.590000 ;
      RECT 466.500000 448.410000 499.500000 449.590000 ;
      RECT 457.500000 448.410000 458.500000 449.590000 ;
      RECT 416.500000 448.410000 449.500000 449.590000 ;
      RECT 407.500000 448.410000 408.500000 449.590000 ;
      RECT 366.500000 448.410000 399.500000 449.590000 ;
      RECT 357.500000 448.410000 358.500000 449.590000 ;
      RECT 316.500000 448.410000 349.500000 449.590000 ;
      RECT 307.500000 448.410000 308.500000 449.590000 ;
      RECT 216.500000 448.410000 299.500000 449.590000 ;
      RECT 207.500000 448.410000 208.500000 449.590000 ;
      RECT 116.500000 448.410000 199.500000 449.590000 ;
      RECT 107.500000 448.410000 108.500000 449.590000 ;
      RECT 66.500000 448.410000 99.500000 449.590000 ;
      RECT 57.500000 448.410000 58.500000 449.590000 ;
      RECT 29.500000 448.410000 49.500000 449.590000 ;
      RECT 15.500000 448.410000 16.500000 449.590000 ;
      RECT 0.000000 448.410000 2.500000 451.590000 ;
      RECT 1139.000000 447.590000 1158.500000 448.410000 ;
      RECT 722.500000 447.590000 739.000000 448.410000 ;
      RECT 666.500000 447.590000 708.500000 448.410000 ;
      RECT 616.500000 447.590000 658.500000 448.410000 ;
      RECT 566.500000 447.590000 608.500000 448.410000 ;
      RECT 516.500000 447.590000 558.500000 448.410000 ;
      RECT 466.500000 447.590000 508.500000 448.410000 ;
      RECT 416.500000 447.590000 458.500000 448.410000 ;
      RECT 366.500000 447.590000 408.500000 448.410000 ;
      RECT 316.500000 447.590000 358.500000 448.410000 ;
      RECT 216.500000 447.590000 308.500000 448.410000 ;
      RECT 116.500000 447.590000 208.500000 448.410000 ;
      RECT 66.500000 447.590000 108.500000 448.410000 ;
      RECT 29.500000 447.590000 58.500000 448.410000 ;
      RECT 0.000000 447.590000 16.500000 448.410000 ;
      RECT 1166.500000 446.410000 1186.000000 449.590000 ;
      RECT 1157.500000 446.410000 1158.500000 447.590000 ;
      RECT 722.500000 446.410000 723.500000 447.590000 ;
      RECT 707.500000 446.410000 708.500000 447.590000 ;
      RECT 666.500000 446.410000 699.500000 447.590000 ;
      RECT 657.500000 446.410000 658.500000 447.590000 ;
      RECT 616.500000 446.410000 649.500000 447.590000 ;
      RECT 607.500000 446.410000 608.500000 447.590000 ;
      RECT 566.500000 446.410000 599.500000 447.590000 ;
      RECT 557.500000 446.410000 558.500000 447.590000 ;
      RECT 516.500000 446.410000 549.500000 447.590000 ;
      RECT 507.500000 446.410000 508.500000 447.590000 ;
      RECT 466.500000 446.410000 499.500000 447.590000 ;
      RECT 457.500000 446.410000 458.500000 447.590000 ;
      RECT 416.500000 446.410000 449.500000 447.590000 ;
      RECT 407.500000 446.410000 408.500000 447.590000 ;
      RECT 366.500000 446.410000 399.500000 447.590000 ;
      RECT 357.500000 446.410000 358.500000 447.590000 ;
      RECT 316.500000 446.410000 349.500000 447.590000 ;
      RECT 307.500000 446.410000 308.500000 447.590000 ;
      RECT 216.500000 446.410000 299.500000 447.590000 ;
      RECT 207.500000 446.410000 208.500000 447.590000 ;
      RECT 116.500000 446.410000 199.500000 447.590000 ;
      RECT 107.500000 446.410000 108.500000 447.590000 ;
      RECT 66.500000 446.410000 99.500000 447.590000 ;
      RECT 57.500000 446.410000 58.500000 447.590000 ;
      RECT 29.500000 446.410000 49.500000 447.590000 ;
      RECT 15.500000 446.410000 16.500000 447.590000 ;
      RECT 1139.000000 446.000000 1149.500000 447.590000 ;
      RECT 736.500000 446.000000 739.000000 447.590000 ;
      RECT 1157.500000 445.590000 1186.000000 446.410000 ;
      RECT 736.500000 445.590000 1149.500000 446.000000 ;
      RECT 707.500000 445.590000 723.500000 446.410000 ;
      RECT 657.500000 445.590000 699.500000 446.410000 ;
      RECT 607.500000 445.590000 649.500000 446.410000 ;
      RECT 557.500000 445.590000 599.500000 446.410000 ;
      RECT 507.500000 445.590000 549.500000 446.410000 ;
      RECT 457.500000 445.590000 499.500000 446.410000 ;
      RECT 407.500000 445.590000 449.500000 446.410000 ;
      RECT 357.500000 445.590000 399.500000 446.410000 ;
      RECT 307.500000 445.590000 349.500000 446.410000 ;
      RECT 207.500000 445.590000 299.500000 446.410000 ;
      RECT 107.500000 445.590000 199.500000 446.410000 ;
      RECT 57.500000 445.590000 99.500000 446.410000 ;
      RECT 15.500000 445.590000 49.500000 446.410000 ;
      RECT 1157.500000 444.410000 1158.500000 445.590000 ;
      RECT 1116.500000 444.410000 1149.500000 445.590000 ;
      RECT 736.500000 444.410000 758.500000 445.590000 ;
      RECT 722.500000 444.410000 723.500000 445.590000 ;
      RECT 707.500000 444.410000 708.500000 445.590000 ;
      RECT 666.500000 444.410000 699.500000 445.590000 ;
      RECT 657.500000 444.410000 658.500000 445.590000 ;
      RECT 616.500000 444.410000 649.500000 445.590000 ;
      RECT 607.500000 444.410000 608.500000 445.590000 ;
      RECT 566.500000 444.410000 599.500000 445.590000 ;
      RECT 557.500000 444.410000 558.500000 445.590000 ;
      RECT 516.500000 444.410000 549.500000 445.590000 ;
      RECT 507.500000 444.410000 508.500000 445.590000 ;
      RECT 466.500000 444.410000 499.500000 445.590000 ;
      RECT 457.500000 444.410000 458.500000 445.590000 ;
      RECT 416.500000 444.410000 449.500000 445.590000 ;
      RECT 407.500000 444.410000 408.500000 445.590000 ;
      RECT 366.500000 444.410000 399.500000 445.590000 ;
      RECT 357.500000 444.410000 358.500000 445.590000 ;
      RECT 316.500000 444.410000 349.500000 445.590000 ;
      RECT 307.500000 444.410000 308.500000 445.590000 ;
      RECT 216.500000 444.410000 299.500000 445.590000 ;
      RECT 207.500000 444.410000 208.500000 445.590000 ;
      RECT 116.500000 444.410000 199.500000 445.590000 ;
      RECT 107.500000 444.410000 108.500000 445.590000 ;
      RECT 66.500000 444.410000 99.500000 445.590000 ;
      RECT 57.500000 444.410000 58.500000 445.590000 ;
      RECT 29.500000 444.410000 49.500000 445.590000 ;
      RECT 15.500000 444.410000 16.500000 445.590000 ;
      RECT 0.000000 444.410000 2.500000 447.590000 ;
      RECT 1166.500000 443.590000 1186.000000 445.590000 ;
      RECT 1116.500000 443.590000 1158.500000 444.410000 ;
      RECT 1066.500000 443.590000 1108.500000 445.590000 ;
      RECT 1016.500000 443.590000 1058.500000 445.590000 ;
      RECT 966.500000 443.590000 1008.500000 445.590000 ;
      RECT 916.500000 443.590000 958.500000 445.590000 ;
      RECT 866.500000 443.590000 908.500000 445.590000 ;
      RECT 816.500000 443.590000 858.500000 445.590000 ;
      RECT 766.500000 443.590000 808.500000 445.590000 ;
      RECT 722.500000 443.590000 758.500000 444.410000 ;
      RECT 666.500000 443.590000 708.500000 444.410000 ;
      RECT 616.500000 443.590000 658.500000 444.410000 ;
      RECT 566.500000 443.590000 608.500000 444.410000 ;
      RECT 516.500000 443.590000 558.500000 444.410000 ;
      RECT 466.500000 443.590000 508.500000 444.410000 ;
      RECT 416.500000 443.590000 458.500000 444.410000 ;
      RECT 366.500000 443.590000 408.500000 444.410000 ;
      RECT 316.500000 443.590000 358.500000 444.410000 ;
      RECT 216.500000 443.590000 308.500000 444.410000 ;
      RECT 116.500000 443.590000 208.500000 444.410000 ;
      RECT 66.500000 443.590000 108.500000 444.410000 ;
      RECT 29.500000 443.590000 58.500000 444.410000 ;
      RECT 0.000000 443.590000 16.500000 444.410000 ;
      RECT 1166.500000 442.410000 1170.500000 443.590000 ;
      RECT 1157.500000 442.410000 1158.500000 443.590000 ;
      RECT 1116.500000 442.410000 1149.500000 443.590000 ;
      RECT 1107.500000 442.410000 1108.500000 443.590000 ;
      RECT 1066.500000 442.410000 1099.500000 443.590000 ;
      RECT 1057.500000 442.410000 1058.500000 443.590000 ;
      RECT 1016.500000 442.410000 1049.500000 443.590000 ;
      RECT 1007.500000 442.410000 1008.500000 443.590000 ;
      RECT 966.500000 442.410000 999.500000 443.590000 ;
      RECT 957.500000 442.410000 958.500000 443.590000 ;
      RECT 916.500000 442.410000 949.500000 443.590000 ;
      RECT 907.500000 442.410000 908.500000 443.590000 ;
      RECT 866.500000 442.410000 899.500000 443.590000 ;
      RECT 857.500000 442.410000 858.500000 443.590000 ;
      RECT 816.500000 442.410000 849.500000 443.590000 ;
      RECT 807.500000 442.410000 808.500000 443.590000 ;
      RECT 766.500000 442.410000 799.500000 443.590000 ;
      RECT 757.500000 442.410000 758.500000 443.590000 ;
      RECT 722.500000 442.410000 723.500000 443.590000 ;
      RECT 707.500000 442.410000 708.500000 443.590000 ;
      RECT 666.500000 442.410000 699.500000 443.590000 ;
      RECT 657.500000 442.410000 658.500000 443.590000 ;
      RECT 616.500000 442.410000 649.500000 443.590000 ;
      RECT 607.500000 442.410000 608.500000 443.590000 ;
      RECT 566.500000 442.410000 599.500000 443.590000 ;
      RECT 557.500000 442.410000 558.500000 443.590000 ;
      RECT 516.500000 442.410000 549.500000 443.590000 ;
      RECT 507.500000 442.410000 508.500000 443.590000 ;
      RECT 466.500000 442.410000 499.500000 443.590000 ;
      RECT 457.500000 442.410000 458.500000 443.590000 ;
      RECT 416.500000 442.410000 449.500000 443.590000 ;
      RECT 407.500000 442.410000 408.500000 443.590000 ;
      RECT 366.500000 442.410000 399.500000 443.590000 ;
      RECT 357.500000 442.410000 358.500000 443.590000 ;
      RECT 316.500000 442.410000 349.500000 443.590000 ;
      RECT 307.500000 442.410000 308.500000 443.590000 ;
      RECT 216.500000 442.410000 299.500000 443.590000 ;
      RECT 207.500000 442.410000 208.500000 443.590000 ;
      RECT 116.500000 442.410000 199.500000 443.590000 ;
      RECT 107.500000 442.410000 108.500000 443.590000 ;
      RECT 66.500000 442.410000 99.500000 443.590000 ;
      RECT 57.500000 442.410000 58.500000 443.590000 ;
      RECT 29.500000 442.410000 49.500000 443.590000 ;
      RECT 15.500000 442.410000 16.500000 443.590000 ;
      RECT 1157.500000 441.590000 1170.500000 442.410000 ;
      RECT 1107.500000 441.590000 1149.500000 442.410000 ;
      RECT 1057.500000 441.590000 1099.500000 442.410000 ;
      RECT 1007.500000 441.590000 1049.500000 442.410000 ;
      RECT 957.500000 441.590000 999.500000 442.410000 ;
      RECT 907.500000 441.590000 949.500000 442.410000 ;
      RECT 857.500000 441.590000 899.500000 442.410000 ;
      RECT 807.500000 441.590000 849.500000 442.410000 ;
      RECT 757.500000 441.590000 799.500000 442.410000 ;
      RECT 707.500000 441.590000 723.500000 442.410000 ;
      RECT 657.500000 441.590000 699.500000 442.410000 ;
      RECT 607.500000 441.590000 649.500000 442.410000 ;
      RECT 557.500000 441.590000 599.500000 442.410000 ;
      RECT 507.500000 441.590000 549.500000 442.410000 ;
      RECT 457.500000 441.590000 499.500000 442.410000 ;
      RECT 407.500000 441.590000 449.500000 442.410000 ;
      RECT 357.500000 441.590000 399.500000 442.410000 ;
      RECT 307.500000 441.590000 349.500000 442.410000 ;
      RECT 207.500000 441.590000 299.500000 442.410000 ;
      RECT 107.500000 441.590000 199.500000 442.410000 ;
      RECT 57.500000 441.590000 99.500000 442.410000 ;
      RECT 15.500000 441.590000 49.500000 442.410000 ;
      RECT 1183.500000 440.410000 1186.000000 443.590000 ;
      RECT 1166.500000 440.410000 1170.500000 441.590000 ;
      RECT 1157.500000 440.410000 1158.500000 441.590000 ;
      RECT 1116.500000 440.410000 1149.500000 441.590000 ;
      RECT 1107.500000 440.410000 1108.500000 441.590000 ;
      RECT 1066.500000 440.410000 1099.500000 441.590000 ;
      RECT 1057.500000 440.410000 1058.500000 441.590000 ;
      RECT 1016.500000 440.410000 1049.500000 441.590000 ;
      RECT 1007.500000 440.410000 1008.500000 441.590000 ;
      RECT 966.500000 440.410000 999.500000 441.590000 ;
      RECT 957.500000 440.410000 958.500000 441.590000 ;
      RECT 916.500000 440.410000 949.500000 441.590000 ;
      RECT 907.500000 440.410000 908.500000 441.590000 ;
      RECT 866.500000 440.410000 899.500000 441.590000 ;
      RECT 857.500000 440.410000 858.500000 441.590000 ;
      RECT 816.500000 440.410000 849.500000 441.590000 ;
      RECT 807.500000 440.410000 808.500000 441.590000 ;
      RECT 766.500000 440.410000 799.500000 441.590000 ;
      RECT 757.500000 440.410000 758.500000 441.590000 ;
      RECT 736.500000 440.410000 749.500000 443.590000 ;
      RECT 722.500000 440.410000 723.500000 441.590000 ;
      RECT 707.500000 440.410000 708.500000 441.590000 ;
      RECT 666.500000 440.410000 699.500000 441.590000 ;
      RECT 657.500000 440.410000 658.500000 441.590000 ;
      RECT 616.500000 440.410000 649.500000 441.590000 ;
      RECT 607.500000 440.410000 608.500000 441.590000 ;
      RECT 566.500000 440.410000 599.500000 441.590000 ;
      RECT 557.500000 440.410000 558.500000 441.590000 ;
      RECT 516.500000 440.410000 549.500000 441.590000 ;
      RECT 507.500000 440.410000 508.500000 441.590000 ;
      RECT 466.500000 440.410000 499.500000 441.590000 ;
      RECT 457.500000 440.410000 458.500000 441.590000 ;
      RECT 416.500000 440.410000 449.500000 441.590000 ;
      RECT 407.500000 440.410000 408.500000 441.590000 ;
      RECT 366.500000 440.410000 399.500000 441.590000 ;
      RECT 357.500000 440.410000 358.500000 441.590000 ;
      RECT 316.500000 440.410000 349.500000 441.590000 ;
      RECT 307.500000 440.410000 308.500000 441.590000 ;
      RECT 216.500000 440.410000 299.500000 441.590000 ;
      RECT 207.500000 440.410000 208.500000 441.590000 ;
      RECT 116.500000 440.410000 199.500000 441.590000 ;
      RECT 107.500000 440.410000 108.500000 441.590000 ;
      RECT 66.500000 440.410000 99.500000 441.590000 ;
      RECT 57.500000 440.410000 58.500000 441.590000 ;
      RECT 29.500000 440.410000 49.500000 441.590000 ;
      RECT 15.500000 440.410000 16.500000 441.590000 ;
      RECT 0.000000 440.410000 2.500000 443.590000 ;
      RECT 1166.500000 439.590000 1186.000000 440.410000 ;
      RECT 1116.500000 439.590000 1158.500000 440.410000 ;
      RECT 1066.500000 439.590000 1108.500000 440.410000 ;
      RECT 1016.500000 439.590000 1058.500000 440.410000 ;
      RECT 966.500000 439.590000 1008.500000 440.410000 ;
      RECT 916.500000 439.590000 958.500000 440.410000 ;
      RECT 866.500000 439.590000 908.500000 440.410000 ;
      RECT 816.500000 439.590000 858.500000 440.410000 ;
      RECT 766.500000 439.590000 808.500000 440.410000 ;
      RECT 722.500000 439.590000 758.500000 440.410000 ;
      RECT 666.500000 439.590000 708.500000 440.410000 ;
      RECT 616.500000 439.590000 658.500000 440.410000 ;
      RECT 566.500000 439.590000 608.500000 440.410000 ;
      RECT 516.500000 439.590000 558.500000 440.410000 ;
      RECT 466.500000 439.590000 508.500000 440.410000 ;
      RECT 416.500000 439.590000 458.500000 440.410000 ;
      RECT 366.500000 439.590000 408.500000 440.410000 ;
      RECT 316.500000 439.590000 358.500000 440.410000 ;
      RECT 216.500000 439.590000 308.500000 440.410000 ;
      RECT 116.500000 439.590000 208.500000 440.410000 ;
      RECT 66.500000 439.590000 108.500000 440.410000 ;
      RECT 29.500000 439.590000 58.500000 440.410000 ;
      RECT 0.000000 439.590000 16.500000 440.410000 ;
      RECT 1166.500000 438.410000 1170.500000 439.590000 ;
      RECT 1157.500000 438.410000 1158.500000 439.590000 ;
      RECT 1116.500000 438.410000 1149.500000 439.590000 ;
      RECT 1107.500000 438.410000 1108.500000 439.590000 ;
      RECT 1066.500000 438.410000 1099.500000 439.590000 ;
      RECT 1057.500000 438.410000 1058.500000 439.590000 ;
      RECT 1016.500000 438.410000 1049.500000 439.590000 ;
      RECT 1007.500000 438.410000 1008.500000 439.590000 ;
      RECT 966.500000 438.410000 999.500000 439.590000 ;
      RECT 957.500000 438.410000 958.500000 439.590000 ;
      RECT 916.500000 438.410000 949.500000 439.590000 ;
      RECT 907.500000 438.410000 908.500000 439.590000 ;
      RECT 866.500000 438.410000 899.500000 439.590000 ;
      RECT 857.500000 438.410000 858.500000 439.590000 ;
      RECT 816.500000 438.410000 849.500000 439.590000 ;
      RECT 807.500000 438.410000 808.500000 439.590000 ;
      RECT 766.500000 438.410000 799.500000 439.590000 ;
      RECT 757.500000 438.410000 758.500000 439.590000 ;
      RECT 722.500000 438.410000 723.500000 439.590000 ;
      RECT 707.500000 438.410000 708.500000 439.590000 ;
      RECT 666.500000 438.410000 699.500000 439.590000 ;
      RECT 657.500000 438.410000 658.500000 439.590000 ;
      RECT 616.500000 438.410000 649.500000 439.590000 ;
      RECT 607.500000 438.410000 608.500000 439.590000 ;
      RECT 566.500000 438.410000 599.500000 439.590000 ;
      RECT 557.500000 438.410000 558.500000 439.590000 ;
      RECT 516.500000 438.410000 549.500000 439.590000 ;
      RECT 507.500000 438.410000 508.500000 439.590000 ;
      RECT 466.500000 438.410000 499.500000 439.590000 ;
      RECT 457.500000 438.410000 458.500000 439.590000 ;
      RECT 416.500000 438.410000 449.500000 439.590000 ;
      RECT 407.500000 438.410000 408.500000 439.590000 ;
      RECT 366.500000 438.410000 399.500000 439.590000 ;
      RECT 357.500000 438.410000 358.500000 439.590000 ;
      RECT 316.500000 438.410000 349.500000 439.590000 ;
      RECT 307.500000 438.410000 308.500000 439.590000 ;
      RECT 216.500000 438.410000 299.500000 439.590000 ;
      RECT 207.500000 438.410000 208.500000 439.590000 ;
      RECT 116.500000 438.410000 199.500000 439.590000 ;
      RECT 107.500000 438.410000 108.500000 439.590000 ;
      RECT 66.500000 438.410000 99.500000 439.590000 ;
      RECT 57.500000 438.410000 58.500000 439.590000 ;
      RECT 29.500000 438.410000 49.500000 439.590000 ;
      RECT 15.500000 438.410000 16.500000 439.590000 ;
      RECT 1157.500000 437.590000 1170.500000 438.410000 ;
      RECT 1107.500000 437.590000 1149.500000 438.410000 ;
      RECT 1057.500000 437.590000 1099.500000 438.410000 ;
      RECT 1007.500000 437.590000 1049.500000 438.410000 ;
      RECT 957.500000 437.590000 999.500000 438.410000 ;
      RECT 907.500000 437.590000 949.500000 438.410000 ;
      RECT 857.500000 437.590000 899.500000 438.410000 ;
      RECT 807.500000 437.590000 849.500000 438.410000 ;
      RECT 757.500000 437.590000 799.500000 438.410000 ;
      RECT 707.500000 437.590000 723.500000 438.410000 ;
      RECT 657.500000 437.590000 699.500000 438.410000 ;
      RECT 607.500000 437.590000 649.500000 438.410000 ;
      RECT 557.500000 437.590000 599.500000 438.410000 ;
      RECT 507.500000 437.590000 549.500000 438.410000 ;
      RECT 457.500000 437.590000 499.500000 438.410000 ;
      RECT 407.500000 437.590000 449.500000 438.410000 ;
      RECT 357.500000 437.590000 399.500000 438.410000 ;
      RECT 307.500000 437.590000 349.500000 438.410000 ;
      RECT 207.500000 437.590000 299.500000 438.410000 ;
      RECT 107.500000 437.590000 199.500000 438.410000 ;
      RECT 57.500000 437.590000 99.500000 438.410000 ;
      RECT 15.500000 437.590000 49.500000 438.410000 ;
      RECT 1183.500000 436.410000 1186.000000 439.590000 ;
      RECT 1166.500000 436.410000 1170.500000 437.590000 ;
      RECT 1157.500000 436.410000 1158.500000 437.590000 ;
      RECT 1116.500000 436.410000 1149.500000 437.590000 ;
      RECT 1107.500000 436.410000 1108.500000 437.590000 ;
      RECT 1066.500000 436.410000 1099.500000 437.590000 ;
      RECT 1057.500000 436.410000 1058.500000 437.590000 ;
      RECT 1016.500000 436.410000 1049.500000 437.590000 ;
      RECT 1007.500000 436.410000 1008.500000 437.590000 ;
      RECT 966.500000 436.410000 999.500000 437.590000 ;
      RECT 957.500000 436.410000 958.500000 437.590000 ;
      RECT 916.500000 436.410000 949.500000 437.590000 ;
      RECT 907.500000 436.410000 908.500000 437.590000 ;
      RECT 866.500000 436.410000 899.500000 437.590000 ;
      RECT 857.500000 436.410000 858.500000 437.590000 ;
      RECT 816.500000 436.410000 849.500000 437.590000 ;
      RECT 807.500000 436.410000 808.500000 437.590000 ;
      RECT 766.500000 436.410000 799.500000 437.590000 ;
      RECT 757.500000 436.410000 758.500000 437.590000 ;
      RECT 736.500000 436.410000 749.500000 439.590000 ;
      RECT 722.500000 436.410000 723.500000 437.590000 ;
      RECT 707.500000 436.410000 708.500000 437.590000 ;
      RECT 666.500000 436.410000 699.500000 437.590000 ;
      RECT 657.500000 436.410000 658.500000 437.590000 ;
      RECT 616.500000 436.410000 649.500000 437.590000 ;
      RECT 607.500000 436.410000 608.500000 437.590000 ;
      RECT 566.500000 436.410000 599.500000 437.590000 ;
      RECT 557.500000 436.410000 558.500000 437.590000 ;
      RECT 516.500000 436.410000 549.500000 437.590000 ;
      RECT 507.500000 436.410000 508.500000 437.590000 ;
      RECT 466.500000 436.410000 499.500000 437.590000 ;
      RECT 457.500000 436.410000 458.500000 437.590000 ;
      RECT 416.500000 436.410000 449.500000 437.590000 ;
      RECT 407.500000 436.410000 408.500000 437.590000 ;
      RECT 366.500000 436.410000 399.500000 437.590000 ;
      RECT 357.500000 436.410000 358.500000 437.590000 ;
      RECT 316.500000 436.410000 349.500000 437.590000 ;
      RECT 307.500000 436.410000 308.500000 437.590000 ;
      RECT 216.500000 436.410000 299.500000 437.590000 ;
      RECT 207.500000 436.410000 208.500000 437.590000 ;
      RECT 116.500000 436.410000 199.500000 437.590000 ;
      RECT 107.500000 436.410000 108.500000 437.590000 ;
      RECT 66.500000 436.410000 99.500000 437.590000 ;
      RECT 57.500000 436.410000 58.500000 437.590000 ;
      RECT 29.500000 436.410000 49.500000 437.590000 ;
      RECT 15.500000 436.410000 16.500000 437.590000 ;
      RECT 0.000000 436.410000 2.500000 439.590000 ;
      RECT 1166.500000 435.590000 1186.000000 436.410000 ;
      RECT 1116.500000 435.590000 1158.500000 436.410000 ;
      RECT 1066.500000 435.590000 1108.500000 436.410000 ;
      RECT 1016.500000 435.590000 1058.500000 436.410000 ;
      RECT 966.500000 435.590000 1008.500000 436.410000 ;
      RECT 916.500000 435.590000 958.500000 436.410000 ;
      RECT 866.500000 435.590000 908.500000 436.410000 ;
      RECT 816.500000 435.590000 858.500000 436.410000 ;
      RECT 766.500000 435.590000 808.500000 436.410000 ;
      RECT 722.500000 435.590000 758.500000 436.410000 ;
      RECT 666.500000 435.590000 708.500000 436.410000 ;
      RECT 616.500000 435.590000 658.500000 436.410000 ;
      RECT 566.500000 435.590000 608.500000 436.410000 ;
      RECT 516.500000 435.590000 558.500000 436.410000 ;
      RECT 466.500000 435.590000 508.500000 436.410000 ;
      RECT 416.500000 435.590000 458.500000 436.410000 ;
      RECT 366.500000 435.590000 408.500000 436.410000 ;
      RECT 316.500000 435.590000 358.500000 436.410000 ;
      RECT 216.500000 435.590000 308.500000 436.410000 ;
      RECT 116.500000 435.590000 208.500000 436.410000 ;
      RECT 66.500000 435.590000 108.500000 436.410000 ;
      RECT 29.500000 435.590000 58.500000 436.410000 ;
      RECT 0.000000 435.590000 16.500000 436.410000 ;
      RECT 1166.500000 434.410000 1170.500000 435.590000 ;
      RECT 1157.500000 434.410000 1158.500000 435.590000 ;
      RECT 1116.500000 434.410000 1149.500000 435.590000 ;
      RECT 1107.500000 434.410000 1108.500000 435.590000 ;
      RECT 1066.500000 434.410000 1099.500000 435.590000 ;
      RECT 1057.500000 434.410000 1058.500000 435.590000 ;
      RECT 1016.500000 434.410000 1049.500000 435.590000 ;
      RECT 1007.500000 434.410000 1008.500000 435.590000 ;
      RECT 966.500000 434.410000 999.500000 435.590000 ;
      RECT 957.500000 434.410000 958.500000 435.590000 ;
      RECT 916.500000 434.410000 949.500000 435.590000 ;
      RECT 907.500000 434.410000 908.500000 435.590000 ;
      RECT 866.500000 434.410000 899.500000 435.590000 ;
      RECT 857.500000 434.410000 858.500000 435.590000 ;
      RECT 816.500000 434.410000 849.500000 435.590000 ;
      RECT 807.500000 434.410000 808.500000 435.590000 ;
      RECT 766.500000 434.410000 799.500000 435.590000 ;
      RECT 757.500000 434.410000 758.500000 435.590000 ;
      RECT 722.500000 434.410000 723.500000 435.590000 ;
      RECT 707.500000 434.410000 708.500000 435.590000 ;
      RECT 666.500000 434.410000 699.500000 435.590000 ;
      RECT 657.500000 434.410000 658.500000 435.590000 ;
      RECT 616.500000 434.410000 649.500000 435.590000 ;
      RECT 607.500000 434.410000 608.500000 435.590000 ;
      RECT 566.500000 434.410000 599.500000 435.590000 ;
      RECT 557.500000 434.410000 558.500000 435.590000 ;
      RECT 516.500000 434.410000 549.500000 435.590000 ;
      RECT 507.500000 434.410000 508.500000 435.590000 ;
      RECT 466.500000 434.410000 499.500000 435.590000 ;
      RECT 457.500000 434.410000 458.500000 435.590000 ;
      RECT 416.500000 434.410000 449.500000 435.590000 ;
      RECT 407.500000 434.410000 408.500000 435.590000 ;
      RECT 366.500000 434.410000 399.500000 435.590000 ;
      RECT 357.500000 434.410000 358.500000 435.590000 ;
      RECT 316.500000 434.410000 349.500000 435.590000 ;
      RECT 307.500000 434.410000 308.500000 435.590000 ;
      RECT 216.500000 434.410000 299.500000 435.590000 ;
      RECT 207.500000 434.410000 208.500000 435.590000 ;
      RECT 116.500000 434.410000 199.500000 435.590000 ;
      RECT 107.500000 434.410000 108.500000 435.590000 ;
      RECT 66.500000 434.410000 99.500000 435.590000 ;
      RECT 57.500000 434.410000 58.500000 435.590000 ;
      RECT 29.500000 434.410000 49.500000 435.590000 ;
      RECT 15.500000 434.410000 16.500000 435.590000 ;
      RECT 1157.500000 433.590000 1170.500000 434.410000 ;
      RECT 1107.500000 433.590000 1149.500000 434.410000 ;
      RECT 1057.500000 433.590000 1099.500000 434.410000 ;
      RECT 1007.500000 433.590000 1049.500000 434.410000 ;
      RECT 957.500000 433.590000 999.500000 434.410000 ;
      RECT 907.500000 433.590000 949.500000 434.410000 ;
      RECT 857.500000 433.590000 899.500000 434.410000 ;
      RECT 807.500000 433.590000 849.500000 434.410000 ;
      RECT 757.500000 433.590000 799.500000 434.410000 ;
      RECT 707.500000 433.590000 723.500000 434.410000 ;
      RECT 657.500000 433.590000 699.500000 434.410000 ;
      RECT 607.500000 433.590000 649.500000 434.410000 ;
      RECT 557.500000 433.590000 599.500000 434.410000 ;
      RECT 507.500000 433.590000 549.500000 434.410000 ;
      RECT 457.500000 433.590000 499.500000 434.410000 ;
      RECT 407.500000 433.590000 449.500000 434.410000 ;
      RECT 357.500000 433.590000 399.500000 434.410000 ;
      RECT 307.500000 433.590000 349.500000 434.410000 ;
      RECT 207.500000 433.590000 299.500000 434.410000 ;
      RECT 107.500000 433.590000 199.500000 434.410000 ;
      RECT 57.500000 433.590000 99.500000 434.410000 ;
      RECT 15.500000 433.590000 49.500000 434.410000 ;
      RECT 1183.500000 432.410000 1186.000000 435.590000 ;
      RECT 1166.500000 432.410000 1170.500000 433.590000 ;
      RECT 1157.500000 432.410000 1158.500000 433.590000 ;
      RECT 1116.500000 432.410000 1149.500000 433.590000 ;
      RECT 1107.500000 432.410000 1108.500000 433.590000 ;
      RECT 1066.500000 432.410000 1099.500000 433.590000 ;
      RECT 1057.500000 432.410000 1058.500000 433.590000 ;
      RECT 1016.500000 432.410000 1049.500000 433.590000 ;
      RECT 1007.500000 432.410000 1008.500000 433.590000 ;
      RECT 966.500000 432.410000 999.500000 433.590000 ;
      RECT 957.500000 432.410000 958.500000 433.590000 ;
      RECT 916.500000 432.410000 949.500000 433.590000 ;
      RECT 907.500000 432.410000 908.500000 433.590000 ;
      RECT 866.500000 432.410000 899.500000 433.590000 ;
      RECT 857.500000 432.410000 858.500000 433.590000 ;
      RECT 816.500000 432.410000 849.500000 433.590000 ;
      RECT 807.500000 432.410000 808.500000 433.590000 ;
      RECT 766.500000 432.410000 799.500000 433.590000 ;
      RECT 757.500000 432.410000 758.500000 433.590000 ;
      RECT 736.500000 432.410000 749.500000 435.590000 ;
      RECT 722.500000 432.410000 723.500000 433.590000 ;
      RECT 707.500000 432.410000 708.500000 433.590000 ;
      RECT 666.500000 432.410000 699.500000 433.590000 ;
      RECT 657.500000 432.410000 658.500000 433.590000 ;
      RECT 616.500000 432.410000 649.500000 433.590000 ;
      RECT 607.500000 432.410000 608.500000 433.590000 ;
      RECT 566.500000 432.410000 599.500000 433.590000 ;
      RECT 557.500000 432.410000 558.500000 433.590000 ;
      RECT 516.500000 432.410000 549.500000 433.590000 ;
      RECT 507.500000 432.410000 508.500000 433.590000 ;
      RECT 466.500000 432.410000 499.500000 433.590000 ;
      RECT 457.500000 432.410000 458.500000 433.590000 ;
      RECT 416.500000 432.410000 449.500000 433.590000 ;
      RECT 407.500000 432.410000 408.500000 433.590000 ;
      RECT 366.500000 432.410000 399.500000 433.590000 ;
      RECT 357.500000 432.410000 358.500000 433.590000 ;
      RECT 316.500000 432.410000 349.500000 433.590000 ;
      RECT 307.500000 432.410000 308.500000 433.590000 ;
      RECT 216.500000 432.410000 299.500000 433.590000 ;
      RECT 207.500000 432.410000 208.500000 433.590000 ;
      RECT 116.500000 432.410000 199.500000 433.590000 ;
      RECT 107.500000 432.410000 108.500000 433.590000 ;
      RECT 66.500000 432.410000 99.500000 433.590000 ;
      RECT 57.500000 432.410000 58.500000 433.590000 ;
      RECT 29.500000 432.410000 49.500000 433.590000 ;
      RECT 15.500000 432.410000 16.500000 433.590000 ;
      RECT 0.000000 432.410000 2.500000 435.590000 ;
      RECT 1166.500000 431.590000 1186.000000 432.410000 ;
      RECT 1116.500000 431.590000 1158.500000 432.410000 ;
      RECT 1066.500000 431.590000 1108.500000 432.410000 ;
      RECT 1016.500000 431.590000 1058.500000 432.410000 ;
      RECT 966.500000 431.590000 1008.500000 432.410000 ;
      RECT 916.500000 431.590000 958.500000 432.410000 ;
      RECT 866.500000 431.590000 908.500000 432.410000 ;
      RECT 816.500000 431.590000 858.500000 432.410000 ;
      RECT 766.500000 431.590000 808.500000 432.410000 ;
      RECT 722.500000 431.590000 758.500000 432.410000 ;
      RECT 666.500000 431.590000 708.500000 432.410000 ;
      RECT 616.500000 431.590000 658.500000 432.410000 ;
      RECT 566.500000 431.590000 608.500000 432.410000 ;
      RECT 516.500000 431.590000 558.500000 432.410000 ;
      RECT 466.500000 431.590000 508.500000 432.410000 ;
      RECT 416.500000 431.590000 458.500000 432.410000 ;
      RECT 366.500000 431.590000 408.500000 432.410000 ;
      RECT 316.500000 431.590000 358.500000 432.410000 ;
      RECT 216.500000 431.590000 308.500000 432.410000 ;
      RECT 116.500000 431.590000 208.500000 432.410000 ;
      RECT 66.500000 431.590000 108.500000 432.410000 ;
      RECT 29.500000 431.590000 58.500000 432.410000 ;
      RECT 0.000000 431.590000 16.500000 432.410000 ;
      RECT 1166.500000 430.410000 1170.500000 431.590000 ;
      RECT 1157.500000 430.410000 1158.500000 431.590000 ;
      RECT 1116.500000 430.410000 1149.500000 431.590000 ;
      RECT 1107.500000 430.410000 1108.500000 431.590000 ;
      RECT 1066.500000 430.410000 1099.500000 431.590000 ;
      RECT 1057.500000 430.410000 1058.500000 431.590000 ;
      RECT 1016.500000 430.410000 1049.500000 431.590000 ;
      RECT 1007.500000 430.410000 1008.500000 431.590000 ;
      RECT 966.500000 430.410000 999.500000 431.590000 ;
      RECT 957.500000 430.410000 958.500000 431.590000 ;
      RECT 916.500000 430.410000 949.500000 431.590000 ;
      RECT 907.500000 430.410000 908.500000 431.590000 ;
      RECT 866.500000 430.410000 899.500000 431.590000 ;
      RECT 857.500000 430.410000 858.500000 431.590000 ;
      RECT 816.500000 430.410000 849.500000 431.590000 ;
      RECT 807.500000 430.410000 808.500000 431.590000 ;
      RECT 766.500000 430.410000 799.500000 431.590000 ;
      RECT 757.500000 430.410000 758.500000 431.590000 ;
      RECT 722.500000 430.410000 749.500000 431.590000 ;
      RECT 707.500000 430.410000 708.500000 431.590000 ;
      RECT 666.500000 430.410000 699.500000 431.590000 ;
      RECT 657.500000 430.410000 658.500000 431.590000 ;
      RECT 616.500000 430.410000 649.500000 431.590000 ;
      RECT 607.500000 430.410000 608.500000 431.590000 ;
      RECT 566.500000 430.410000 599.500000 431.590000 ;
      RECT 557.500000 430.410000 558.500000 431.590000 ;
      RECT 516.500000 430.410000 549.500000 431.590000 ;
      RECT 507.500000 430.410000 508.500000 431.590000 ;
      RECT 466.500000 430.410000 499.500000 431.590000 ;
      RECT 457.500000 430.410000 458.500000 431.590000 ;
      RECT 416.500000 430.410000 449.500000 431.590000 ;
      RECT 407.500000 430.410000 408.500000 431.590000 ;
      RECT 366.500000 430.410000 399.500000 431.590000 ;
      RECT 357.500000 430.410000 358.500000 431.590000 ;
      RECT 316.500000 430.410000 349.500000 431.590000 ;
      RECT 307.500000 430.410000 308.500000 431.590000 ;
      RECT 216.500000 430.410000 299.500000 431.590000 ;
      RECT 207.500000 430.410000 208.500000 431.590000 ;
      RECT 116.500000 430.410000 199.500000 431.590000 ;
      RECT 107.500000 430.410000 108.500000 431.590000 ;
      RECT 66.500000 430.410000 99.500000 431.590000 ;
      RECT 57.500000 430.410000 58.500000 431.590000 ;
      RECT 29.500000 430.410000 49.500000 431.590000 ;
      RECT 15.500000 430.410000 16.500000 431.590000 ;
      RECT 1157.500000 429.590000 1170.500000 430.410000 ;
      RECT 1107.500000 429.590000 1149.500000 430.410000 ;
      RECT 1057.500000 429.590000 1099.500000 430.410000 ;
      RECT 1007.500000 429.590000 1049.500000 430.410000 ;
      RECT 957.500000 429.590000 999.500000 430.410000 ;
      RECT 907.500000 429.590000 949.500000 430.410000 ;
      RECT 857.500000 429.590000 899.500000 430.410000 ;
      RECT 807.500000 429.590000 849.500000 430.410000 ;
      RECT 757.500000 429.590000 799.500000 430.410000 ;
      RECT 707.500000 429.590000 749.500000 430.410000 ;
      RECT 657.500000 429.590000 699.500000 430.410000 ;
      RECT 607.500000 429.590000 649.500000 430.410000 ;
      RECT 557.500000 429.590000 599.500000 430.410000 ;
      RECT 507.500000 429.590000 549.500000 430.410000 ;
      RECT 457.500000 429.590000 499.500000 430.410000 ;
      RECT 407.500000 429.590000 449.500000 430.410000 ;
      RECT 357.500000 429.590000 399.500000 430.410000 ;
      RECT 307.500000 429.590000 349.500000 430.410000 ;
      RECT 207.500000 429.590000 299.500000 430.410000 ;
      RECT 107.500000 429.590000 199.500000 430.410000 ;
      RECT 57.500000 429.590000 99.500000 430.410000 ;
      RECT 15.500000 429.590000 49.500000 430.410000 ;
      RECT 1183.500000 428.410000 1186.000000 431.590000 ;
      RECT 1169.500000 428.410000 1170.500000 429.590000 ;
      RECT 1116.500000 428.410000 1149.500000 429.590000 ;
      RECT 1107.500000 428.410000 1108.500000 429.590000 ;
      RECT 1066.500000 428.410000 1099.500000 429.590000 ;
      RECT 1057.500000 428.410000 1058.500000 429.590000 ;
      RECT 1016.500000 428.410000 1049.500000 429.590000 ;
      RECT 1007.500000 428.410000 1008.500000 429.590000 ;
      RECT 966.500000 428.410000 999.500000 429.590000 ;
      RECT 957.500000 428.410000 958.500000 429.590000 ;
      RECT 916.500000 428.410000 949.500000 429.590000 ;
      RECT 907.500000 428.410000 908.500000 429.590000 ;
      RECT 866.500000 428.410000 899.500000 429.590000 ;
      RECT 857.500000 428.410000 858.500000 429.590000 ;
      RECT 816.500000 428.410000 849.500000 429.590000 ;
      RECT 807.500000 428.410000 808.500000 429.590000 ;
      RECT 766.500000 428.410000 799.500000 429.590000 ;
      RECT 757.500000 428.410000 758.500000 429.590000 ;
      RECT 722.500000 428.410000 749.500000 429.590000 ;
      RECT 707.500000 428.410000 709.500000 429.590000 ;
      RECT 666.500000 428.410000 699.500000 429.590000 ;
      RECT 657.500000 428.410000 658.500000 429.590000 ;
      RECT 616.500000 428.410000 649.500000 429.590000 ;
      RECT 607.500000 428.410000 608.500000 429.590000 ;
      RECT 566.500000 428.410000 599.500000 429.590000 ;
      RECT 557.500000 428.410000 558.500000 429.590000 ;
      RECT 516.500000 428.410000 549.500000 429.590000 ;
      RECT 507.500000 428.410000 508.500000 429.590000 ;
      RECT 466.500000 428.410000 499.500000 429.590000 ;
      RECT 457.500000 428.410000 458.500000 429.590000 ;
      RECT 416.500000 428.410000 449.500000 429.590000 ;
      RECT 407.500000 428.410000 408.500000 429.590000 ;
      RECT 366.500000 428.410000 399.500000 429.590000 ;
      RECT 357.500000 428.410000 358.500000 429.590000 ;
      RECT 316.500000 428.410000 349.500000 429.590000 ;
      RECT 307.500000 428.410000 308.500000 429.590000 ;
      RECT 216.500000 428.410000 299.500000 429.590000 ;
      RECT 207.500000 428.410000 208.500000 429.590000 ;
      RECT 116.500000 428.410000 199.500000 429.590000 ;
      RECT 107.500000 428.410000 108.500000 429.590000 ;
      RECT 66.500000 428.410000 99.500000 429.590000 ;
      RECT 57.500000 428.410000 58.500000 429.590000 ;
      RECT 29.500000 428.410000 49.500000 429.590000 ;
      RECT 15.500000 428.410000 16.500000 429.590000 ;
      RECT 0.000000 428.410000 2.500000 431.590000 ;
      RECT 1169.500000 427.590000 1186.000000 428.410000 ;
      RECT 1116.500000 427.590000 1156.500000 428.410000 ;
      RECT 1066.500000 427.590000 1108.500000 428.410000 ;
      RECT 1016.500000 427.590000 1058.500000 428.410000 ;
      RECT 966.500000 427.590000 1008.500000 428.410000 ;
      RECT 916.500000 427.590000 958.500000 428.410000 ;
      RECT 866.500000 427.590000 908.500000 428.410000 ;
      RECT 816.500000 427.590000 858.500000 428.410000 ;
      RECT 766.500000 427.590000 808.500000 428.410000 ;
      RECT 722.500000 427.590000 758.500000 428.410000 ;
      RECT 666.500000 427.590000 709.500000 428.410000 ;
      RECT 616.500000 427.590000 658.500000 428.410000 ;
      RECT 566.500000 427.590000 608.500000 428.410000 ;
      RECT 516.500000 427.590000 558.500000 428.410000 ;
      RECT 466.500000 427.590000 508.500000 428.410000 ;
      RECT 416.500000 427.590000 458.500000 428.410000 ;
      RECT 366.500000 427.590000 408.500000 428.410000 ;
      RECT 316.500000 427.590000 358.500000 428.410000 ;
      RECT 216.500000 427.590000 308.500000 428.410000 ;
      RECT 116.500000 427.590000 208.500000 428.410000 ;
      RECT 66.500000 427.590000 108.500000 428.410000 ;
      RECT 29.500000 427.590000 58.500000 428.410000 ;
      RECT 0.000000 427.590000 16.500000 428.410000 ;
      RECT 1169.500000 426.410000 1170.500000 427.590000 ;
      RECT 1116.500000 426.410000 1149.500000 427.590000 ;
      RECT 1107.500000 426.410000 1108.500000 427.590000 ;
      RECT 1066.500000 426.410000 1099.500000 427.590000 ;
      RECT 1057.500000 426.410000 1058.500000 427.590000 ;
      RECT 1016.500000 426.410000 1049.500000 427.590000 ;
      RECT 1007.500000 426.410000 1008.500000 427.590000 ;
      RECT 966.500000 426.410000 999.500000 427.590000 ;
      RECT 957.500000 426.410000 958.500000 427.590000 ;
      RECT 916.500000 426.410000 949.500000 427.590000 ;
      RECT 907.500000 426.410000 908.500000 427.590000 ;
      RECT 866.500000 426.410000 899.500000 427.590000 ;
      RECT 857.500000 426.410000 858.500000 427.590000 ;
      RECT 816.500000 426.410000 849.500000 427.590000 ;
      RECT 807.500000 426.410000 808.500000 427.590000 ;
      RECT 766.500000 426.410000 799.500000 427.590000 ;
      RECT 757.500000 426.410000 758.500000 427.590000 ;
      RECT 722.500000 426.410000 749.500000 427.590000 ;
      RECT 707.500000 426.410000 709.500000 427.590000 ;
      RECT 666.500000 426.410000 699.500000 427.590000 ;
      RECT 657.500000 426.410000 658.500000 427.590000 ;
      RECT 616.500000 426.410000 649.500000 427.590000 ;
      RECT 607.500000 426.410000 608.500000 427.590000 ;
      RECT 566.500000 426.410000 599.500000 427.590000 ;
      RECT 557.500000 426.410000 558.500000 427.590000 ;
      RECT 516.500000 426.410000 549.500000 427.590000 ;
      RECT 507.500000 426.410000 508.500000 427.590000 ;
      RECT 466.500000 426.410000 499.500000 427.590000 ;
      RECT 457.500000 426.410000 458.500000 427.590000 ;
      RECT 416.500000 426.410000 449.500000 427.590000 ;
      RECT 407.500000 426.410000 408.500000 427.590000 ;
      RECT 366.500000 426.410000 399.500000 427.590000 ;
      RECT 357.500000 426.410000 358.500000 427.590000 ;
      RECT 316.500000 426.410000 349.500000 427.590000 ;
      RECT 307.500000 426.410000 308.500000 427.590000 ;
      RECT 216.500000 426.410000 299.500000 427.590000 ;
      RECT 207.500000 426.410000 208.500000 427.590000 ;
      RECT 116.500000 426.410000 199.500000 427.590000 ;
      RECT 107.500000 426.410000 108.500000 427.590000 ;
      RECT 66.500000 426.410000 99.500000 427.590000 ;
      RECT 57.500000 426.410000 58.500000 427.590000 ;
      RECT 29.500000 426.410000 49.500000 427.590000 ;
      RECT 15.500000 426.410000 16.500000 427.590000 ;
      RECT 1157.500000 425.590000 1170.500000 426.410000 ;
      RECT 1107.500000 425.590000 1149.500000 426.410000 ;
      RECT 1057.500000 425.590000 1099.500000 426.410000 ;
      RECT 1007.500000 425.590000 1049.500000 426.410000 ;
      RECT 957.500000 425.590000 999.500000 426.410000 ;
      RECT 907.500000 425.590000 949.500000 426.410000 ;
      RECT 857.500000 425.590000 899.500000 426.410000 ;
      RECT 807.500000 425.590000 849.500000 426.410000 ;
      RECT 757.500000 425.590000 799.500000 426.410000 ;
      RECT 707.500000 425.590000 749.500000 426.410000 ;
      RECT 657.500000 425.590000 699.500000 426.410000 ;
      RECT 607.500000 425.590000 649.500000 426.410000 ;
      RECT 557.500000 425.590000 599.500000 426.410000 ;
      RECT 507.500000 425.590000 549.500000 426.410000 ;
      RECT 457.500000 425.590000 499.500000 426.410000 ;
      RECT 407.500000 425.590000 449.500000 426.410000 ;
      RECT 357.500000 425.590000 399.500000 426.410000 ;
      RECT 307.500000 425.590000 349.500000 426.410000 ;
      RECT 207.500000 425.590000 299.500000 426.410000 ;
      RECT 107.500000 425.590000 199.500000 426.410000 ;
      RECT 57.500000 425.590000 99.500000 426.410000 ;
      RECT 15.500000 425.590000 49.500000 426.410000 ;
      RECT 1183.500000 424.410000 1186.000000 427.590000 ;
      RECT 1169.500000 424.410000 1170.500000 425.590000 ;
      RECT 1116.500000 424.410000 1149.500000 425.590000 ;
      RECT 1107.500000 424.410000 1108.500000 425.590000 ;
      RECT 1066.500000 424.410000 1099.500000 425.590000 ;
      RECT 1057.500000 424.410000 1058.500000 425.590000 ;
      RECT 1016.500000 424.410000 1049.500000 425.590000 ;
      RECT 1007.500000 424.410000 1008.500000 425.590000 ;
      RECT 966.500000 424.410000 999.500000 425.590000 ;
      RECT 957.500000 424.410000 958.500000 425.590000 ;
      RECT 916.500000 424.410000 949.500000 425.590000 ;
      RECT 907.500000 424.410000 908.500000 425.590000 ;
      RECT 866.500000 424.410000 899.500000 425.590000 ;
      RECT 857.500000 424.410000 858.500000 425.590000 ;
      RECT 816.500000 424.410000 849.500000 425.590000 ;
      RECT 807.500000 424.410000 808.500000 425.590000 ;
      RECT 766.500000 424.410000 799.500000 425.590000 ;
      RECT 757.500000 424.410000 758.500000 425.590000 ;
      RECT 722.500000 424.410000 749.500000 425.590000 ;
      RECT 707.500000 424.410000 709.500000 425.590000 ;
      RECT 666.500000 424.410000 699.500000 425.590000 ;
      RECT 657.500000 424.410000 658.500000 425.590000 ;
      RECT 616.500000 424.410000 649.500000 425.590000 ;
      RECT 607.500000 424.410000 608.500000 425.590000 ;
      RECT 566.500000 424.410000 599.500000 425.590000 ;
      RECT 557.500000 424.410000 558.500000 425.590000 ;
      RECT 516.500000 424.410000 549.500000 425.590000 ;
      RECT 507.500000 424.410000 508.500000 425.590000 ;
      RECT 466.500000 424.410000 499.500000 425.590000 ;
      RECT 457.500000 424.410000 458.500000 425.590000 ;
      RECT 416.500000 424.410000 449.500000 425.590000 ;
      RECT 407.500000 424.410000 408.500000 425.590000 ;
      RECT 366.500000 424.410000 399.500000 425.590000 ;
      RECT 357.500000 424.410000 358.500000 425.590000 ;
      RECT 316.500000 424.410000 349.500000 425.590000 ;
      RECT 307.500000 424.410000 308.500000 425.590000 ;
      RECT 216.500000 424.410000 299.500000 425.590000 ;
      RECT 207.500000 424.410000 208.500000 425.590000 ;
      RECT 116.500000 424.410000 199.500000 425.590000 ;
      RECT 107.500000 424.410000 108.500000 425.590000 ;
      RECT 66.500000 424.410000 99.500000 425.590000 ;
      RECT 57.500000 424.410000 58.500000 425.590000 ;
      RECT 29.500000 424.410000 49.500000 425.590000 ;
      RECT 15.500000 424.410000 16.500000 425.590000 ;
      RECT 0.000000 424.410000 2.500000 427.590000 ;
      RECT 1169.500000 423.590000 1186.000000 424.410000 ;
      RECT 1116.500000 423.590000 1156.500000 424.410000 ;
      RECT 1066.500000 423.590000 1108.500000 424.410000 ;
      RECT 1016.500000 423.590000 1058.500000 424.410000 ;
      RECT 966.500000 423.590000 1008.500000 424.410000 ;
      RECT 916.500000 423.590000 958.500000 424.410000 ;
      RECT 866.500000 423.590000 908.500000 424.410000 ;
      RECT 816.500000 423.590000 858.500000 424.410000 ;
      RECT 766.500000 423.590000 808.500000 424.410000 ;
      RECT 722.500000 423.590000 758.500000 424.410000 ;
      RECT 666.500000 423.590000 709.500000 424.410000 ;
      RECT 616.500000 423.590000 658.500000 424.410000 ;
      RECT 566.500000 423.590000 608.500000 424.410000 ;
      RECT 516.500000 423.590000 558.500000 424.410000 ;
      RECT 466.500000 423.590000 508.500000 424.410000 ;
      RECT 416.500000 423.590000 458.500000 424.410000 ;
      RECT 366.500000 423.590000 408.500000 424.410000 ;
      RECT 316.500000 423.590000 358.500000 424.410000 ;
      RECT 216.500000 423.590000 308.500000 424.410000 ;
      RECT 116.500000 423.590000 208.500000 424.410000 ;
      RECT 66.500000 423.590000 108.500000 424.410000 ;
      RECT 29.500000 423.590000 58.500000 424.410000 ;
      RECT 0.000000 423.590000 16.500000 424.410000 ;
      RECT 1169.500000 422.410000 1170.500000 423.590000 ;
      RECT 1116.500000 422.410000 1149.500000 423.590000 ;
      RECT 1107.500000 422.410000 1108.500000 423.590000 ;
      RECT 1066.500000 422.410000 1099.500000 423.590000 ;
      RECT 1057.500000 422.410000 1058.500000 423.590000 ;
      RECT 1016.500000 422.410000 1049.500000 423.590000 ;
      RECT 1007.500000 422.410000 1008.500000 423.590000 ;
      RECT 966.500000 422.410000 999.500000 423.590000 ;
      RECT 957.500000 422.410000 958.500000 423.590000 ;
      RECT 916.500000 422.410000 949.500000 423.590000 ;
      RECT 907.500000 422.410000 908.500000 423.590000 ;
      RECT 866.500000 422.410000 899.500000 423.590000 ;
      RECT 857.500000 422.410000 858.500000 423.590000 ;
      RECT 816.500000 422.410000 849.500000 423.590000 ;
      RECT 807.500000 422.410000 808.500000 423.590000 ;
      RECT 766.500000 422.410000 799.500000 423.590000 ;
      RECT 757.500000 422.410000 758.500000 423.590000 ;
      RECT 722.500000 422.410000 749.500000 423.590000 ;
      RECT 707.500000 422.410000 709.500000 423.590000 ;
      RECT 666.500000 422.410000 699.500000 423.590000 ;
      RECT 657.500000 422.410000 658.500000 423.590000 ;
      RECT 616.500000 422.410000 649.500000 423.590000 ;
      RECT 607.500000 422.410000 608.500000 423.590000 ;
      RECT 566.500000 422.410000 599.500000 423.590000 ;
      RECT 557.500000 422.410000 558.500000 423.590000 ;
      RECT 516.500000 422.410000 549.500000 423.590000 ;
      RECT 507.500000 422.410000 508.500000 423.590000 ;
      RECT 466.500000 422.410000 499.500000 423.590000 ;
      RECT 457.500000 422.410000 458.500000 423.590000 ;
      RECT 416.500000 422.410000 449.500000 423.590000 ;
      RECT 407.500000 422.410000 408.500000 423.590000 ;
      RECT 366.500000 422.410000 399.500000 423.590000 ;
      RECT 357.500000 422.410000 358.500000 423.590000 ;
      RECT 316.500000 422.410000 349.500000 423.590000 ;
      RECT 307.500000 422.410000 308.500000 423.590000 ;
      RECT 216.500000 422.410000 299.500000 423.590000 ;
      RECT 207.500000 422.410000 208.500000 423.590000 ;
      RECT 116.500000 422.410000 199.500000 423.590000 ;
      RECT 107.500000 422.410000 108.500000 423.590000 ;
      RECT 66.500000 422.410000 99.500000 423.590000 ;
      RECT 57.500000 422.410000 58.500000 423.590000 ;
      RECT 29.500000 422.410000 49.500000 423.590000 ;
      RECT 15.500000 422.410000 16.500000 423.590000 ;
      RECT 1157.500000 421.590000 1170.500000 422.410000 ;
      RECT 1107.500000 421.590000 1149.500000 422.410000 ;
      RECT 1057.500000 421.590000 1099.500000 422.410000 ;
      RECT 1007.500000 421.590000 1049.500000 422.410000 ;
      RECT 957.500000 421.590000 999.500000 422.410000 ;
      RECT 907.500000 421.590000 949.500000 422.410000 ;
      RECT 857.500000 421.590000 899.500000 422.410000 ;
      RECT 807.500000 421.590000 849.500000 422.410000 ;
      RECT 757.500000 421.590000 799.500000 422.410000 ;
      RECT 707.500000 421.590000 749.500000 422.410000 ;
      RECT 657.500000 421.590000 699.500000 422.410000 ;
      RECT 607.500000 421.590000 649.500000 422.410000 ;
      RECT 557.500000 421.590000 599.500000 422.410000 ;
      RECT 507.500000 421.590000 549.500000 422.410000 ;
      RECT 457.500000 421.590000 499.500000 422.410000 ;
      RECT 407.500000 421.590000 449.500000 422.410000 ;
      RECT 357.500000 421.590000 399.500000 422.410000 ;
      RECT 307.500000 421.590000 349.500000 422.410000 ;
      RECT 207.500000 421.590000 299.500000 422.410000 ;
      RECT 107.500000 421.590000 199.500000 422.410000 ;
      RECT 57.500000 421.590000 99.500000 422.410000 ;
      RECT 15.500000 421.590000 49.500000 422.410000 ;
      RECT 1183.500000 420.410000 1186.000000 423.590000 ;
      RECT 1169.500000 420.410000 1170.500000 421.590000 ;
      RECT 1116.500000 420.410000 1149.500000 421.590000 ;
      RECT 1107.500000 420.410000 1108.500000 421.590000 ;
      RECT 1066.500000 420.410000 1099.500000 421.590000 ;
      RECT 1057.500000 420.410000 1058.500000 421.590000 ;
      RECT 1016.500000 420.410000 1049.500000 421.590000 ;
      RECT 1007.500000 420.410000 1008.500000 421.590000 ;
      RECT 966.500000 420.410000 999.500000 421.590000 ;
      RECT 957.500000 420.410000 958.500000 421.590000 ;
      RECT 916.500000 420.410000 949.500000 421.590000 ;
      RECT 907.500000 420.410000 908.500000 421.590000 ;
      RECT 866.500000 420.410000 899.500000 421.590000 ;
      RECT 857.500000 420.410000 858.500000 421.590000 ;
      RECT 816.500000 420.410000 849.500000 421.590000 ;
      RECT 807.500000 420.410000 808.500000 421.590000 ;
      RECT 766.500000 420.410000 799.500000 421.590000 ;
      RECT 757.500000 420.410000 758.500000 421.590000 ;
      RECT 722.500000 420.410000 749.500000 421.590000 ;
      RECT 707.500000 420.410000 709.500000 421.590000 ;
      RECT 666.500000 420.410000 699.500000 421.590000 ;
      RECT 657.500000 420.410000 658.500000 421.590000 ;
      RECT 616.500000 420.410000 649.500000 421.590000 ;
      RECT 607.500000 420.410000 608.500000 421.590000 ;
      RECT 566.500000 420.410000 599.500000 421.590000 ;
      RECT 557.500000 420.410000 558.500000 421.590000 ;
      RECT 516.500000 420.410000 549.500000 421.590000 ;
      RECT 507.500000 420.410000 508.500000 421.590000 ;
      RECT 466.500000 420.410000 499.500000 421.590000 ;
      RECT 457.500000 420.410000 458.500000 421.590000 ;
      RECT 416.500000 420.410000 449.500000 421.590000 ;
      RECT 407.500000 420.410000 408.500000 421.590000 ;
      RECT 366.500000 420.410000 399.500000 421.590000 ;
      RECT 357.500000 420.410000 358.500000 421.590000 ;
      RECT 316.500000 420.410000 349.500000 421.590000 ;
      RECT 307.500000 420.410000 308.500000 421.590000 ;
      RECT 216.500000 420.410000 299.500000 421.590000 ;
      RECT 207.500000 420.410000 208.500000 421.590000 ;
      RECT 116.500000 420.410000 199.500000 421.590000 ;
      RECT 107.500000 420.410000 108.500000 421.590000 ;
      RECT 66.500000 420.410000 99.500000 421.590000 ;
      RECT 57.500000 420.410000 58.500000 421.590000 ;
      RECT 29.500000 420.410000 49.500000 421.590000 ;
      RECT 15.500000 420.410000 16.500000 421.590000 ;
      RECT 0.000000 420.410000 2.500000 423.590000 ;
      RECT 1169.500000 419.590000 1186.000000 420.410000 ;
      RECT 1116.500000 419.590000 1156.500000 420.410000 ;
      RECT 1066.500000 419.590000 1108.500000 420.410000 ;
      RECT 1016.500000 419.590000 1058.500000 420.410000 ;
      RECT 966.500000 419.590000 1008.500000 420.410000 ;
      RECT 916.500000 419.590000 958.500000 420.410000 ;
      RECT 866.500000 419.590000 908.500000 420.410000 ;
      RECT 816.500000 419.590000 858.500000 420.410000 ;
      RECT 766.500000 419.590000 808.500000 420.410000 ;
      RECT 722.500000 419.590000 758.500000 420.410000 ;
      RECT 666.500000 419.590000 709.500000 420.410000 ;
      RECT 616.500000 419.590000 658.500000 420.410000 ;
      RECT 566.500000 419.590000 608.500000 420.410000 ;
      RECT 516.500000 419.590000 558.500000 420.410000 ;
      RECT 466.500000 419.590000 508.500000 420.410000 ;
      RECT 366.500000 419.590000 408.500000 420.410000 ;
      RECT 316.500000 419.590000 358.500000 420.410000 ;
      RECT 216.500000 419.590000 308.500000 420.410000 ;
      RECT 116.500000 419.590000 208.500000 420.410000 ;
      RECT 66.500000 419.590000 108.500000 420.410000 ;
      RECT 29.500000 419.590000 58.500000 420.410000 ;
      RECT 0.000000 419.590000 16.500000 420.410000 ;
      RECT 416.500000 418.605000 458.500000 420.410000 ;
      RECT 1169.500000 418.410000 1170.500000 419.590000 ;
      RECT 1116.500000 418.410000 1149.500000 419.590000 ;
      RECT 1107.500000 418.410000 1108.500000 419.590000 ;
      RECT 1066.500000 418.410000 1099.500000 419.590000 ;
      RECT 1057.500000 418.410000 1058.500000 419.590000 ;
      RECT 1016.500000 418.410000 1049.500000 419.590000 ;
      RECT 1007.500000 418.410000 1008.500000 419.590000 ;
      RECT 966.500000 418.410000 999.500000 419.590000 ;
      RECT 957.500000 418.410000 958.500000 419.590000 ;
      RECT 916.500000 418.410000 949.500000 419.590000 ;
      RECT 907.500000 418.410000 908.500000 419.590000 ;
      RECT 866.500000 418.410000 899.500000 419.590000 ;
      RECT 857.500000 418.410000 858.500000 419.590000 ;
      RECT 816.500000 418.410000 849.500000 419.590000 ;
      RECT 807.500000 418.410000 808.500000 419.590000 ;
      RECT 766.500000 418.410000 799.500000 419.590000 ;
      RECT 757.500000 418.410000 758.500000 419.590000 ;
      RECT 722.500000 418.410000 749.500000 419.590000 ;
      RECT 707.500000 418.410000 709.500000 419.590000 ;
      RECT 666.500000 418.410000 699.500000 419.590000 ;
      RECT 657.500000 418.410000 658.500000 419.590000 ;
      RECT 616.500000 418.410000 649.500000 419.590000 ;
      RECT 607.500000 418.410000 608.500000 419.590000 ;
      RECT 566.500000 418.410000 599.500000 419.590000 ;
      RECT 557.500000 418.410000 558.500000 419.590000 ;
      RECT 516.500000 418.410000 549.500000 419.590000 ;
      RECT 507.500000 418.410000 508.500000 419.590000 ;
      RECT 466.500000 418.410000 499.500000 419.590000 ;
      RECT 457.500000 418.410000 458.500000 418.605000 ;
      RECT 416.500000 418.410000 449.500000 418.605000 ;
      RECT 407.500000 418.410000 408.500000 419.590000 ;
      RECT 366.500000 418.410000 399.500000 419.590000 ;
      RECT 357.500000 418.410000 358.500000 419.590000 ;
      RECT 316.500000 418.410000 349.500000 419.590000 ;
      RECT 307.500000 418.410000 308.500000 419.590000 ;
      RECT 216.500000 418.410000 299.500000 419.590000 ;
      RECT 207.500000 418.410000 208.500000 419.590000 ;
      RECT 116.500000 418.410000 199.500000 419.590000 ;
      RECT 107.500000 418.410000 108.500000 419.590000 ;
      RECT 66.500000 418.410000 99.500000 419.590000 ;
      RECT 57.500000 418.410000 58.500000 419.590000 ;
      RECT 29.500000 418.410000 49.500000 419.590000 ;
      RECT 15.500000 418.410000 16.500000 419.590000 ;
      RECT 1157.500000 417.590000 1170.500000 418.410000 ;
      RECT 1107.500000 417.590000 1149.500000 418.410000 ;
      RECT 1057.500000 417.590000 1099.500000 418.410000 ;
      RECT 1007.500000 417.590000 1049.500000 418.410000 ;
      RECT 957.500000 417.590000 999.500000 418.410000 ;
      RECT 907.500000 417.590000 949.500000 418.410000 ;
      RECT 857.500000 417.590000 899.500000 418.410000 ;
      RECT 807.500000 417.590000 849.500000 418.410000 ;
      RECT 757.500000 417.590000 799.500000 418.410000 ;
      RECT 707.500000 417.590000 749.500000 418.410000 ;
      RECT 657.500000 417.590000 699.500000 418.410000 ;
      RECT 607.500000 417.590000 649.500000 418.410000 ;
      RECT 557.500000 417.590000 599.500000 418.410000 ;
      RECT 507.500000 417.590000 549.500000 418.410000 ;
      RECT 407.500000 417.590000 449.500000 418.410000 ;
      RECT 357.500000 417.590000 399.500000 418.410000 ;
      RECT 307.500000 417.590000 349.500000 418.410000 ;
      RECT 207.500000 417.590000 299.500000 418.410000 ;
      RECT 107.500000 417.590000 199.500000 418.410000 ;
      RECT 57.500000 417.590000 99.500000 418.410000 ;
      RECT 15.500000 417.590000 49.500000 418.410000 ;
      RECT 1183.500000 416.410000 1186.000000 419.590000 ;
      RECT 1169.500000 416.410000 1170.500000 417.590000 ;
      RECT 1116.500000 416.410000 1149.500000 417.590000 ;
      RECT 1107.500000 416.410000 1108.500000 417.590000 ;
      RECT 1066.500000 416.410000 1099.500000 417.590000 ;
      RECT 1057.500000 416.410000 1058.500000 417.590000 ;
      RECT 1016.500000 416.410000 1049.500000 417.590000 ;
      RECT 1007.500000 416.410000 1008.500000 417.590000 ;
      RECT 966.500000 416.410000 999.500000 417.590000 ;
      RECT 957.500000 416.410000 958.500000 417.590000 ;
      RECT 916.500000 416.410000 949.500000 417.590000 ;
      RECT 907.500000 416.410000 908.500000 417.590000 ;
      RECT 866.500000 416.410000 899.500000 417.590000 ;
      RECT 857.500000 416.410000 858.500000 417.590000 ;
      RECT 816.500000 416.410000 849.500000 417.590000 ;
      RECT 807.500000 416.410000 808.500000 417.590000 ;
      RECT 766.500000 416.410000 799.500000 417.590000 ;
      RECT 757.500000 416.410000 758.500000 417.590000 ;
      RECT 720.000000 416.410000 749.500000 417.590000 ;
      RECT 707.500000 416.410000 712.000000 417.590000 ;
      RECT 666.500000 416.410000 699.500000 417.590000 ;
      RECT 657.500000 416.410000 658.500000 417.590000 ;
      RECT 616.500000 416.410000 649.500000 417.590000 ;
      RECT 607.500000 416.410000 608.500000 417.590000 ;
      RECT 566.500000 416.410000 599.500000 417.590000 ;
      RECT 557.500000 416.410000 558.500000 417.590000 ;
      RECT 516.500000 416.410000 549.500000 417.590000 ;
      RECT 507.500000 416.410000 508.500000 417.590000 ;
      RECT 457.500000 416.410000 499.500000 418.410000 ;
      RECT 407.500000 416.410000 408.500000 417.590000 ;
      RECT 366.500000 416.410000 399.500000 417.590000 ;
      RECT 357.500000 416.410000 358.500000 417.590000 ;
      RECT 316.500000 416.410000 349.500000 417.590000 ;
      RECT 307.500000 416.410000 308.500000 417.590000 ;
      RECT 216.500000 416.410000 299.500000 417.590000 ;
      RECT 207.500000 416.410000 208.500000 417.590000 ;
      RECT 116.500000 416.410000 199.500000 417.590000 ;
      RECT 107.500000 416.410000 108.500000 417.590000 ;
      RECT 66.500000 416.410000 99.500000 417.590000 ;
      RECT 57.500000 416.410000 58.500000 417.590000 ;
      RECT 29.500000 416.410000 49.500000 417.590000 ;
      RECT 15.500000 416.410000 16.500000 417.590000 ;
      RECT 0.000000 416.410000 2.500000 419.590000 ;
      RECT 1169.500000 415.590000 1186.000000 416.410000 ;
      RECT 1116.500000 415.590000 1156.500000 416.410000 ;
      RECT 1066.500000 415.590000 1108.500000 416.410000 ;
      RECT 1016.500000 415.590000 1058.500000 416.410000 ;
      RECT 966.500000 415.590000 1008.500000 416.410000 ;
      RECT 916.500000 415.590000 958.500000 416.410000 ;
      RECT 866.500000 415.590000 908.500000 416.410000 ;
      RECT 816.500000 415.590000 858.500000 416.410000 ;
      RECT 766.500000 415.590000 808.500000 416.410000 ;
      RECT 720.000000 415.590000 758.500000 416.410000 ;
      RECT 666.500000 415.590000 712.000000 416.410000 ;
      RECT 616.500000 415.590000 658.500000 416.410000 ;
      RECT 566.500000 415.590000 608.500000 416.410000 ;
      RECT 516.500000 415.590000 558.500000 416.410000 ;
      RECT 457.500000 415.590000 508.500000 416.410000 ;
      RECT 366.500000 415.590000 408.500000 416.410000 ;
      RECT 316.500000 415.590000 358.500000 416.410000 ;
      RECT 216.500000 415.590000 308.500000 416.410000 ;
      RECT 116.500000 415.590000 208.500000 416.410000 ;
      RECT 66.500000 415.590000 108.500000 416.410000 ;
      RECT 29.500000 415.590000 58.500000 416.410000 ;
      RECT 0.000000 415.590000 16.500000 416.410000 ;
      RECT 457.500000 414.605000 499.500000 415.590000 ;
      RECT 416.500000 414.605000 449.500000 417.590000 ;
      RECT 1169.500000 414.410000 1170.500000 415.590000 ;
      RECT 1116.500000 414.410000 1149.500000 415.590000 ;
      RECT 1107.500000 414.410000 1108.500000 415.590000 ;
      RECT 1066.500000 414.410000 1099.500000 415.590000 ;
      RECT 1057.500000 414.410000 1058.500000 415.590000 ;
      RECT 1016.500000 414.410000 1049.500000 415.590000 ;
      RECT 1007.500000 414.410000 1008.500000 415.590000 ;
      RECT 966.500000 414.410000 999.500000 415.590000 ;
      RECT 957.500000 414.410000 958.500000 415.590000 ;
      RECT 916.500000 414.410000 949.500000 415.590000 ;
      RECT 907.500000 414.410000 908.500000 415.590000 ;
      RECT 866.500000 414.410000 899.500000 415.590000 ;
      RECT 857.500000 414.410000 858.500000 415.590000 ;
      RECT 816.500000 414.410000 849.500000 415.590000 ;
      RECT 807.500000 414.410000 808.500000 415.590000 ;
      RECT 766.500000 414.410000 799.500000 415.590000 ;
      RECT 757.500000 414.410000 758.500000 415.590000 ;
      RECT 720.000000 414.410000 749.500000 415.590000 ;
      RECT 707.500000 414.410000 712.000000 415.590000 ;
      RECT 666.500000 414.410000 699.500000 415.590000 ;
      RECT 657.500000 414.410000 658.500000 415.590000 ;
      RECT 616.500000 414.410000 649.500000 415.590000 ;
      RECT 607.500000 414.410000 608.500000 415.590000 ;
      RECT 566.500000 414.410000 599.500000 415.590000 ;
      RECT 557.500000 414.410000 558.500000 415.590000 ;
      RECT 516.500000 414.410000 549.500000 415.590000 ;
      RECT 507.500000 414.410000 508.500000 415.590000 ;
      RECT 416.500000 414.410000 499.500000 414.605000 ;
      RECT 407.500000 414.410000 408.500000 415.590000 ;
      RECT 366.500000 414.410000 399.500000 415.590000 ;
      RECT 357.500000 414.410000 358.500000 415.590000 ;
      RECT 316.500000 414.410000 349.500000 415.590000 ;
      RECT 307.500000 414.410000 308.500000 415.590000 ;
      RECT 216.500000 414.410000 299.500000 415.590000 ;
      RECT 207.500000 414.410000 208.500000 415.590000 ;
      RECT 116.500000 414.410000 199.500000 415.590000 ;
      RECT 107.500000 414.410000 108.500000 415.590000 ;
      RECT 66.500000 414.410000 99.500000 415.590000 ;
      RECT 57.500000 414.410000 58.500000 415.590000 ;
      RECT 29.500000 414.410000 49.500000 415.590000 ;
      RECT 15.500000 414.410000 16.500000 415.590000 ;
      RECT 1157.500000 413.590000 1170.500000 414.410000 ;
      RECT 1107.500000 413.590000 1149.500000 414.410000 ;
      RECT 1057.500000 413.590000 1099.500000 414.410000 ;
      RECT 1007.500000 413.590000 1049.500000 414.410000 ;
      RECT 957.500000 413.590000 999.500000 414.410000 ;
      RECT 907.500000 413.590000 949.500000 414.410000 ;
      RECT 857.500000 413.590000 899.500000 414.410000 ;
      RECT 807.500000 413.590000 849.500000 414.410000 ;
      RECT 757.500000 413.590000 799.500000 414.410000 ;
      RECT 707.500000 413.590000 749.500000 414.410000 ;
      RECT 657.500000 413.590000 699.500000 414.410000 ;
      RECT 607.500000 413.590000 649.500000 414.410000 ;
      RECT 557.500000 413.590000 599.500000 414.410000 ;
      RECT 507.500000 413.590000 549.500000 414.410000 ;
      RECT 407.500000 413.590000 499.500000 414.410000 ;
      RECT 357.500000 413.590000 399.500000 414.410000 ;
      RECT 307.500000 413.590000 349.500000 414.410000 ;
      RECT 207.500000 413.590000 299.500000 414.410000 ;
      RECT 107.500000 413.590000 199.500000 414.410000 ;
      RECT 57.500000 413.590000 99.500000 414.410000 ;
      RECT 15.500000 413.590000 49.500000 414.410000 ;
      RECT 1183.500000 412.410000 1186.000000 415.590000 ;
      RECT 1169.500000 412.410000 1170.500000 413.590000 ;
      RECT 1116.500000 412.410000 1149.500000 413.590000 ;
      RECT 1107.500000 412.410000 1108.500000 413.590000 ;
      RECT 1066.500000 412.410000 1099.500000 413.590000 ;
      RECT 1057.500000 412.410000 1058.500000 413.590000 ;
      RECT 1016.500000 412.410000 1049.500000 413.590000 ;
      RECT 1007.500000 412.410000 1008.500000 413.590000 ;
      RECT 966.500000 412.410000 999.500000 413.590000 ;
      RECT 957.500000 412.410000 958.500000 413.590000 ;
      RECT 916.500000 412.410000 949.500000 413.590000 ;
      RECT 907.500000 412.410000 908.500000 413.590000 ;
      RECT 866.500000 412.410000 899.500000 413.590000 ;
      RECT 857.500000 412.410000 858.500000 413.590000 ;
      RECT 816.500000 412.410000 849.500000 413.590000 ;
      RECT 807.500000 412.410000 808.500000 413.590000 ;
      RECT 766.500000 412.410000 799.500000 413.590000 ;
      RECT 757.500000 412.410000 758.500000 413.590000 ;
      RECT 720.000000 412.410000 749.500000 413.590000 ;
      RECT 707.500000 412.410000 708.500000 413.590000 ;
      RECT 666.500000 412.410000 699.500000 413.590000 ;
      RECT 657.500000 412.410000 658.500000 413.590000 ;
      RECT 616.500000 412.410000 649.500000 413.590000 ;
      RECT 607.500000 412.410000 608.500000 413.590000 ;
      RECT 566.500000 412.410000 599.500000 413.590000 ;
      RECT 557.500000 412.410000 558.500000 413.590000 ;
      RECT 516.500000 412.410000 549.500000 413.590000 ;
      RECT 507.500000 412.410000 508.500000 413.590000 ;
      RECT 416.500000 412.410000 499.500000 413.590000 ;
      RECT 407.500000 412.410000 408.500000 413.590000 ;
      RECT 366.500000 412.410000 399.500000 413.590000 ;
      RECT 357.500000 412.410000 358.500000 413.590000 ;
      RECT 316.500000 412.410000 349.500000 413.590000 ;
      RECT 307.500000 412.410000 308.500000 413.590000 ;
      RECT 216.500000 412.410000 299.500000 413.590000 ;
      RECT 207.500000 412.410000 208.500000 413.590000 ;
      RECT 116.500000 412.410000 199.500000 413.590000 ;
      RECT 107.500000 412.410000 108.500000 413.590000 ;
      RECT 66.500000 412.410000 99.500000 413.590000 ;
      RECT 57.500000 412.410000 58.500000 413.590000 ;
      RECT 29.500000 412.410000 49.500000 413.590000 ;
      RECT 15.500000 412.410000 16.500000 413.590000 ;
      RECT 0.000000 412.410000 2.500000 415.590000 ;
      RECT 1169.500000 411.590000 1186.000000 412.410000 ;
      RECT 1116.500000 411.590000 1156.500000 412.410000 ;
      RECT 1066.500000 411.590000 1108.500000 412.410000 ;
      RECT 1016.500000 411.590000 1058.500000 412.410000 ;
      RECT 966.500000 411.590000 1008.500000 412.410000 ;
      RECT 916.500000 411.590000 958.500000 412.410000 ;
      RECT 866.500000 411.590000 908.500000 412.410000 ;
      RECT 816.500000 411.590000 858.500000 412.410000 ;
      RECT 766.500000 411.590000 808.500000 412.410000 ;
      RECT 720.000000 411.590000 758.500000 412.410000 ;
      RECT 666.500000 411.590000 708.500000 412.410000 ;
      RECT 616.500000 411.590000 658.500000 412.410000 ;
      RECT 566.500000 411.590000 608.500000 412.410000 ;
      RECT 516.500000 411.590000 558.500000 412.410000 ;
      RECT 416.500000 411.590000 508.500000 412.410000 ;
      RECT 366.500000 411.590000 408.500000 412.410000 ;
      RECT 316.500000 411.590000 358.500000 412.410000 ;
      RECT 216.500000 411.590000 308.500000 412.410000 ;
      RECT 116.500000 411.590000 208.500000 412.410000 ;
      RECT 66.500000 411.590000 108.500000 412.410000 ;
      RECT 29.500000 411.590000 58.500000 412.410000 ;
      RECT 0.000000 411.590000 16.500000 412.410000 ;
      RECT 1169.500000 410.410000 1170.500000 411.590000 ;
      RECT 1116.500000 410.410000 1149.500000 411.590000 ;
      RECT 1107.500000 410.410000 1108.500000 411.590000 ;
      RECT 1066.500000 410.410000 1099.500000 411.590000 ;
      RECT 1057.500000 410.410000 1058.500000 411.590000 ;
      RECT 1016.500000 410.410000 1049.500000 411.590000 ;
      RECT 1007.500000 410.410000 1008.500000 411.590000 ;
      RECT 966.500000 410.410000 999.500000 411.590000 ;
      RECT 957.500000 410.410000 958.500000 411.590000 ;
      RECT 916.500000 410.410000 949.500000 411.590000 ;
      RECT 907.500000 410.410000 908.500000 411.590000 ;
      RECT 866.500000 410.410000 899.500000 411.590000 ;
      RECT 857.500000 410.410000 858.500000 411.590000 ;
      RECT 816.500000 410.410000 849.500000 411.590000 ;
      RECT 807.500000 410.410000 808.500000 411.590000 ;
      RECT 766.500000 410.410000 799.500000 411.590000 ;
      RECT 757.500000 410.410000 758.500000 411.590000 ;
      RECT 720.000000 410.410000 749.500000 411.590000 ;
      RECT 707.500000 410.410000 708.500000 411.590000 ;
      RECT 666.500000 410.410000 699.500000 411.590000 ;
      RECT 657.500000 410.410000 658.500000 411.590000 ;
      RECT 616.500000 410.410000 649.500000 411.590000 ;
      RECT 607.500000 410.410000 608.500000 411.590000 ;
      RECT 566.500000 410.410000 599.500000 411.590000 ;
      RECT 557.500000 410.410000 558.500000 411.590000 ;
      RECT 516.500000 410.410000 549.500000 411.590000 ;
      RECT 507.500000 410.410000 508.500000 411.590000 ;
      RECT 416.500000 410.410000 499.500000 411.590000 ;
      RECT 407.500000 410.410000 408.500000 411.590000 ;
      RECT 366.500000 410.410000 399.500000 411.590000 ;
      RECT 357.500000 410.410000 358.500000 411.590000 ;
      RECT 316.500000 410.410000 349.500000 411.590000 ;
      RECT 307.500000 410.410000 308.500000 411.590000 ;
      RECT 216.500000 410.410000 299.500000 411.590000 ;
      RECT 207.500000 410.410000 208.500000 411.590000 ;
      RECT 116.500000 410.410000 199.500000 411.590000 ;
      RECT 107.500000 410.410000 108.500000 411.590000 ;
      RECT 66.500000 410.410000 99.500000 411.590000 ;
      RECT 57.500000 410.410000 58.500000 411.590000 ;
      RECT 29.500000 410.410000 49.500000 411.590000 ;
      RECT 15.500000 410.410000 16.500000 411.590000 ;
      RECT 1157.500000 409.590000 1170.500000 410.410000 ;
      RECT 1107.500000 409.590000 1149.500000 410.410000 ;
      RECT 1057.500000 409.590000 1099.500000 410.410000 ;
      RECT 1007.500000 409.590000 1049.500000 410.410000 ;
      RECT 957.500000 409.590000 999.500000 410.410000 ;
      RECT 907.500000 409.590000 949.500000 410.410000 ;
      RECT 857.500000 409.590000 899.500000 410.410000 ;
      RECT 807.500000 409.590000 849.500000 410.410000 ;
      RECT 757.500000 409.590000 799.500000 410.410000 ;
      RECT 707.500000 409.590000 749.500000 410.410000 ;
      RECT 657.500000 409.590000 699.500000 410.410000 ;
      RECT 607.500000 409.590000 649.500000 410.410000 ;
      RECT 557.500000 409.590000 599.500000 410.410000 ;
      RECT 507.500000 409.590000 549.500000 410.410000 ;
      RECT 407.500000 409.590000 499.500000 410.410000 ;
      RECT 357.500000 409.590000 399.500000 410.410000 ;
      RECT 307.500000 409.590000 349.500000 410.410000 ;
      RECT 207.500000 409.590000 299.500000 410.410000 ;
      RECT 107.500000 409.590000 199.500000 410.410000 ;
      RECT 57.500000 409.590000 99.500000 410.410000 ;
      RECT 15.500000 409.590000 49.500000 410.410000 ;
      RECT 1183.500000 408.410000 1186.000000 411.590000 ;
      RECT 1169.500000 408.410000 1170.500000 409.590000 ;
      RECT 1116.500000 408.410000 1149.500000 409.590000 ;
      RECT 1107.500000 408.410000 1108.500000 409.590000 ;
      RECT 1066.500000 408.410000 1099.500000 409.590000 ;
      RECT 1057.500000 408.410000 1058.500000 409.590000 ;
      RECT 1016.500000 408.410000 1049.500000 409.590000 ;
      RECT 1007.500000 408.410000 1008.500000 409.590000 ;
      RECT 966.500000 408.410000 999.500000 409.590000 ;
      RECT 957.500000 408.410000 958.500000 409.590000 ;
      RECT 916.500000 408.410000 949.500000 409.590000 ;
      RECT 907.500000 408.410000 908.500000 409.590000 ;
      RECT 866.500000 408.410000 899.500000 409.590000 ;
      RECT 857.500000 408.410000 858.500000 409.590000 ;
      RECT 816.500000 408.410000 849.500000 409.590000 ;
      RECT 807.500000 408.410000 808.500000 409.590000 ;
      RECT 766.500000 408.410000 799.500000 409.590000 ;
      RECT 757.500000 408.410000 758.500000 409.590000 ;
      RECT 716.500000 408.410000 749.500000 409.590000 ;
      RECT 707.500000 408.410000 708.500000 409.590000 ;
      RECT 666.500000 408.410000 699.500000 409.590000 ;
      RECT 657.500000 408.410000 658.500000 409.590000 ;
      RECT 616.500000 408.410000 649.500000 409.590000 ;
      RECT 607.500000 408.410000 608.500000 409.590000 ;
      RECT 566.500000 408.410000 599.500000 409.590000 ;
      RECT 557.500000 408.410000 558.500000 409.590000 ;
      RECT 516.500000 408.410000 549.500000 409.590000 ;
      RECT 507.500000 408.410000 508.500000 409.590000 ;
      RECT 416.500000 408.410000 499.500000 409.590000 ;
      RECT 407.500000 408.410000 408.500000 409.590000 ;
      RECT 366.500000 408.410000 399.500000 409.590000 ;
      RECT 357.500000 408.410000 358.500000 409.590000 ;
      RECT 316.500000 408.410000 349.500000 409.590000 ;
      RECT 307.500000 408.410000 308.500000 409.590000 ;
      RECT 266.500000 408.410000 299.500000 409.590000 ;
      RECT 207.500000 408.410000 208.500000 409.590000 ;
      RECT 166.500000 408.410000 199.500000 409.590000 ;
      RECT 107.500000 408.410000 108.500000 409.590000 ;
      RECT 66.500000 408.410000 99.500000 409.590000 ;
      RECT 57.500000 408.410000 58.500000 409.590000 ;
      RECT 29.500000 408.410000 49.500000 409.590000 ;
      RECT 15.500000 408.410000 16.500000 409.590000 ;
      RECT 0.000000 408.410000 2.500000 411.590000 ;
      RECT 1169.500000 407.590000 1186.000000 408.410000 ;
      RECT 1116.500000 407.590000 1156.500000 408.410000 ;
      RECT 1066.500000 407.590000 1108.500000 408.410000 ;
      RECT 1016.500000 407.590000 1058.500000 408.410000 ;
      RECT 966.500000 407.590000 1008.500000 408.410000 ;
      RECT 916.500000 407.590000 958.500000 408.410000 ;
      RECT 866.500000 407.590000 908.500000 408.410000 ;
      RECT 816.500000 407.590000 858.500000 408.410000 ;
      RECT 766.500000 407.590000 808.500000 408.410000 ;
      RECT 716.500000 407.590000 758.500000 408.410000 ;
      RECT 666.500000 407.590000 708.500000 408.410000 ;
      RECT 616.500000 407.590000 658.500000 408.410000 ;
      RECT 566.500000 407.590000 608.500000 408.410000 ;
      RECT 516.500000 407.590000 558.500000 408.410000 ;
      RECT 416.500000 407.590000 508.500000 408.410000 ;
      RECT 366.500000 407.590000 408.500000 408.410000 ;
      RECT 316.500000 407.590000 358.500000 408.410000 ;
      RECT 266.500000 407.590000 308.500000 408.410000 ;
      RECT 216.500000 407.590000 258.500000 409.590000 ;
      RECT 166.500000 407.590000 208.500000 408.410000 ;
      RECT 116.500000 407.590000 158.500000 409.590000 ;
      RECT 66.500000 407.590000 108.500000 408.410000 ;
      RECT 29.500000 407.590000 58.500000 408.410000 ;
      RECT 0.000000 407.590000 16.500000 408.410000 ;
      RECT 1169.500000 406.410000 1170.500000 407.590000 ;
      RECT 1116.500000 406.410000 1149.500000 407.590000 ;
      RECT 1107.500000 406.410000 1108.500000 407.590000 ;
      RECT 1066.500000 406.410000 1099.500000 407.590000 ;
      RECT 1057.500000 406.410000 1058.500000 407.590000 ;
      RECT 1016.500000 406.410000 1049.500000 407.590000 ;
      RECT 1007.500000 406.410000 1008.500000 407.590000 ;
      RECT 966.500000 406.410000 999.500000 407.590000 ;
      RECT 957.500000 406.410000 958.500000 407.590000 ;
      RECT 916.500000 406.410000 949.500000 407.590000 ;
      RECT 907.500000 406.410000 908.500000 407.590000 ;
      RECT 866.500000 406.410000 899.500000 407.590000 ;
      RECT 857.500000 406.410000 858.500000 407.590000 ;
      RECT 816.500000 406.410000 849.500000 407.590000 ;
      RECT 807.500000 406.410000 808.500000 407.590000 ;
      RECT 766.500000 406.410000 799.500000 407.590000 ;
      RECT 757.500000 406.410000 758.500000 407.590000 ;
      RECT 716.500000 406.410000 749.500000 407.590000 ;
      RECT 707.500000 406.410000 708.500000 407.590000 ;
      RECT 666.500000 406.410000 699.500000 407.590000 ;
      RECT 657.500000 406.410000 658.500000 407.590000 ;
      RECT 616.500000 406.410000 649.500000 407.590000 ;
      RECT 607.500000 406.410000 608.500000 407.590000 ;
      RECT 566.500000 406.410000 599.500000 407.590000 ;
      RECT 557.500000 406.410000 558.500000 407.590000 ;
      RECT 516.500000 406.410000 549.500000 407.590000 ;
      RECT 507.500000 406.410000 508.500000 407.590000 ;
      RECT 416.500000 406.410000 499.500000 407.590000 ;
      RECT 407.500000 406.410000 408.500000 407.590000 ;
      RECT 366.500000 406.410000 399.500000 407.590000 ;
      RECT 357.500000 406.410000 358.500000 407.590000 ;
      RECT 316.500000 406.410000 349.500000 407.590000 ;
      RECT 307.500000 406.410000 308.500000 407.590000 ;
      RECT 266.500000 406.410000 299.500000 407.590000 ;
      RECT 257.500000 406.410000 258.500000 407.590000 ;
      RECT 216.500000 406.410000 249.500000 407.590000 ;
      RECT 207.500000 406.410000 208.500000 407.590000 ;
      RECT 166.500000 406.410000 199.500000 407.590000 ;
      RECT 157.500000 406.410000 158.500000 407.590000 ;
      RECT 116.500000 406.410000 149.500000 407.590000 ;
      RECT 107.500000 406.410000 108.500000 407.590000 ;
      RECT 66.500000 406.410000 99.500000 407.590000 ;
      RECT 57.500000 406.410000 58.500000 407.590000 ;
      RECT 29.500000 406.410000 49.500000 407.590000 ;
      RECT 15.500000 406.410000 16.500000 407.590000 ;
      RECT 1157.500000 405.590000 1170.500000 406.410000 ;
      RECT 1107.500000 405.590000 1149.500000 406.410000 ;
      RECT 1057.500000 405.590000 1099.500000 406.410000 ;
      RECT 1007.500000 405.590000 1049.500000 406.410000 ;
      RECT 957.500000 405.590000 999.500000 406.410000 ;
      RECT 907.500000 405.590000 949.500000 406.410000 ;
      RECT 857.500000 405.590000 899.500000 406.410000 ;
      RECT 807.500000 405.590000 849.500000 406.410000 ;
      RECT 757.500000 405.590000 799.500000 406.410000 ;
      RECT 707.500000 405.590000 749.500000 406.410000 ;
      RECT 657.500000 405.590000 699.500000 406.410000 ;
      RECT 607.500000 405.590000 649.500000 406.410000 ;
      RECT 557.500000 405.590000 599.500000 406.410000 ;
      RECT 507.500000 405.590000 549.500000 406.410000 ;
      RECT 407.500000 405.590000 499.500000 406.410000 ;
      RECT 357.500000 405.590000 399.500000 406.410000 ;
      RECT 307.500000 405.590000 349.500000 406.410000 ;
      RECT 257.500000 405.590000 299.500000 406.410000 ;
      RECT 207.500000 405.590000 249.500000 406.410000 ;
      RECT 157.500000 405.590000 199.500000 406.410000 ;
      RECT 107.500000 405.590000 149.500000 406.410000 ;
      RECT 57.500000 405.590000 99.500000 406.410000 ;
      RECT 15.500000 405.590000 49.500000 406.410000 ;
      RECT 1183.500000 404.410000 1186.000000 407.590000 ;
      RECT 1169.500000 404.410000 1170.500000 405.590000 ;
      RECT 1116.500000 404.410000 1149.500000 405.590000 ;
      RECT 1107.500000 404.410000 1108.500000 405.590000 ;
      RECT 1066.500000 404.410000 1099.500000 405.590000 ;
      RECT 1057.500000 404.410000 1058.500000 405.590000 ;
      RECT 1016.500000 404.410000 1049.500000 405.590000 ;
      RECT 1007.500000 404.410000 1008.500000 405.590000 ;
      RECT 966.500000 404.410000 999.500000 405.590000 ;
      RECT 957.500000 404.410000 958.500000 405.590000 ;
      RECT 916.500000 404.410000 949.500000 405.590000 ;
      RECT 907.500000 404.410000 908.500000 405.590000 ;
      RECT 866.500000 404.410000 899.500000 405.590000 ;
      RECT 857.500000 404.410000 858.500000 405.590000 ;
      RECT 816.500000 404.410000 849.500000 405.590000 ;
      RECT 807.500000 404.410000 808.500000 405.590000 ;
      RECT 766.500000 404.410000 799.500000 405.590000 ;
      RECT 757.500000 404.410000 758.500000 405.590000 ;
      RECT 716.500000 404.410000 749.500000 405.590000 ;
      RECT 707.500000 404.410000 708.500000 405.590000 ;
      RECT 666.500000 404.410000 699.500000 405.590000 ;
      RECT 657.500000 404.410000 658.500000 405.590000 ;
      RECT 616.500000 404.410000 649.500000 405.590000 ;
      RECT 607.500000 404.410000 608.500000 405.590000 ;
      RECT 566.500000 404.410000 599.500000 405.590000 ;
      RECT 557.500000 404.410000 558.500000 405.590000 ;
      RECT 516.500000 404.410000 549.500000 405.590000 ;
      RECT 507.500000 404.410000 508.500000 405.590000 ;
      RECT 416.500000 404.410000 499.500000 405.590000 ;
      RECT 407.500000 404.410000 408.500000 405.590000 ;
      RECT 366.500000 404.410000 399.500000 405.590000 ;
      RECT 357.500000 404.410000 358.500000 405.590000 ;
      RECT 316.500000 404.410000 349.500000 405.590000 ;
      RECT 307.500000 404.410000 308.500000 405.590000 ;
      RECT 266.500000 404.410000 299.500000 405.590000 ;
      RECT 257.500000 404.410000 258.500000 405.590000 ;
      RECT 216.500000 404.410000 249.500000 405.590000 ;
      RECT 207.500000 404.410000 208.500000 405.590000 ;
      RECT 166.500000 404.410000 199.500000 405.590000 ;
      RECT 157.500000 404.410000 158.500000 405.590000 ;
      RECT 116.500000 404.410000 149.500000 405.590000 ;
      RECT 107.500000 404.410000 108.500000 405.590000 ;
      RECT 66.500000 404.410000 99.500000 405.590000 ;
      RECT 57.500000 404.410000 58.500000 405.590000 ;
      RECT 29.500000 404.410000 49.500000 405.590000 ;
      RECT 15.500000 404.410000 16.500000 405.590000 ;
      RECT 0.000000 404.410000 2.500000 407.590000 ;
      RECT 416.500000 403.730000 508.500000 404.410000 ;
      RECT 1169.500000 403.590000 1186.000000 404.410000 ;
      RECT 1116.500000 403.590000 1156.500000 404.410000 ;
      RECT 1066.500000 403.590000 1108.500000 404.410000 ;
      RECT 1016.500000 403.590000 1058.500000 404.410000 ;
      RECT 966.500000 403.590000 1008.500000 404.410000 ;
      RECT 916.500000 403.590000 958.500000 404.410000 ;
      RECT 866.500000 403.590000 908.500000 404.410000 ;
      RECT 816.500000 403.590000 858.500000 404.410000 ;
      RECT 766.500000 403.590000 808.500000 404.410000 ;
      RECT 716.500000 403.590000 758.500000 404.410000 ;
      RECT 666.500000 403.590000 708.500000 404.410000 ;
      RECT 616.500000 403.590000 658.500000 404.410000 ;
      RECT 566.500000 403.590000 608.500000 404.410000 ;
      RECT 516.500000 403.590000 558.500000 404.410000 ;
      RECT 466.500000 403.590000 508.500000 403.730000 ;
      RECT 366.500000 403.590000 408.500000 404.410000 ;
      RECT 316.500000 403.590000 358.500000 404.410000 ;
      RECT 266.500000 403.590000 308.500000 404.410000 ;
      RECT 216.500000 403.590000 258.500000 404.410000 ;
      RECT 166.500000 403.590000 208.500000 404.410000 ;
      RECT 116.500000 403.590000 158.500000 404.410000 ;
      RECT 66.500000 403.590000 108.500000 404.410000 ;
      RECT 29.500000 403.590000 58.500000 404.410000 ;
      RECT 0.000000 403.590000 16.500000 404.410000 ;
      RECT 1169.500000 402.410000 1170.500000 403.590000 ;
      RECT 1116.500000 402.410000 1149.500000 403.590000 ;
      RECT 1107.500000 402.410000 1108.500000 403.590000 ;
      RECT 1066.500000 402.410000 1099.500000 403.590000 ;
      RECT 1057.500000 402.410000 1058.500000 403.590000 ;
      RECT 1016.500000 402.410000 1049.500000 403.590000 ;
      RECT 1007.500000 402.410000 1008.500000 403.590000 ;
      RECT 966.500000 402.410000 999.500000 403.590000 ;
      RECT 957.500000 402.410000 958.500000 403.590000 ;
      RECT 916.500000 402.410000 949.500000 403.590000 ;
      RECT 907.500000 402.410000 908.500000 403.590000 ;
      RECT 866.500000 402.410000 899.500000 403.590000 ;
      RECT 857.500000 402.410000 858.500000 403.590000 ;
      RECT 816.500000 402.410000 849.500000 403.590000 ;
      RECT 807.500000 402.410000 808.500000 403.590000 ;
      RECT 766.500000 402.410000 799.500000 403.590000 ;
      RECT 757.500000 402.410000 758.500000 403.590000 ;
      RECT 716.500000 402.410000 749.500000 403.590000 ;
      RECT 707.500000 402.410000 708.500000 403.590000 ;
      RECT 666.500000 402.410000 699.500000 403.590000 ;
      RECT 657.500000 402.410000 658.500000 403.590000 ;
      RECT 616.500000 402.410000 649.500000 403.590000 ;
      RECT 607.500000 402.410000 608.500000 403.590000 ;
      RECT 566.500000 402.410000 599.500000 403.590000 ;
      RECT 557.500000 402.410000 558.500000 403.590000 ;
      RECT 516.500000 402.410000 549.500000 403.590000 ;
      RECT 507.500000 402.410000 508.500000 403.590000 ;
      RECT 416.500000 402.410000 458.500000 403.730000 ;
      RECT 407.500000 402.410000 408.500000 403.590000 ;
      RECT 366.500000 402.410000 399.500000 403.590000 ;
      RECT 357.500000 402.410000 358.500000 403.590000 ;
      RECT 316.500000 402.410000 349.500000 403.590000 ;
      RECT 307.500000 402.410000 308.500000 403.590000 ;
      RECT 266.500000 402.410000 299.500000 403.590000 ;
      RECT 257.500000 402.410000 258.500000 403.590000 ;
      RECT 216.500000 402.410000 249.500000 403.590000 ;
      RECT 207.500000 402.410000 208.500000 403.590000 ;
      RECT 166.500000 402.410000 199.500000 403.590000 ;
      RECT 157.500000 402.410000 158.500000 403.590000 ;
      RECT 116.500000 402.410000 149.500000 403.590000 ;
      RECT 107.500000 402.410000 108.500000 403.590000 ;
      RECT 66.500000 402.410000 99.500000 403.590000 ;
      RECT 57.500000 402.410000 58.500000 403.590000 ;
      RECT 29.500000 402.410000 49.500000 403.590000 ;
      RECT 15.500000 402.410000 16.500000 403.590000 ;
      RECT 1157.500000 401.590000 1170.500000 402.410000 ;
      RECT 1107.500000 401.590000 1149.500000 402.410000 ;
      RECT 1057.500000 401.590000 1099.500000 402.410000 ;
      RECT 1007.500000 401.590000 1049.500000 402.410000 ;
      RECT 957.500000 401.590000 999.500000 402.410000 ;
      RECT 907.500000 401.590000 949.500000 402.410000 ;
      RECT 857.500000 401.590000 899.500000 402.410000 ;
      RECT 807.500000 401.590000 849.500000 402.410000 ;
      RECT 757.500000 401.590000 799.500000 402.410000 ;
      RECT 707.500000 401.590000 749.500000 402.410000 ;
      RECT 657.500000 401.590000 699.500000 402.410000 ;
      RECT 607.500000 401.590000 649.500000 402.410000 ;
      RECT 557.500000 401.590000 599.500000 402.410000 ;
      RECT 507.500000 401.590000 549.500000 402.410000 ;
      RECT 407.500000 401.590000 458.500000 402.410000 ;
      RECT 357.500000 401.590000 399.500000 402.410000 ;
      RECT 307.500000 401.590000 349.500000 402.410000 ;
      RECT 257.500000 401.590000 299.500000 402.410000 ;
      RECT 207.500000 401.590000 249.500000 402.410000 ;
      RECT 157.500000 401.590000 199.500000 402.410000 ;
      RECT 107.500000 401.590000 149.500000 402.410000 ;
      RECT 57.500000 401.590000 99.500000 402.410000 ;
      RECT 15.500000 401.590000 49.500000 402.410000 ;
      RECT 1183.500000 400.410000 1186.000000 403.590000 ;
      RECT 1169.500000 400.410000 1170.500000 401.590000 ;
      RECT 1116.500000 400.410000 1149.500000 401.590000 ;
      RECT 1107.500000 400.410000 1108.500000 401.590000 ;
      RECT 1066.500000 400.410000 1099.500000 401.590000 ;
      RECT 1057.500000 400.410000 1058.500000 401.590000 ;
      RECT 1016.500000 400.410000 1049.500000 401.590000 ;
      RECT 1007.500000 400.410000 1008.500000 401.590000 ;
      RECT 966.500000 400.410000 999.500000 401.590000 ;
      RECT 957.500000 400.410000 958.500000 401.590000 ;
      RECT 916.500000 400.410000 949.500000 401.590000 ;
      RECT 907.500000 400.410000 908.500000 401.590000 ;
      RECT 866.500000 400.410000 899.500000 401.590000 ;
      RECT 857.500000 400.410000 858.500000 401.590000 ;
      RECT 816.500000 400.410000 849.500000 401.590000 ;
      RECT 807.500000 400.410000 808.500000 401.590000 ;
      RECT 766.500000 400.410000 799.500000 401.590000 ;
      RECT 757.500000 400.410000 758.500000 401.590000 ;
      RECT 716.500000 400.410000 749.500000 401.590000 ;
      RECT 707.500000 400.410000 708.500000 401.590000 ;
      RECT 666.500000 400.410000 699.500000 401.590000 ;
      RECT 657.500000 400.410000 658.500000 401.590000 ;
      RECT 616.500000 400.410000 649.500000 401.590000 ;
      RECT 607.500000 400.410000 608.500000 401.590000 ;
      RECT 566.500000 400.410000 599.500000 401.590000 ;
      RECT 557.500000 400.410000 558.500000 401.590000 ;
      RECT 516.500000 400.410000 549.500000 401.590000 ;
      RECT 507.500000 400.410000 508.500000 401.590000 ;
      RECT 466.500000 400.410000 499.500000 403.590000 ;
      RECT 407.500000 400.410000 408.500000 401.590000 ;
      RECT 366.500000 400.410000 399.500000 401.590000 ;
      RECT 357.500000 400.410000 358.500000 401.590000 ;
      RECT 316.500000 400.410000 349.500000 401.590000 ;
      RECT 307.500000 400.410000 308.500000 401.590000 ;
      RECT 266.500000 400.410000 299.500000 401.590000 ;
      RECT 257.500000 400.410000 258.500000 401.590000 ;
      RECT 216.500000 400.410000 249.500000 401.590000 ;
      RECT 207.500000 400.410000 208.500000 401.590000 ;
      RECT 166.500000 400.410000 199.500000 401.590000 ;
      RECT 157.500000 400.410000 158.500000 401.590000 ;
      RECT 116.500000 400.410000 149.500000 401.590000 ;
      RECT 107.500000 400.410000 108.500000 401.590000 ;
      RECT 66.500000 400.410000 99.500000 401.590000 ;
      RECT 57.500000 400.410000 58.500000 401.590000 ;
      RECT 29.500000 400.410000 49.500000 401.590000 ;
      RECT 15.500000 400.410000 16.500000 401.590000 ;
      RECT 0.000000 400.410000 2.500000 403.590000 ;
      RECT 466.500000 399.730000 508.500000 400.410000 ;
      RECT 416.500000 399.730000 458.500000 401.590000 ;
      RECT 1169.500000 399.590000 1186.000000 400.410000 ;
      RECT 1116.500000 399.590000 1156.500000 400.410000 ;
      RECT 1066.500000 399.590000 1108.500000 400.410000 ;
      RECT 1016.500000 399.590000 1058.500000 400.410000 ;
      RECT 966.500000 399.590000 1008.500000 400.410000 ;
      RECT 916.500000 399.590000 958.500000 400.410000 ;
      RECT 866.500000 399.590000 908.500000 400.410000 ;
      RECT 816.500000 399.590000 858.500000 400.410000 ;
      RECT 766.500000 399.590000 808.500000 400.410000 ;
      RECT 716.500000 399.590000 758.500000 400.410000 ;
      RECT 666.500000 399.590000 708.500000 400.410000 ;
      RECT 616.500000 399.590000 658.500000 400.410000 ;
      RECT 566.500000 399.590000 608.500000 400.410000 ;
      RECT 516.500000 399.590000 558.500000 400.410000 ;
      RECT 416.500000 399.590000 508.500000 399.730000 ;
      RECT 366.500000 399.590000 408.500000 400.410000 ;
      RECT 316.500000 399.590000 358.500000 400.410000 ;
      RECT 266.500000 399.590000 308.500000 400.410000 ;
      RECT 216.500000 399.590000 258.500000 400.410000 ;
      RECT 166.500000 399.590000 208.500000 400.410000 ;
      RECT 116.500000 399.590000 158.500000 400.410000 ;
      RECT 66.500000 399.590000 108.500000 400.410000 ;
      RECT 29.500000 399.590000 58.500000 400.410000 ;
      RECT 0.000000 399.590000 16.500000 400.410000 ;
      RECT 1169.500000 398.410000 1170.500000 399.590000 ;
      RECT 1116.500000 398.410000 1149.500000 399.590000 ;
      RECT 1107.500000 398.410000 1108.500000 399.590000 ;
      RECT 1066.500000 398.410000 1099.500000 399.590000 ;
      RECT 1057.500000 398.410000 1058.500000 399.590000 ;
      RECT 1016.500000 398.410000 1049.500000 399.590000 ;
      RECT 1007.500000 398.410000 1008.500000 399.590000 ;
      RECT 966.500000 398.410000 999.500000 399.590000 ;
      RECT 957.500000 398.410000 958.500000 399.590000 ;
      RECT 916.500000 398.410000 949.500000 399.590000 ;
      RECT 907.500000 398.410000 908.500000 399.590000 ;
      RECT 866.500000 398.410000 899.500000 399.590000 ;
      RECT 857.500000 398.410000 858.500000 399.590000 ;
      RECT 816.500000 398.410000 849.500000 399.590000 ;
      RECT 807.500000 398.410000 808.500000 399.590000 ;
      RECT 766.500000 398.410000 799.500000 399.590000 ;
      RECT 757.500000 398.410000 758.500000 399.590000 ;
      RECT 716.500000 398.410000 749.500000 399.590000 ;
      RECT 707.500000 398.410000 708.500000 399.590000 ;
      RECT 666.500000 398.410000 699.500000 399.590000 ;
      RECT 657.500000 398.410000 658.500000 399.590000 ;
      RECT 616.500000 398.410000 649.500000 399.590000 ;
      RECT 607.500000 398.410000 608.500000 399.590000 ;
      RECT 566.500000 398.410000 599.500000 399.590000 ;
      RECT 557.500000 398.410000 558.500000 399.590000 ;
      RECT 516.500000 398.410000 549.500000 399.590000 ;
      RECT 507.500000 398.410000 508.500000 399.590000 ;
      RECT 416.500000 398.410000 449.500000 399.590000 ;
      RECT 407.500000 398.410000 408.500000 399.590000 ;
      RECT 366.500000 398.410000 399.500000 399.590000 ;
      RECT 357.500000 398.410000 358.500000 399.590000 ;
      RECT 316.500000 398.410000 349.500000 399.590000 ;
      RECT 307.500000 398.410000 308.500000 399.590000 ;
      RECT 266.500000 398.410000 299.500000 399.590000 ;
      RECT 257.500000 398.410000 258.500000 399.590000 ;
      RECT 216.500000 398.410000 249.500000 399.590000 ;
      RECT 207.500000 398.410000 208.500000 399.590000 ;
      RECT 166.500000 398.410000 199.500000 399.590000 ;
      RECT 157.500000 398.410000 158.500000 399.590000 ;
      RECT 116.500000 398.410000 149.500000 399.590000 ;
      RECT 107.500000 398.410000 108.500000 399.590000 ;
      RECT 66.500000 398.410000 99.500000 399.590000 ;
      RECT 57.500000 398.410000 58.500000 399.590000 ;
      RECT 29.500000 398.410000 49.500000 399.590000 ;
      RECT 15.500000 398.410000 16.500000 399.590000 ;
      RECT 1157.500000 397.590000 1170.500000 398.410000 ;
      RECT 1107.500000 397.590000 1149.500000 398.410000 ;
      RECT 1057.500000 397.590000 1099.500000 398.410000 ;
      RECT 1007.500000 397.590000 1049.500000 398.410000 ;
      RECT 957.500000 397.590000 999.500000 398.410000 ;
      RECT 907.500000 397.590000 949.500000 398.410000 ;
      RECT 857.500000 397.590000 899.500000 398.410000 ;
      RECT 807.500000 397.590000 849.500000 398.410000 ;
      RECT 757.500000 397.590000 799.500000 398.410000 ;
      RECT 707.500000 397.590000 749.500000 398.410000 ;
      RECT 657.500000 397.590000 699.500000 398.410000 ;
      RECT 607.500000 397.590000 649.500000 398.410000 ;
      RECT 557.500000 397.590000 599.500000 398.410000 ;
      RECT 507.500000 397.590000 549.500000 398.410000 ;
      RECT 457.500000 397.590000 499.500000 399.590000 ;
      RECT 407.500000 397.590000 449.500000 398.410000 ;
      RECT 357.500000 397.590000 399.500000 398.410000 ;
      RECT 307.500000 397.590000 349.500000 398.410000 ;
      RECT 257.500000 397.590000 299.500000 398.410000 ;
      RECT 207.500000 397.590000 249.500000 398.410000 ;
      RECT 157.500000 397.590000 199.500000 398.410000 ;
      RECT 107.500000 397.590000 149.500000 398.410000 ;
      RECT 57.500000 397.590000 99.500000 398.410000 ;
      RECT 15.500000 397.590000 49.500000 398.410000 ;
      RECT 1183.500000 396.410000 1186.000000 399.590000 ;
      RECT 1169.500000 396.410000 1170.500000 397.590000 ;
      RECT 1116.500000 396.410000 1149.500000 397.590000 ;
      RECT 1107.500000 396.410000 1108.500000 397.590000 ;
      RECT 1066.500000 396.410000 1099.500000 397.590000 ;
      RECT 1057.500000 396.410000 1058.500000 397.590000 ;
      RECT 1016.500000 396.410000 1049.500000 397.590000 ;
      RECT 1007.500000 396.410000 1008.500000 397.590000 ;
      RECT 966.500000 396.410000 999.500000 397.590000 ;
      RECT 957.500000 396.410000 958.500000 397.590000 ;
      RECT 916.500000 396.410000 949.500000 397.590000 ;
      RECT 907.500000 396.410000 908.500000 397.590000 ;
      RECT 866.500000 396.410000 899.500000 397.590000 ;
      RECT 857.500000 396.410000 858.500000 397.590000 ;
      RECT 816.500000 396.410000 849.500000 397.590000 ;
      RECT 807.500000 396.410000 808.500000 397.590000 ;
      RECT 766.500000 396.410000 799.500000 397.590000 ;
      RECT 757.500000 396.410000 758.500000 397.590000 ;
      RECT 716.500000 396.410000 749.500000 397.590000 ;
      RECT 707.500000 396.410000 708.500000 397.590000 ;
      RECT 666.500000 396.410000 699.500000 397.590000 ;
      RECT 657.500000 396.410000 658.500000 397.590000 ;
      RECT 616.500000 396.410000 649.500000 397.590000 ;
      RECT 607.500000 396.410000 608.500000 397.590000 ;
      RECT 566.500000 396.410000 599.500000 397.590000 ;
      RECT 557.500000 396.410000 558.500000 397.590000 ;
      RECT 516.500000 396.410000 549.500000 397.590000 ;
      RECT 507.500000 396.410000 508.500000 397.590000 ;
      RECT 466.500000 396.410000 499.500000 397.590000 ;
      RECT 457.500000 396.410000 458.500000 397.590000 ;
      RECT 416.500000 396.410000 449.500000 397.590000 ;
      RECT 407.500000 396.410000 408.500000 397.590000 ;
      RECT 366.500000 396.410000 399.500000 397.590000 ;
      RECT 357.500000 396.410000 358.500000 397.590000 ;
      RECT 316.500000 396.410000 349.500000 397.590000 ;
      RECT 307.500000 396.410000 308.500000 397.590000 ;
      RECT 266.500000 396.410000 299.500000 397.590000 ;
      RECT 257.500000 396.410000 258.500000 397.590000 ;
      RECT 216.500000 396.410000 249.500000 397.590000 ;
      RECT 207.500000 396.410000 208.500000 397.590000 ;
      RECT 166.500000 396.410000 199.500000 397.590000 ;
      RECT 157.500000 396.410000 158.500000 397.590000 ;
      RECT 116.500000 396.410000 149.500000 397.590000 ;
      RECT 107.500000 396.410000 108.500000 397.590000 ;
      RECT 66.500000 396.410000 99.500000 397.590000 ;
      RECT 57.500000 396.410000 58.500000 397.590000 ;
      RECT 29.500000 396.410000 49.500000 397.590000 ;
      RECT 15.500000 396.410000 16.500000 397.590000 ;
      RECT 0.000000 396.410000 2.500000 399.590000 ;
      RECT 1169.500000 395.590000 1186.000000 396.410000 ;
      RECT 1116.500000 395.590000 1156.500000 396.410000 ;
      RECT 1066.500000 395.590000 1108.500000 396.410000 ;
      RECT 1016.500000 395.590000 1058.500000 396.410000 ;
      RECT 966.500000 395.590000 1008.500000 396.410000 ;
      RECT 916.500000 395.590000 958.500000 396.410000 ;
      RECT 866.500000 395.590000 908.500000 396.410000 ;
      RECT 816.500000 395.590000 858.500000 396.410000 ;
      RECT 766.500000 395.590000 808.500000 396.410000 ;
      RECT 716.500000 395.590000 758.500000 396.410000 ;
      RECT 666.500000 395.590000 708.500000 396.410000 ;
      RECT 616.500000 395.590000 658.500000 396.410000 ;
      RECT 566.500000 395.590000 608.500000 396.410000 ;
      RECT 516.500000 395.590000 558.500000 396.410000 ;
      RECT 466.500000 395.590000 508.500000 396.410000 ;
      RECT 416.500000 395.590000 458.500000 396.410000 ;
      RECT 366.500000 395.590000 408.500000 396.410000 ;
      RECT 316.500000 395.590000 358.500000 396.410000 ;
      RECT 266.500000 395.590000 308.500000 396.410000 ;
      RECT 216.500000 395.590000 258.500000 396.410000 ;
      RECT 166.500000 395.590000 208.500000 396.410000 ;
      RECT 116.500000 395.590000 158.500000 396.410000 ;
      RECT 66.500000 395.590000 108.500000 396.410000 ;
      RECT 29.500000 395.590000 58.500000 396.410000 ;
      RECT 0.000000 395.590000 16.500000 396.410000 ;
      RECT 1169.500000 394.410000 1170.500000 395.590000 ;
      RECT 1116.500000 394.410000 1149.500000 395.590000 ;
      RECT 1107.500000 394.410000 1108.500000 395.590000 ;
      RECT 1066.500000 394.410000 1099.500000 395.590000 ;
      RECT 1057.500000 394.410000 1058.500000 395.590000 ;
      RECT 1016.500000 394.410000 1049.500000 395.590000 ;
      RECT 1007.500000 394.410000 1008.500000 395.590000 ;
      RECT 966.500000 394.410000 999.500000 395.590000 ;
      RECT 957.500000 394.410000 958.500000 395.590000 ;
      RECT 916.500000 394.410000 949.500000 395.590000 ;
      RECT 907.500000 394.410000 908.500000 395.590000 ;
      RECT 866.500000 394.410000 899.500000 395.590000 ;
      RECT 857.500000 394.410000 858.500000 395.590000 ;
      RECT 816.500000 394.410000 849.500000 395.590000 ;
      RECT 807.500000 394.410000 808.500000 395.590000 ;
      RECT 766.500000 394.410000 799.500000 395.590000 ;
      RECT 757.500000 394.410000 758.500000 395.590000 ;
      RECT 716.500000 394.410000 749.500000 395.590000 ;
      RECT 707.500000 394.410000 708.500000 395.590000 ;
      RECT 666.500000 394.410000 699.500000 395.590000 ;
      RECT 657.500000 394.410000 658.500000 395.590000 ;
      RECT 616.500000 394.410000 649.500000 395.590000 ;
      RECT 607.500000 394.410000 608.500000 395.590000 ;
      RECT 566.500000 394.410000 599.500000 395.590000 ;
      RECT 557.500000 394.410000 558.500000 395.590000 ;
      RECT 516.500000 394.410000 549.500000 395.590000 ;
      RECT 507.500000 394.410000 508.500000 395.590000 ;
      RECT 466.500000 394.410000 499.500000 395.590000 ;
      RECT 457.500000 394.410000 458.500000 395.590000 ;
      RECT 416.500000 394.410000 449.500000 395.590000 ;
      RECT 407.500000 394.410000 408.500000 395.590000 ;
      RECT 366.500000 394.410000 399.500000 395.590000 ;
      RECT 357.500000 394.410000 358.500000 395.590000 ;
      RECT 316.500000 394.410000 349.500000 395.590000 ;
      RECT 307.500000 394.410000 308.500000 395.590000 ;
      RECT 266.500000 394.410000 299.500000 395.590000 ;
      RECT 257.500000 394.410000 258.500000 395.590000 ;
      RECT 216.500000 394.410000 249.500000 395.590000 ;
      RECT 207.500000 394.410000 208.500000 395.590000 ;
      RECT 166.500000 394.410000 199.500000 395.590000 ;
      RECT 157.500000 394.410000 158.500000 395.590000 ;
      RECT 116.500000 394.410000 149.500000 395.590000 ;
      RECT 107.500000 394.410000 108.500000 395.590000 ;
      RECT 66.500000 394.410000 99.500000 395.590000 ;
      RECT 57.500000 394.410000 58.500000 395.590000 ;
      RECT 29.500000 394.410000 49.500000 395.590000 ;
      RECT 15.500000 394.410000 16.500000 395.590000 ;
      RECT 1157.500000 393.590000 1170.500000 394.410000 ;
      RECT 1107.500000 393.590000 1149.500000 394.410000 ;
      RECT 1057.500000 393.590000 1099.500000 394.410000 ;
      RECT 1007.500000 393.590000 1049.500000 394.410000 ;
      RECT 957.500000 393.590000 999.500000 394.410000 ;
      RECT 907.500000 393.590000 949.500000 394.410000 ;
      RECT 857.500000 393.590000 899.500000 394.410000 ;
      RECT 807.500000 393.590000 849.500000 394.410000 ;
      RECT 757.500000 393.590000 799.500000 394.410000 ;
      RECT 707.500000 393.590000 749.500000 394.410000 ;
      RECT 657.500000 393.590000 699.500000 394.410000 ;
      RECT 607.500000 393.590000 649.500000 394.410000 ;
      RECT 557.500000 393.590000 599.500000 394.410000 ;
      RECT 507.500000 393.590000 549.500000 394.410000 ;
      RECT 457.500000 393.590000 499.500000 394.410000 ;
      RECT 407.500000 393.590000 449.500000 394.410000 ;
      RECT 357.500000 393.590000 399.500000 394.410000 ;
      RECT 307.500000 393.590000 349.500000 394.410000 ;
      RECT 257.500000 393.590000 299.500000 394.410000 ;
      RECT 207.500000 393.590000 249.500000 394.410000 ;
      RECT 157.500000 393.590000 199.500000 394.410000 ;
      RECT 107.500000 393.590000 149.500000 394.410000 ;
      RECT 57.500000 393.590000 99.500000 394.410000 ;
      RECT 15.500000 393.590000 49.500000 394.410000 ;
      RECT 1183.500000 392.410000 1186.000000 395.590000 ;
      RECT 1169.500000 392.410000 1170.500000 393.590000 ;
      RECT 1116.500000 392.410000 1149.500000 393.590000 ;
      RECT 1107.500000 392.410000 1108.500000 393.590000 ;
      RECT 1066.500000 392.410000 1099.500000 393.590000 ;
      RECT 1057.500000 392.410000 1058.500000 393.590000 ;
      RECT 1016.500000 392.410000 1049.500000 393.590000 ;
      RECT 1007.500000 392.410000 1008.500000 393.590000 ;
      RECT 966.500000 392.410000 999.500000 393.590000 ;
      RECT 957.500000 392.410000 958.500000 393.590000 ;
      RECT 916.500000 392.410000 949.500000 393.590000 ;
      RECT 907.500000 392.410000 908.500000 393.590000 ;
      RECT 866.500000 392.410000 899.500000 393.590000 ;
      RECT 857.500000 392.410000 858.500000 393.590000 ;
      RECT 816.500000 392.410000 849.500000 393.590000 ;
      RECT 807.500000 392.410000 808.500000 393.590000 ;
      RECT 766.500000 392.410000 799.500000 393.590000 ;
      RECT 757.500000 392.410000 758.500000 393.590000 ;
      RECT 716.500000 392.410000 749.500000 393.590000 ;
      RECT 707.500000 392.410000 708.500000 393.590000 ;
      RECT 666.500000 392.410000 699.500000 393.590000 ;
      RECT 657.500000 392.410000 658.500000 393.590000 ;
      RECT 616.500000 392.410000 649.500000 393.590000 ;
      RECT 607.500000 392.410000 608.500000 393.590000 ;
      RECT 566.500000 392.410000 599.500000 393.590000 ;
      RECT 557.500000 392.410000 558.500000 393.590000 ;
      RECT 516.500000 392.410000 549.500000 393.590000 ;
      RECT 507.500000 392.410000 508.500000 393.590000 ;
      RECT 466.500000 392.410000 499.500000 393.590000 ;
      RECT 457.500000 392.410000 458.500000 393.590000 ;
      RECT 416.500000 392.410000 449.500000 393.590000 ;
      RECT 407.500000 392.410000 408.500000 393.590000 ;
      RECT 366.500000 392.410000 399.500000 393.590000 ;
      RECT 357.500000 392.410000 358.500000 393.590000 ;
      RECT 316.500000 392.410000 349.500000 393.590000 ;
      RECT 307.500000 392.410000 308.500000 393.590000 ;
      RECT 266.500000 392.410000 299.500000 393.590000 ;
      RECT 257.500000 392.410000 258.500000 393.590000 ;
      RECT 216.500000 392.410000 249.500000 393.590000 ;
      RECT 207.500000 392.410000 208.500000 393.590000 ;
      RECT 166.500000 392.410000 199.500000 393.590000 ;
      RECT 157.500000 392.410000 158.500000 393.590000 ;
      RECT 116.500000 392.410000 149.500000 393.590000 ;
      RECT 107.500000 392.410000 108.500000 393.590000 ;
      RECT 66.500000 392.410000 99.500000 393.590000 ;
      RECT 57.500000 392.410000 58.500000 393.590000 ;
      RECT 29.500000 392.410000 49.500000 393.590000 ;
      RECT 15.500000 392.410000 16.500000 393.590000 ;
      RECT 0.000000 392.410000 2.500000 395.590000 ;
      RECT 1169.500000 391.590000 1186.000000 392.410000 ;
      RECT 1116.500000 391.590000 1156.500000 392.410000 ;
      RECT 1066.500000 391.590000 1108.500000 392.410000 ;
      RECT 1016.500000 391.590000 1058.500000 392.410000 ;
      RECT 966.500000 391.590000 1008.500000 392.410000 ;
      RECT 916.500000 391.590000 958.500000 392.410000 ;
      RECT 866.500000 391.590000 908.500000 392.410000 ;
      RECT 816.500000 391.590000 858.500000 392.410000 ;
      RECT 766.500000 391.590000 808.500000 392.410000 ;
      RECT 716.500000 391.590000 758.500000 392.410000 ;
      RECT 666.500000 391.590000 708.500000 392.410000 ;
      RECT 616.500000 391.590000 658.500000 392.410000 ;
      RECT 566.500000 391.590000 608.500000 392.410000 ;
      RECT 516.500000 391.590000 558.500000 392.410000 ;
      RECT 466.500000 391.590000 508.500000 392.410000 ;
      RECT 416.500000 391.590000 458.500000 392.410000 ;
      RECT 366.500000 391.590000 408.500000 392.410000 ;
      RECT 316.500000 391.590000 358.500000 392.410000 ;
      RECT 266.500000 391.590000 308.500000 392.410000 ;
      RECT 216.500000 391.590000 258.500000 392.410000 ;
      RECT 166.500000 391.590000 208.500000 392.410000 ;
      RECT 116.500000 391.590000 158.500000 392.410000 ;
      RECT 66.500000 391.590000 108.500000 392.410000 ;
      RECT 29.500000 391.590000 58.500000 392.410000 ;
      RECT 0.000000 391.590000 16.500000 392.410000 ;
      RECT 1169.500000 390.410000 1170.500000 391.590000 ;
      RECT 1116.500000 390.410000 1149.500000 391.590000 ;
      RECT 1107.500000 390.410000 1108.500000 391.590000 ;
      RECT 1066.500000 390.410000 1099.500000 391.590000 ;
      RECT 1057.500000 390.410000 1058.500000 391.590000 ;
      RECT 1016.500000 390.410000 1049.500000 391.590000 ;
      RECT 1007.500000 390.410000 1008.500000 391.590000 ;
      RECT 966.500000 390.410000 999.500000 391.590000 ;
      RECT 957.500000 390.410000 958.500000 391.590000 ;
      RECT 916.500000 390.410000 949.500000 391.590000 ;
      RECT 907.500000 390.410000 908.500000 391.590000 ;
      RECT 866.500000 390.410000 899.500000 391.590000 ;
      RECT 857.500000 390.410000 858.500000 391.590000 ;
      RECT 816.500000 390.410000 849.500000 391.590000 ;
      RECT 807.500000 390.410000 808.500000 391.590000 ;
      RECT 766.500000 390.410000 799.500000 391.590000 ;
      RECT 757.500000 390.410000 758.500000 391.590000 ;
      RECT 716.500000 390.410000 749.500000 391.590000 ;
      RECT 707.500000 390.410000 708.500000 391.590000 ;
      RECT 666.500000 390.410000 699.500000 391.590000 ;
      RECT 657.500000 390.410000 658.500000 391.590000 ;
      RECT 616.500000 390.410000 649.500000 391.590000 ;
      RECT 607.500000 390.410000 608.500000 391.590000 ;
      RECT 566.500000 390.410000 599.500000 391.590000 ;
      RECT 557.500000 390.410000 558.500000 391.590000 ;
      RECT 516.500000 390.410000 549.500000 391.590000 ;
      RECT 507.500000 390.410000 508.500000 391.590000 ;
      RECT 466.500000 390.410000 499.500000 391.590000 ;
      RECT 457.500000 390.410000 458.500000 391.590000 ;
      RECT 416.500000 390.410000 449.500000 391.590000 ;
      RECT 407.500000 390.410000 408.500000 391.590000 ;
      RECT 366.500000 390.410000 399.500000 391.590000 ;
      RECT 357.500000 390.410000 358.500000 391.590000 ;
      RECT 316.500000 390.410000 349.500000 391.590000 ;
      RECT 307.500000 390.410000 308.500000 391.590000 ;
      RECT 266.500000 390.410000 299.500000 391.590000 ;
      RECT 257.500000 390.410000 258.500000 391.590000 ;
      RECT 216.500000 390.410000 249.500000 391.590000 ;
      RECT 207.500000 390.410000 208.500000 391.590000 ;
      RECT 166.500000 390.410000 199.500000 391.590000 ;
      RECT 157.500000 390.410000 158.500000 391.590000 ;
      RECT 116.500000 390.410000 149.500000 391.590000 ;
      RECT 107.500000 390.410000 108.500000 391.590000 ;
      RECT 66.500000 390.410000 99.500000 391.590000 ;
      RECT 57.500000 390.410000 58.500000 391.590000 ;
      RECT 29.500000 390.410000 49.500000 391.590000 ;
      RECT 15.500000 390.410000 16.500000 391.590000 ;
      RECT 1157.500000 389.590000 1170.500000 390.410000 ;
      RECT 1107.500000 389.590000 1149.500000 390.410000 ;
      RECT 1057.500000 389.590000 1099.500000 390.410000 ;
      RECT 1007.500000 389.590000 1049.500000 390.410000 ;
      RECT 957.500000 389.590000 999.500000 390.410000 ;
      RECT 907.500000 389.590000 949.500000 390.410000 ;
      RECT 857.500000 389.590000 899.500000 390.410000 ;
      RECT 807.500000 389.590000 849.500000 390.410000 ;
      RECT 757.500000 389.590000 799.500000 390.410000 ;
      RECT 707.500000 389.590000 749.500000 390.410000 ;
      RECT 657.500000 389.590000 699.500000 390.410000 ;
      RECT 607.500000 389.590000 649.500000 390.410000 ;
      RECT 557.500000 389.590000 599.500000 390.410000 ;
      RECT 507.500000 389.590000 549.500000 390.410000 ;
      RECT 457.500000 389.590000 499.500000 390.410000 ;
      RECT 407.500000 389.590000 449.500000 390.410000 ;
      RECT 357.500000 389.590000 399.500000 390.410000 ;
      RECT 307.500000 389.590000 349.500000 390.410000 ;
      RECT 257.500000 389.590000 299.500000 390.410000 ;
      RECT 207.500000 389.590000 249.500000 390.410000 ;
      RECT 157.500000 389.590000 199.500000 390.410000 ;
      RECT 107.500000 389.590000 149.500000 390.410000 ;
      RECT 57.500000 389.590000 99.500000 390.410000 ;
      RECT 15.500000 389.590000 49.500000 390.410000 ;
      RECT 1183.500000 388.410000 1186.000000 391.590000 ;
      RECT 1169.500000 388.410000 1170.500000 389.590000 ;
      RECT 1116.500000 388.410000 1149.500000 389.590000 ;
      RECT 1107.500000 388.410000 1108.500000 389.590000 ;
      RECT 1066.500000 388.410000 1099.500000 389.590000 ;
      RECT 1057.500000 388.410000 1058.500000 389.590000 ;
      RECT 1016.500000 388.410000 1049.500000 389.590000 ;
      RECT 1007.500000 388.410000 1008.500000 389.590000 ;
      RECT 966.500000 388.410000 999.500000 389.590000 ;
      RECT 957.500000 388.410000 958.500000 389.590000 ;
      RECT 916.500000 388.410000 949.500000 389.590000 ;
      RECT 907.500000 388.410000 908.500000 389.590000 ;
      RECT 866.500000 388.410000 899.500000 389.590000 ;
      RECT 857.500000 388.410000 858.500000 389.590000 ;
      RECT 816.500000 388.410000 849.500000 389.590000 ;
      RECT 807.500000 388.410000 808.500000 389.590000 ;
      RECT 766.500000 388.410000 799.500000 389.590000 ;
      RECT 757.500000 388.410000 758.500000 389.590000 ;
      RECT 716.500000 388.410000 749.500000 389.590000 ;
      RECT 707.500000 388.410000 708.500000 389.590000 ;
      RECT 666.500000 388.410000 699.500000 389.590000 ;
      RECT 657.500000 388.410000 658.500000 389.590000 ;
      RECT 616.500000 388.410000 649.500000 389.590000 ;
      RECT 607.500000 388.410000 608.500000 389.590000 ;
      RECT 566.500000 388.410000 599.500000 389.590000 ;
      RECT 557.500000 388.410000 558.500000 389.590000 ;
      RECT 516.500000 388.410000 549.500000 389.590000 ;
      RECT 507.500000 388.410000 508.500000 389.590000 ;
      RECT 466.500000 388.410000 499.500000 389.590000 ;
      RECT 457.500000 388.410000 458.500000 389.590000 ;
      RECT 416.500000 388.410000 449.500000 389.590000 ;
      RECT 407.500000 388.410000 408.500000 389.590000 ;
      RECT 366.500000 388.410000 399.500000 389.590000 ;
      RECT 357.500000 388.410000 358.500000 389.590000 ;
      RECT 316.500000 388.410000 349.500000 389.590000 ;
      RECT 307.500000 388.410000 308.500000 389.590000 ;
      RECT 266.500000 388.410000 299.500000 389.590000 ;
      RECT 257.500000 388.410000 258.500000 389.590000 ;
      RECT 216.500000 388.410000 249.500000 389.590000 ;
      RECT 207.500000 388.410000 208.500000 389.590000 ;
      RECT 166.500000 388.410000 199.500000 389.590000 ;
      RECT 157.500000 388.410000 158.500000 389.590000 ;
      RECT 116.500000 388.410000 149.500000 389.590000 ;
      RECT 107.500000 388.410000 108.500000 389.590000 ;
      RECT 66.500000 388.410000 99.500000 389.590000 ;
      RECT 57.500000 388.410000 58.500000 389.590000 ;
      RECT 29.500000 388.410000 49.500000 389.590000 ;
      RECT 15.500000 388.410000 16.500000 389.590000 ;
      RECT 0.000000 388.410000 2.500000 391.590000 ;
      RECT 1169.500000 387.590000 1186.000000 388.410000 ;
      RECT 1116.500000 387.590000 1156.500000 388.410000 ;
      RECT 1066.500000 387.590000 1108.500000 388.410000 ;
      RECT 1016.500000 387.590000 1058.500000 388.410000 ;
      RECT 966.500000 387.590000 1008.500000 388.410000 ;
      RECT 916.500000 387.590000 958.500000 388.410000 ;
      RECT 866.500000 387.590000 908.500000 388.410000 ;
      RECT 816.500000 387.590000 858.500000 388.410000 ;
      RECT 766.500000 387.590000 808.500000 388.410000 ;
      RECT 716.500000 387.590000 758.500000 388.410000 ;
      RECT 666.500000 387.590000 708.500000 388.410000 ;
      RECT 616.500000 387.590000 658.500000 388.410000 ;
      RECT 566.500000 387.590000 608.500000 388.410000 ;
      RECT 516.500000 387.590000 558.500000 388.410000 ;
      RECT 466.500000 387.590000 508.500000 388.410000 ;
      RECT 416.500000 387.590000 458.500000 388.410000 ;
      RECT 366.500000 387.590000 408.500000 388.410000 ;
      RECT 316.500000 387.590000 358.500000 388.410000 ;
      RECT 266.500000 387.590000 308.500000 388.410000 ;
      RECT 216.500000 387.590000 258.500000 388.410000 ;
      RECT 166.500000 387.590000 208.500000 388.410000 ;
      RECT 116.500000 387.590000 158.500000 388.410000 ;
      RECT 66.500000 387.590000 108.500000 388.410000 ;
      RECT 29.500000 387.590000 58.500000 388.410000 ;
      RECT 0.000000 387.590000 16.500000 388.410000 ;
      RECT 1169.500000 386.410000 1170.500000 387.590000 ;
      RECT 1116.500000 386.410000 1149.500000 387.590000 ;
      RECT 1107.500000 386.410000 1108.500000 387.590000 ;
      RECT 1066.500000 386.410000 1099.500000 387.590000 ;
      RECT 1057.500000 386.410000 1058.500000 387.590000 ;
      RECT 1016.500000 386.410000 1049.500000 387.590000 ;
      RECT 1007.500000 386.410000 1008.500000 387.590000 ;
      RECT 966.500000 386.410000 999.500000 387.590000 ;
      RECT 957.500000 386.410000 958.500000 387.590000 ;
      RECT 916.500000 386.410000 949.500000 387.590000 ;
      RECT 907.500000 386.410000 908.500000 387.590000 ;
      RECT 866.500000 386.410000 899.500000 387.590000 ;
      RECT 857.500000 386.410000 858.500000 387.590000 ;
      RECT 816.500000 386.410000 849.500000 387.590000 ;
      RECT 807.500000 386.410000 808.500000 387.590000 ;
      RECT 766.500000 386.410000 799.500000 387.590000 ;
      RECT 757.500000 386.410000 758.500000 387.590000 ;
      RECT 716.500000 386.410000 749.500000 387.590000 ;
      RECT 707.500000 386.410000 708.500000 387.590000 ;
      RECT 666.500000 386.410000 699.500000 387.590000 ;
      RECT 657.500000 386.410000 658.500000 387.590000 ;
      RECT 616.500000 386.410000 649.500000 387.590000 ;
      RECT 607.500000 386.410000 608.500000 387.590000 ;
      RECT 566.500000 386.410000 599.500000 387.590000 ;
      RECT 557.500000 386.410000 558.500000 387.590000 ;
      RECT 516.500000 386.410000 549.500000 387.590000 ;
      RECT 507.500000 386.410000 508.500000 387.590000 ;
      RECT 466.500000 386.410000 499.500000 387.590000 ;
      RECT 457.500000 386.410000 458.500000 387.590000 ;
      RECT 416.500000 386.410000 449.500000 387.590000 ;
      RECT 407.500000 386.410000 408.500000 387.590000 ;
      RECT 366.500000 386.410000 399.500000 387.590000 ;
      RECT 357.500000 386.410000 358.500000 387.590000 ;
      RECT 316.500000 386.410000 349.500000 387.590000 ;
      RECT 307.500000 386.410000 308.500000 387.590000 ;
      RECT 266.500000 386.410000 299.500000 387.590000 ;
      RECT 257.500000 386.410000 258.500000 387.590000 ;
      RECT 216.500000 386.410000 249.500000 387.590000 ;
      RECT 207.500000 386.410000 208.500000 387.590000 ;
      RECT 166.500000 386.410000 199.500000 387.590000 ;
      RECT 157.500000 386.410000 158.500000 387.590000 ;
      RECT 116.500000 386.410000 149.500000 387.590000 ;
      RECT 107.500000 386.410000 108.500000 387.590000 ;
      RECT 66.500000 386.410000 99.500000 387.590000 ;
      RECT 57.500000 386.410000 58.500000 387.590000 ;
      RECT 29.500000 386.410000 49.500000 387.590000 ;
      RECT 15.500000 386.410000 16.500000 387.590000 ;
      RECT 1157.500000 385.590000 1170.500000 386.410000 ;
      RECT 1107.500000 385.590000 1149.500000 386.410000 ;
      RECT 1057.500000 385.590000 1099.500000 386.410000 ;
      RECT 1007.500000 385.590000 1049.500000 386.410000 ;
      RECT 957.500000 385.590000 999.500000 386.410000 ;
      RECT 907.500000 385.590000 949.500000 386.410000 ;
      RECT 857.500000 385.590000 899.500000 386.410000 ;
      RECT 807.500000 385.590000 849.500000 386.410000 ;
      RECT 757.500000 385.590000 799.500000 386.410000 ;
      RECT 707.500000 385.590000 749.500000 386.410000 ;
      RECT 657.500000 385.590000 699.500000 386.410000 ;
      RECT 607.500000 385.590000 649.500000 386.410000 ;
      RECT 557.500000 385.590000 599.500000 386.410000 ;
      RECT 507.500000 385.590000 549.500000 386.410000 ;
      RECT 457.500000 385.590000 499.500000 386.410000 ;
      RECT 407.500000 385.590000 449.500000 386.410000 ;
      RECT 357.500000 385.590000 399.500000 386.410000 ;
      RECT 307.500000 385.590000 349.500000 386.410000 ;
      RECT 257.500000 385.590000 299.500000 386.410000 ;
      RECT 207.500000 385.590000 249.500000 386.410000 ;
      RECT 157.500000 385.590000 199.500000 386.410000 ;
      RECT 107.500000 385.590000 149.500000 386.410000 ;
      RECT 57.500000 385.590000 99.500000 386.410000 ;
      RECT 15.500000 385.590000 49.500000 386.410000 ;
      RECT 1183.500000 384.410000 1186.000000 387.590000 ;
      RECT 1169.500000 384.410000 1170.500000 385.590000 ;
      RECT 1116.500000 384.410000 1149.500000 385.590000 ;
      RECT 1107.500000 384.410000 1108.500000 385.590000 ;
      RECT 1066.500000 384.410000 1099.500000 385.590000 ;
      RECT 1057.500000 384.410000 1058.500000 385.590000 ;
      RECT 1016.500000 384.410000 1049.500000 385.590000 ;
      RECT 1007.500000 384.410000 1008.500000 385.590000 ;
      RECT 966.500000 384.410000 999.500000 385.590000 ;
      RECT 957.500000 384.410000 958.500000 385.590000 ;
      RECT 916.500000 384.410000 949.500000 385.590000 ;
      RECT 907.500000 384.410000 908.500000 385.590000 ;
      RECT 866.500000 384.410000 899.500000 385.590000 ;
      RECT 857.500000 384.410000 858.500000 385.590000 ;
      RECT 816.500000 384.410000 849.500000 385.590000 ;
      RECT 807.500000 384.410000 808.500000 385.590000 ;
      RECT 766.500000 384.410000 799.500000 385.590000 ;
      RECT 757.500000 384.410000 758.500000 385.590000 ;
      RECT 716.500000 384.410000 749.500000 385.590000 ;
      RECT 707.500000 384.410000 708.500000 385.590000 ;
      RECT 666.500000 384.410000 699.500000 385.590000 ;
      RECT 657.500000 384.410000 658.500000 385.590000 ;
      RECT 616.500000 384.410000 649.500000 385.590000 ;
      RECT 607.500000 384.410000 608.500000 385.590000 ;
      RECT 566.500000 384.410000 599.500000 385.590000 ;
      RECT 557.500000 384.410000 558.500000 385.590000 ;
      RECT 516.500000 384.410000 549.500000 385.590000 ;
      RECT 507.500000 384.410000 508.500000 385.590000 ;
      RECT 466.500000 384.410000 499.500000 385.590000 ;
      RECT 457.500000 384.410000 458.500000 385.590000 ;
      RECT 416.500000 384.410000 449.500000 385.590000 ;
      RECT 407.500000 384.410000 408.500000 385.590000 ;
      RECT 366.500000 384.410000 399.500000 385.590000 ;
      RECT 357.500000 384.410000 358.500000 385.590000 ;
      RECT 316.500000 384.410000 349.500000 385.590000 ;
      RECT 307.500000 384.410000 308.500000 385.590000 ;
      RECT 266.500000 384.410000 299.500000 385.590000 ;
      RECT 257.500000 384.410000 258.500000 385.590000 ;
      RECT 216.500000 384.410000 249.500000 385.590000 ;
      RECT 207.500000 384.410000 208.500000 385.590000 ;
      RECT 166.500000 384.410000 199.500000 385.590000 ;
      RECT 157.500000 384.410000 158.500000 385.590000 ;
      RECT 116.500000 384.410000 149.500000 385.590000 ;
      RECT 107.500000 384.410000 108.500000 385.590000 ;
      RECT 66.500000 384.410000 99.500000 385.590000 ;
      RECT 57.500000 384.410000 58.500000 385.590000 ;
      RECT 29.500000 384.410000 49.500000 385.590000 ;
      RECT 15.500000 384.410000 16.500000 385.590000 ;
      RECT 0.000000 384.410000 2.500000 387.590000 ;
      RECT 1169.500000 383.590000 1186.000000 384.410000 ;
      RECT 1116.500000 383.590000 1156.500000 384.410000 ;
      RECT 1066.500000 383.590000 1108.500000 384.410000 ;
      RECT 1016.500000 383.590000 1058.500000 384.410000 ;
      RECT 966.500000 383.590000 1008.500000 384.410000 ;
      RECT 916.500000 383.590000 958.500000 384.410000 ;
      RECT 866.500000 383.590000 908.500000 384.410000 ;
      RECT 816.500000 383.590000 858.500000 384.410000 ;
      RECT 766.500000 383.590000 808.500000 384.410000 ;
      RECT 716.500000 383.590000 758.500000 384.410000 ;
      RECT 666.500000 383.590000 708.500000 384.410000 ;
      RECT 616.500000 383.590000 658.500000 384.410000 ;
      RECT 566.500000 383.590000 608.500000 384.410000 ;
      RECT 516.500000 383.590000 558.500000 384.410000 ;
      RECT 466.500000 383.590000 508.500000 384.410000 ;
      RECT 416.500000 383.590000 458.500000 384.410000 ;
      RECT 366.500000 383.590000 408.500000 384.410000 ;
      RECT 316.500000 383.590000 358.500000 384.410000 ;
      RECT 266.500000 383.590000 308.500000 384.410000 ;
      RECT 216.500000 383.590000 258.500000 384.410000 ;
      RECT 166.500000 383.590000 208.500000 384.410000 ;
      RECT 116.500000 383.590000 158.500000 384.410000 ;
      RECT 66.500000 383.590000 108.500000 384.410000 ;
      RECT 29.500000 383.590000 58.500000 384.410000 ;
      RECT 0.000000 383.590000 16.500000 384.410000 ;
      RECT 1169.500000 382.410000 1170.500000 383.590000 ;
      RECT 1116.500000 382.410000 1149.500000 383.590000 ;
      RECT 1107.500000 382.410000 1108.500000 383.590000 ;
      RECT 1066.500000 382.410000 1099.500000 383.590000 ;
      RECT 1057.500000 382.410000 1058.500000 383.590000 ;
      RECT 1016.500000 382.410000 1049.500000 383.590000 ;
      RECT 1007.500000 382.410000 1008.500000 383.590000 ;
      RECT 966.500000 382.410000 999.500000 383.590000 ;
      RECT 957.500000 382.410000 958.500000 383.590000 ;
      RECT 916.500000 382.410000 949.500000 383.590000 ;
      RECT 907.500000 382.410000 908.500000 383.590000 ;
      RECT 866.500000 382.410000 899.500000 383.590000 ;
      RECT 857.500000 382.410000 858.500000 383.590000 ;
      RECT 816.500000 382.410000 849.500000 383.590000 ;
      RECT 807.500000 382.410000 808.500000 383.590000 ;
      RECT 766.500000 382.410000 799.500000 383.590000 ;
      RECT 757.500000 382.410000 758.500000 383.590000 ;
      RECT 716.500000 382.410000 749.500000 383.590000 ;
      RECT 707.500000 382.410000 708.500000 383.590000 ;
      RECT 666.500000 382.410000 699.500000 383.590000 ;
      RECT 657.500000 382.410000 658.500000 383.590000 ;
      RECT 616.500000 382.410000 649.500000 383.590000 ;
      RECT 607.500000 382.410000 608.500000 383.590000 ;
      RECT 566.500000 382.410000 599.500000 383.590000 ;
      RECT 557.500000 382.410000 558.500000 383.590000 ;
      RECT 516.500000 382.410000 549.500000 383.590000 ;
      RECT 507.500000 382.410000 508.500000 383.590000 ;
      RECT 466.500000 382.410000 499.500000 383.590000 ;
      RECT 457.500000 382.410000 458.500000 383.590000 ;
      RECT 416.500000 382.410000 449.500000 383.590000 ;
      RECT 407.500000 382.410000 408.500000 383.590000 ;
      RECT 366.500000 382.410000 399.500000 383.590000 ;
      RECT 357.500000 382.410000 358.500000 383.590000 ;
      RECT 316.500000 382.410000 349.500000 383.590000 ;
      RECT 307.500000 382.410000 308.500000 383.590000 ;
      RECT 266.500000 382.410000 299.500000 383.590000 ;
      RECT 257.500000 382.410000 258.500000 383.590000 ;
      RECT 216.500000 382.410000 249.500000 383.590000 ;
      RECT 207.500000 382.410000 208.500000 383.590000 ;
      RECT 166.500000 382.410000 199.500000 383.590000 ;
      RECT 157.500000 382.410000 158.500000 383.590000 ;
      RECT 116.500000 382.410000 149.500000 383.590000 ;
      RECT 107.500000 382.410000 108.500000 383.590000 ;
      RECT 66.500000 382.410000 99.500000 383.590000 ;
      RECT 57.500000 382.410000 58.500000 383.590000 ;
      RECT 29.500000 382.410000 49.500000 383.590000 ;
      RECT 15.500000 382.410000 16.500000 383.590000 ;
      RECT 1157.500000 381.590000 1170.500000 382.410000 ;
      RECT 1107.500000 381.590000 1149.500000 382.410000 ;
      RECT 1057.500000 381.590000 1099.500000 382.410000 ;
      RECT 1007.500000 381.590000 1049.500000 382.410000 ;
      RECT 957.500000 381.590000 999.500000 382.410000 ;
      RECT 907.500000 381.590000 949.500000 382.410000 ;
      RECT 857.500000 381.590000 899.500000 382.410000 ;
      RECT 807.500000 381.590000 849.500000 382.410000 ;
      RECT 757.500000 381.590000 799.500000 382.410000 ;
      RECT 707.500000 381.590000 749.500000 382.410000 ;
      RECT 657.500000 381.590000 699.500000 382.410000 ;
      RECT 607.500000 381.590000 649.500000 382.410000 ;
      RECT 557.500000 381.590000 599.500000 382.410000 ;
      RECT 507.500000 381.590000 549.500000 382.410000 ;
      RECT 457.500000 381.590000 499.500000 382.410000 ;
      RECT 407.500000 381.590000 449.500000 382.410000 ;
      RECT 357.500000 381.590000 399.500000 382.410000 ;
      RECT 307.500000 381.590000 349.500000 382.410000 ;
      RECT 257.500000 381.590000 299.500000 382.410000 ;
      RECT 207.500000 381.590000 249.500000 382.410000 ;
      RECT 157.500000 381.590000 199.500000 382.410000 ;
      RECT 107.500000 381.590000 149.500000 382.410000 ;
      RECT 57.500000 381.590000 99.500000 382.410000 ;
      RECT 15.500000 381.590000 49.500000 382.410000 ;
      RECT 1183.500000 380.410000 1186.000000 383.590000 ;
      RECT 1169.500000 380.410000 1170.500000 381.590000 ;
      RECT 1116.500000 380.410000 1149.500000 381.590000 ;
      RECT 1107.500000 380.410000 1108.500000 381.590000 ;
      RECT 1066.500000 380.410000 1099.500000 381.590000 ;
      RECT 1057.500000 380.410000 1058.500000 381.590000 ;
      RECT 1016.500000 380.410000 1049.500000 381.590000 ;
      RECT 1007.500000 380.410000 1008.500000 381.590000 ;
      RECT 966.500000 380.410000 999.500000 381.590000 ;
      RECT 957.500000 380.410000 958.500000 381.590000 ;
      RECT 916.500000 380.410000 949.500000 381.590000 ;
      RECT 907.500000 380.410000 908.500000 381.590000 ;
      RECT 866.500000 380.410000 899.500000 381.590000 ;
      RECT 857.500000 380.410000 858.500000 381.590000 ;
      RECT 816.500000 380.410000 849.500000 381.590000 ;
      RECT 807.500000 380.410000 808.500000 381.590000 ;
      RECT 766.500000 380.410000 799.500000 381.590000 ;
      RECT 757.500000 380.410000 758.500000 381.590000 ;
      RECT 716.500000 380.410000 749.500000 381.590000 ;
      RECT 707.500000 380.410000 708.500000 381.590000 ;
      RECT 666.500000 380.410000 699.500000 381.590000 ;
      RECT 657.500000 380.410000 658.500000 381.590000 ;
      RECT 616.500000 380.410000 649.500000 381.590000 ;
      RECT 607.500000 380.410000 608.500000 381.590000 ;
      RECT 566.500000 380.410000 599.500000 381.590000 ;
      RECT 557.500000 380.410000 558.500000 381.590000 ;
      RECT 516.500000 380.410000 549.500000 381.590000 ;
      RECT 507.500000 380.410000 508.500000 381.590000 ;
      RECT 466.500000 380.410000 499.500000 381.590000 ;
      RECT 457.500000 380.410000 458.500000 381.590000 ;
      RECT 416.500000 380.410000 449.500000 381.590000 ;
      RECT 407.500000 380.410000 408.500000 381.590000 ;
      RECT 366.500000 380.410000 399.500000 381.590000 ;
      RECT 357.500000 380.410000 358.500000 381.590000 ;
      RECT 316.500000 380.410000 349.500000 381.590000 ;
      RECT 307.500000 380.410000 308.500000 381.590000 ;
      RECT 266.500000 380.410000 299.500000 381.590000 ;
      RECT 257.500000 380.410000 258.500000 381.590000 ;
      RECT 216.500000 380.410000 249.500000 381.590000 ;
      RECT 207.500000 380.410000 208.500000 381.590000 ;
      RECT 166.500000 380.410000 199.500000 381.590000 ;
      RECT 157.500000 380.410000 158.500000 381.590000 ;
      RECT 116.500000 380.410000 149.500000 381.590000 ;
      RECT 107.500000 380.410000 108.500000 381.590000 ;
      RECT 66.500000 380.410000 99.500000 381.590000 ;
      RECT 57.500000 380.410000 58.500000 381.590000 ;
      RECT 29.500000 380.410000 49.500000 381.590000 ;
      RECT 15.500000 380.410000 16.500000 381.590000 ;
      RECT 0.000000 380.410000 2.500000 383.590000 ;
      RECT 1169.500000 379.590000 1186.000000 380.410000 ;
      RECT 1116.500000 379.590000 1156.500000 380.410000 ;
      RECT 1066.500000 379.590000 1108.500000 380.410000 ;
      RECT 1016.500000 379.590000 1058.500000 380.410000 ;
      RECT 966.500000 379.590000 1008.500000 380.410000 ;
      RECT 916.500000 379.590000 958.500000 380.410000 ;
      RECT 866.500000 379.590000 908.500000 380.410000 ;
      RECT 816.500000 379.590000 858.500000 380.410000 ;
      RECT 766.500000 379.590000 808.500000 380.410000 ;
      RECT 716.500000 379.590000 758.500000 380.410000 ;
      RECT 666.500000 379.590000 708.500000 380.410000 ;
      RECT 616.500000 379.590000 658.500000 380.410000 ;
      RECT 566.500000 379.590000 608.500000 380.410000 ;
      RECT 516.500000 379.590000 558.500000 380.410000 ;
      RECT 466.500000 379.590000 508.500000 380.410000 ;
      RECT 416.500000 379.590000 458.500000 380.410000 ;
      RECT 366.500000 379.590000 408.500000 380.410000 ;
      RECT 316.500000 379.590000 358.500000 380.410000 ;
      RECT 266.500000 379.590000 308.500000 380.410000 ;
      RECT 216.500000 379.590000 258.500000 380.410000 ;
      RECT 166.500000 379.590000 208.500000 380.410000 ;
      RECT 116.500000 379.590000 158.500000 380.410000 ;
      RECT 66.500000 379.590000 108.500000 380.410000 ;
      RECT 29.500000 379.590000 58.500000 380.410000 ;
      RECT 0.000000 379.590000 16.500000 380.410000 ;
      RECT 1169.500000 378.410000 1170.500000 379.590000 ;
      RECT 1116.500000 378.410000 1149.500000 379.590000 ;
      RECT 1107.500000 378.410000 1108.500000 379.590000 ;
      RECT 1066.500000 378.410000 1099.500000 379.590000 ;
      RECT 1057.500000 378.410000 1058.500000 379.590000 ;
      RECT 1016.500000 378.410000 1049.500000 379.590000 ;
      RECT 1007.500000 378.410000 1008.500000 379.590000 ;
      RECT 966.500000 378.410000 999.500000 379.590000 ;
      RECT 957.500000 378.410000 958.500000 379.590000 ;
      RECT 916.500000 378.410000 949.500000 379.590000 ;
      RECT 907.500000 378.410000 908.500000 379.590000 ;
      RECT 866.500000 378.410000 899.500000 379.590000 ;
      RECT 857.500000 378.410000 858.500000 379.590000 ;
      RECT 816.500000 378.410000 849.500000 379.590000 ;
      RECT 807.500000 378.410000 808.500000 379.590000 ;
      RECT 766.500000 378.410000 799.500000 379.590000 ;
      RECT 757.500000 378.410000 758.500000 379.590000 ;
      RECT 716.500000 378.410000 749.500000 379.590000 ;
      RECT 707.500000 378.410000 708.500000 379.590000 ;
      RECT 666.500000 378.410000 699.500000 379.590000 ;
      RECT 657.500000 378.410000 658.500000 379.590000 ;
      RECT 616.500000 378.410000 649.500000 379.590000 ;
      RECT 607.500000 378.410000 608.500000 379.590000 ;
      RECT 566.500000 378.410000 599.500000 379.590000 ;
      RECT 557.500000 378.410000 558.500000 379.590000 ;
      RECT 516.500000 378.410000 549.500000 379.590000 ;
      RECT 507.500000 378.410000 508.500000 379.590000 ;
      RECT 466.500000 378.410000 499.500000 379.590000 ;
      RECT 457.500000 378.410000 458.500000 379.590000 ;
      RECT 416.500000 378.410000 449.500000 379.590000 ;
      RECT 407.500000 378.410000 408.500000 379.590000 ;
      RECT 366.500000 378.410000 399.500000 379.590000 ;
      RECT 357.500000 378.410000 358.500000 379.590000 ;
      RECT 316.500000 378.410000 349.500000 379.590000 ;
      RECT 307.500000 378.410000 308.500000 379.590000 ;
      RECT 266.500000 378.410000 299.500000 379.590000 ;
      RECT 257.500000 378.410000 258.500000 379.590000 ;
      RECT 216.500000 378.410000 249.500000 379.590000 ;
      RECT 207.500000 378.410000 208.500000 379.590000 ;
      RECT 166.500000 378.410000 199.500000 379.590000 ;
      RECT 157.500000 378.410000 158.500000 379.590000 ;
      RECT 116.500000 378.410000 149.500000 379.590000 ;
      RECT 107.500000 378.410000 108.500000 379.590000 ;
      RECT 66.500000 378.410000 99.500000 379.590000 ;
      RECT 57.500000 378.410000 58.500000 379.590000 ;
      RECT 29.500000 378.410000 49.500000 379.590000 ;
      RECT 15.500000 378.410000 16.500000 379.590000 ;
      RECT 1157.500000 377.590000 1170.500000 378.410000 ;
      RECT 1107.500000 377.590000 1149.500000 378.410000 ;
      RECT 1057.500000 377.590000 1099.500000 378.410000 ;
      RECT 1007.500000 377.590000 1049.500000 378.410000 ;
      RECT 957.500000 377.590000 999.500000 378.410000 ;
      RECT 907.500000 377.590000 949.500000 378.410000 ;
      RECT 857.500000 377.590000 899.500000 378.410000 ;
      RECT 807.500000 377.590000 849.500000 378.410000 ;
      RECT 757.500000 377.590000 799.500000 378.410000 ;
      RECT 707.500000 377.590000 749.500000 378.410000 ;
      RECT 657.500000 377.590000 699.500000 378.410000 ;
      RECT 607.500000 377.590000 649.500000 378.410000 ;
      RECT 557.500000 377.590000 599.500000 378.410000 ;
      RECT 507.500000 377.590000 549.500000 378.410000 ;
      RECT 457.500000 377.590000 499.500000 378.410000 ;
      RECT 407.500000 377.590000 449.500000 378.410000 ;
      RECT 357.500000 377.590000 399.500000 378.410000 ;
      RECT 307.500000 377.590000 349.500000 378.410000 ;
      RECT 257.500000 377.590000 299.500000 378.410000 ;
      RECT 207.500000 377.590000 249.500000 378.410000 ;
      RECT 157.500000 377.590000 199.500000 378.410000 ;
      RECT 107.500000 377.590000 149.500000 378.410000 ;
      RECT 57.500000 377.590000 99.500000 378.410000 ;
      RECT 15.500000 377.590000 49.500000 378.410000 ;
      RECT 1183.500000 376.410000 1186.000000 379.590000 ;
      RECT 1169.500000 376.410000 1170.500000 377.590000 ;
      RECT 1116.500000 376.410000 1149.500000 377.590000 ;
      RECT 1107.500000 376.410000 1108.500000 377.590000 ;
      RECT 1066.500000 376.410000 1099.500000 377.590000 ;
      RECT 1057.500000 376.410000 1058.500000 377.590000 ;
      RECT 1016.500000 376.410000 1049.500000 377.590000 ;
      RECT 1007.500000 376.410000 1008.500000 377.590000 ;
      RECT 966.500000 376.410000 999.500000 377.590000 ;
      RECT 957.500000 376.410000 958.500000 377.590000 ;
      RECT 916.500000 376.410000 949.500000 377.590000 ;
      RECT 907.500000 376.410000 908.500000 377.590000 ;
      RECT 866.500000 376.410000 899.500000 377.590000 ;
      RECT 857.500000 376.410000 858.500000 377.590000 ;
      RECT 816.500000 376.410000 849.500000 377.590000 ;
      RECT 807.500000 376.410000 808.500000 377.590000 ;
      RECT 766.500000 376.410000 799.500000 377.590000 ;
      RECT 757.500000 376.410000 758.500000 377.590000 ;
      RECT 716.500000 376.410000 749.500000 377.590000 ;
      RECT 707.500000 376.410000 708.500000 377.590000 ;
      RECT 666.500000 376.410000 699.500000 377.590000 ;
      RECT 657.500000 376.410000 658.500000 377.590000 ;
      RECT 616.500000 376.410000 649.500000 377.590000 ;
      RECT 607.500000 376.410000 608.500000 377.590000 ;
      RECT 566.500000 376.410000 599.500000 377.590000 ;
      RECT 557.500000 376.410000 558.500000 377.590000 ;
      RECT 516.500000 376.410000 549.500000 377.590000 ;
      RECT 507.500000 376.410000 508.500000 377.590000 ;
      RECT 466.500000 376.410000 499.500000 377.590000 ;
      RECT 457.500000 376.410000 458.500000 377.590000 ;
      RECT 416.500000 376.410000 449.500000 377.590000 ;
      RECT 407.500000 376.410000 408.500000 377.590000 ;
      RECT 366.500000 376.410000 399.500000 377.590000 ;
      RECT 357.500000 376.410000 358.500000 377.590000 ;
      RECT 316.500000 376.410000 349.500000 377.590000 ;
      RECT 307.500000 376.410000 308.500000 377.590000 ;
      RECT 266.500000 376.410000 299.500000 377.590000 ;
      RECT 257.500000 376.410000 258.500000 377.590000 ;
      RECT 216.500000 376.410000 249.500000 377.590000 ;
      RECT 207.500000 376.410000 208.500000 377.590000 ;
      RECT 166.500000 376.410000 199.500000 377.590000 ;
      RECT 157.500000 376.410000 158.500000 377.590000 ;
      RECT 116.500000 376.410000 149.500000 377.590000 ;
      RECT 107.500000 376.410000 108.500000 377.590000 ;
      RECT 66.500000 376.410000 99.500000 377.590000 ;
      RECT 57.500000 376.410000 58.500000 377.590000 ;
      RECT 29.500000 376.410000 49.500000 377.590000 ;
      RECT 15.500000 376.410000 16.500000 377.590000 ;
      RECT 0.000000 376.410000 2.500000 379.590000 ;
      RECT 1169.500000 375.590000 1186.000000 376.410000 ;
      RECT 1116.500000 375.590000 1156.500000 376.410000 ;
      RECT 1066.500000 375.590000 1108.500000 376.410000 ;
      RECT 1016.500000 375.590000 1058.500000 376.410000 ;
      RECT 966.500000 375.590000 1008.500000 376.410000 ;
      RECT 916.500000 375.590000 958.500000 376.410000 ;
      RECT 866.500000 375.590000 908.500000 376.410000 ;
      RECT 816.500000 375.590000 858.500000 376.410000 ;
      RECT 766.500000 375.590000 808.500000 376.410000 ;
      RECT 716.500000 375.590000 758.500000 376.410000 ;
      RECT 666.500000 375.590000 708.500000 376.410000 ;
      RECT 616.500000 375.590000 658.500000 376.410000 ;
      RECT 566.500000 375.590000 608.500000 376.410000 ;
      RECT 516.500000 375.590000 558.500000 376.410000 ;
      RECT 466.500000 375.590000 508.500000 376.410000 ;
      RECT 416.500000 375.590000 458.500000 376.410000 ;
      RECT 366.500000 375.590000 408.500000 376.410000 ;
      RECT 316.500000 375.590000 358.500000 376.410000 ;
      RECT 266.500000 375.590000 308.500000 376.410000 ;
      RECT 216.500000 375.590000 258.500000 376.410000 ;
      RECT 166.500000 375.590000 208.500000 376.410000 ;
      RECT 116.500000 375.590000 158.500000 376.410000 ;
      RECT 66.500000 375.590000 108.500000 376.410000 ;
      RECT 29.500000 375.590000 58.500000 376.410000 ;
      RECT 0.000000 375.590000 16.500000 376.410000 ;
      RECT 1169.500000 374.410000 1170.500000 375.590000 ;
      RECT 1116.500000 374.410000 1149.500000 375.590000 ;
      RECT 1107.500000 374.410000 1108.500000 375.590000 ;
      RECT 1066.500000 374.410000 1099.500000 375.590000 ;
      RECT 1057.500000 374.410000 1058.500000 375.590000 ;
      RECT 1016.500000 374.410000 1049.500000 375.590000 ;
      RECT 1007.500000 374.410000 1008.500000 375.590000 ;
      RECT 966.500000 374.410000 999.500000 375.590000 ;
      RECT 957.500000 374.410000 958.500000 375.590000 ;
      RECT 916.500000 374.410000 949.500000 375.590000 ;
      RECT 907.500000 374.410000 908.500000 375.590000 ;
      RECT 866.500000 374.410000 899.500000 375.590000 ;
      RECT 857.500000 374.410000 858.500000 375.590000 ;
      RECT 816.500000 374.410000 849.500000 375.590000 ;
      RECT 807.500000 374.410000 808.500000 375.590000 ;
      RECT 766.500000 374.410000 799.500000 375.590000 ;
      RECT 757.500000 374.410000 758.500000 375.590000 ;
      RECT 716.500000 374.410000 749.500000 375.590000 ;
      RECT 707.500000 374.410000 708.500000 375.590000 ;
      RECT 666.500000 374.410000 699.500000 375.590000 ;
      RECT 657.500000 374.410000 658.500000 375.590000 ;
      RECT 616.500000 374.410000 649.500000 375.590000 ;
      RECT 607.500000 374.410000 608.500000 375.590000 ;
      RECT 566.500000 374.410000 599.500000 375.590000 ;
      RECT 557.500000 374.410000 558.500000 375.590000 ;
      RECT 516.500000 374.410000 549.500000 375.590000 ;
      RECT 507.500000 374.410000 508.500000 375.590000 ;
      RECT 466.500000 374.410000 499.500000 375.590000 ;
      RECT 457.500000 374.410000 458.500000 375.590000 ;
      RECT 416.500000 374.410000 449.500000 375.590000 ;
      RECT 407.500000 374.410000 408.500000 375.590000 ;
      RECT 366.500000 374.410000 399.500000 375.590000 ;
      RECT 357.500000 374.410000 358.500000 375.590000 ;
      RECT 316.500000 374.410000 349.500000 375.590000 ;
      RECT 307.500000 374.410000 308.500000 375.590000 ;
      RECT 266.500000 374.410000 299.500000 375.590000 ;
      RECT 257.500000 374.410000 258.500000 375.590000 ;
      RECT 216.500000 374.410000 249.500000 375.590000 ;
      RECT 207.500000 374.410000 208.500000 375.590000 ;
      RECT 166.500000 374.410000 199.500000 375.590000 ;
      RECT 157.500000 374.410000 158.500000 375.590000 ;
      RECT 116.500000 374.410000 149.500000 375.590000 ;
      RECT 107.500000 374.410000 108.500000 375.590000 ;
      RECT 66.500000 374.410000 99.500000 375.590000 ;
      RECT 57.500000 374.410000 58.500000 375.590000 ;
      RECT 29.500000 374.410000 49.500000 375.590000 ;
      RECT 15.500000 374.410000 16.500000 375.590000 ;
      RECT 1157.500000 373.590000 1170.500000 374.410000 ;
      RECT 1107.500000 373.590000 1149.500000 374.410000 ;
      RECT 1057.500000 373.590000 1099.500000 374.410000 ;
      RECT 1007.500000 373.590000 1049.500000 374.410000 ;
      RECT 957.500000 373.590000 999.500000 374.410000 ;
      RECT 907.500000 373.590000 949.500000 374.410000 ;
      RECT 857.500000 373.590000 899.500000 374.410000 ;
      RECT 807.500000 373.590000 849.500000 374.410000 ;
      RECT 757.500000 373.590000 799.500000 374.410000 ;
      RECT 707.500000 373.590000 749.500000 374.410000 ;
      RECT 657.500000 373.590000 699.500000 374.410000 ;
      RECT 607.500000 373.590000 649.500000 374.410000 ;
      RECT 557.500000 373.590000 599.500000 374.410000 ;
      RECT 507.500000 373.590000 549.500000 374.410000 ;
      RECT 457.500000 373.590000 499.500000 374.410000 ;
      RECT 407.500000 373.590000 449.500000 374.410000 ;
      RECT 357.500000 373.590000 399.500000 374.410000 ;
      RECT 307.500000 373.590000 349.500000 374.410000 ;
      RECT 257.500000 373.590000 299.500000 374.410000 ;
      RECT 207.500000 373.590000 249.500000 374.410000 ;
      RECT 157.500000 373.590000 199.500000 374.410000 ;
      RECT 107.500000 373.590000 149.500000 374.410000 ;
      RECT 57.500000 373.590000 99.500000 374.410000 ;
      RECT 15.500000 373.590000 49.500000 374.410000 ;
      RECT 1183.500000 372.410000 1186.000000 375.590000 ;
      RECT 1169.500000 372.410000 1170.500000 373.590000 ;
      RECT 1116.500000 372.410000 1149.500000 373.590000 ;
      RECT 1107.500000 372.410000 1108.500000 373.590000 ;
      RECT 1066.500000 372.410000 1099.500000 373.590000 ;
      RECT 1057.500000 372.410000 1058.500000 373.590000 ;
      RECT 1016.500000 372.410000 1049.500000 373.590000 ;
      RECT 1007.500000 372.410000 1008.500000 373.590000 ;
      RECT 966.500000 372.410000 999.500000 373.590000 ;
      RECT 957.500000 372.410000 958.500000 373.590000 ;
      RECT 916.500000 372.410000 949.500000 373.590000 ;
      RECT 907.500000 372.410000 908.500000 373.590000 ;
      RECT 866.500000 372.410000 899.500000 373.590000 ;
      RECT 857.500000 372.410000 858.500000 373.590000 ;
      RECT 816.500000 372.410000 849.500000 373.590000 ;
      RECT 807.500000 372.410000 808.500000 373.590000 ;
      RECT 766.500000 372.410000 799.500000 373.590000 ;
      RECT 757.500000 372.410000 758.500000 373.590000 ;
      RECT 716.500000 372.410000 749.500000 373.590000 ;
      RECT 707.500000 372.410000 708.500000 373.590000 ;
      RECT 666.500000 372.410000 699.500000 373.590000 ;
      RECT 657.500000 372.410000 658.500000 373.590000 ;
      RECT 616.500000 372.410000 649.500000 373.590000 ;
      RECT 607.500000 372.410000 608.500000 373.590000 ;
      RECT 566.500000 372.410000 599.500000 373.590000 ;
      RECT 557.500000 372.410000 558.500000 373.590000 ;
      RECT 516.500000 372.410000 549.500000 373.590000 ;
      RECT 507.500000 372.410000 508.500000 373.590000 ;
      RECT 466.500000 372.410000 499.500000 373.590000 ;
      RECT 457.500000 372.410000 458.500000 373.590000 ;
      RECT 416.500000 372.410000 449.500000 373.590000 ;
      RECT 407.500000 372.410000 408.500000 373.590000 ;
      RECT 366.500000 372.410000 399.500000 373.590000 ;
      RECT 357.500000 372.410000 358.500000 373.590000 ;
      RECT 316.500000 372.410000 349.500000 373.590000 ;
      RECT 307.500000 372.410000 308.500000 373.590000 ;
      RECT 266.500000 372.410000 299.500000 373.590000 ;
      RECT 257.500000 372.410000 258.500000 373.590000 ;
      RECT 216.500000 372.410000 249.500000 373.590000 ;
      RECT 207.500000 372.410000 208.500000 373.590000 ;
      RECT 166.500000 372.410000 199.500000 373.590000 ;
      RECT 157.500000 372.410000 158.500000 373.590000 ;
      RECT 116.500000 372.410000 149.500000 373.590000 ;
      RECT 107.500000 372.410000 108.500000 373.590000 ;
      RECT 66.500000 372.410000 99.500000 373.590000 ;
      RECT 57.500000 372.410000 58.500000 373.590000 ;
      RECT 29.500000 372.410000 49.500000 373.590000 ;
      RECT 15.500000 372.410000 16.500000 373.590000 ;
      RECT 0.000000 372.410000 2.500000 375.590000 ;
      RECT 1169.500000 371.590000 1186.000000 372.410000 ;
      RECT 1116.500000 371.590000 1156.500000 372.410000 ;
      RECT 1066.500000 371.590000 1108.500000 372.410000 ;
      RECT 1016.500000 371.590000 1058.500000 372.410000 ;
      RECT 966.500000 371.590000 1008.500000 372.410000 ;
      RECT 916.500000 371.590000 958.500000 372.410000 ;
      RECT 866.500000 371.590000 908.500000 372.410000 ;
      RECT 816.500000 371.590000 858.500000 372.410000 ;
      RECT 766.500000 371.590000 808.500000 372.410000 ;
      RECT 716.500000 371.590000 758.500000 372.410000 ;
      RECT 666.500000 371.590000 708.500000 372.410000 ;
      RECT 616.500000 371.590000 658.500000 372.410000 ;
      RECT 566.500000 371.590000 608.500000 372.410000 ;
      RECT 516.500000 371.590000 558.500000 372.410000 ;
      RECT 466.500000 371.590000 508.500000 372.410000 ;
      RECT 416.500000 371.590000 458.500000 372.410000 ;
      RECT 366.500000 371.590000 408.500000 372.410000 ;
      RECT 316.500000 371.590000 358.500000 372.410000 ;
      RECT 266.500000 371.590000 308.500000 372.410000 ;
      RECT 216.500000 371.590000 258.500000 372.410000 ;
      RECT 166.500000 371.590000 208.500000 372.410000 ;
      RECT 116.500000 371.590000 158.500000 372.410000 ;
      RECT 66.500000 371.590000 108.500000 372.410000 ;
      RECT 29.500000 371.590000 58.500000 372.410000 ;
      RECT 0.000000 371.590000 16.500000 372.410000 ;
      RECT 1169.500000 370.410000 1170.500000 371.590000 ;
      RECT 1116.500000 370.410000 1149.500000 371.590000 ;
      RECT 1107.500000 370.410000 1108.500000 371.590000 ;
      RECT 1066.500000 370.410000 1099.500000 371.590000 ;
      RECT 1057.500000 370.410000 1058.500000 371.590000 ;
      RECT 1016.500000 370.410000 1049.500000 371.590000 ;
      RECT 1007.500000 370.410000 1008.500000 371.590000 ;
      RECT 966.500000 370.410000 999.500000 371.590000 ;
      RECT 957.500000 370.410000 958.500000 371.590000 ;
      RECT 916.500000 370.410000 949.500000 371.590000 ;
      RECT 907.500000 370.410000 908.500000 371.590000 ;
      RECT 866.500000 370.410000 899.500000 371.590000 ;
      RECT 857.500000 370.410000 858.500000 371.590000 ;
      RECT 816.500000 370.410000 849.500000 371.590000 ;
      RECT 807.500000 370.410000 808.500000 371.590000 ;
      RECT 766.500000 370.410000 799.500000 371.590000 ;
      RECT 757.500000 370.410000 758.500000 371.590000 ;
      RECT 716.500000 370.410000 749.500000 371.590000 ;
      RECT 707.500000 370.410000 708.500000 371.590000 ;
      RECT 666.500000 370.410000 699.500000 371.590000 ;
      RECT 657.500000 370.410000 658.500000 371.590000 ;
      RECT 616.500000 370.410000 649.500000 371.590000 ;
      RECT 607.500000 370.410000 608.500000 371.590000 ;
      RECT 566.500000 370.410000 599.500000 371.590000 ;
      RECT 557.500000 370.410000 558.500000 371.590000 ;
      RECT 516.500000 370.410000 549.500000 371.590000 ;
      RECT 507.500000 370.410000 508.500000 371.590000 ;
      RECT 466.500000 370.410000 499.500000 371.590000 ;
      RECT 457.500000 370.410000 458.500000 371.590000 ;
      RECT 416.500000 370.410000 449.500000 371.590000 ;
      RECT 407.500000 370.410000 408.500000 371.590000 ;
      RECT 366.500000 370.410000 399.500000 371.590000 ;
      RECT 357.500000 370.410000 358.500000 371.590000 ;
      RECT 316.500000 370.410000 349.500000 371.590000 ;
      RECT 307.500000 370.410000 308.500000 371.590000 ;
      RECT 266.500000 370.410000 299.500000 371.590000 ;
      RECT 257.500000 370.410000 258.500000 371.590000 ;
      RECT 216.500000 370.410000 249.500000 371.590000 ;
      RECT 207.500000 370.410000 208.500000 371.590000 ;
      RECT 166.500000 370.410000 199.500000 371.590000 ;
      RECT 157.500000 370.410000 158.500000 371.590000 ;
      RECT 116.500000 370.410000 149.500000 371.590000 ;
      RECT 107.500000 370.410000 108.500000 371.590000 ;
      RECT 66.500000 370.410000 99.500000 371.590000 ;
      RECT 57.500000 370.410000 58.500000 371.590000 ;
      RECT 29.500000 370.410000 49.500000 371.590000 ;
      RECT 15.500000 370.410000 16.500000 371.590000 ;
      RECT 1157.500000 369.590000 1170.500000 370.410000 ;
      RECT 1107.500000 369.590000 1149.500000 370.410000 ;
      RECT 1057.500000 369.590000 1099.500000 370.410000 ;
      RECT 1007.500000 369.590000 1049.500000 370.410000 ;
      RECT 957.500000 369.590000 999.500000 370.410000 ;
      RECT 907.500000 369.590000 949.500000 370.410000 ;
      RECT 857.500000 369.590000 899.500000 370.410000 ;
      RECT 807.500000 369.590000 849.500000 370.410000 ;
      RECT 757.500000 369.590000 799.500000 370.410000 ;
      RECT 707.500000 369.590000 749.500000 370.410000 ;
      RECT 657.500000 369.590000 699.500000 370.410000 ;
      RECT 607.500000 369.590000 649.500000 370.410000 ;
      RECT 557.500000 369.590000 599.500000 370.410000 ;
      RECT 507.500000 369.590000 549.500000 370.410000 ;
      RECT 407.500000 369.590000 449.500000 370.410000 ;
      RECT 357.500000 369.590000 399.500000 370.410000 ;
      RECT 307.500000 369.590000 349.500000 370.410000 ;
      RECT 257.500000 369.590000 299.500000 370.410000 ;
      RECT 207.500000 369.590000 249.500000 370.410000 ;
      RECT 157.500000 369.590000 199.500000 370.410000 ;
      RECT 107.500000 369.590000 149.500000 370.410000 ;
      RECT 57.500000 369.590000 99.500000 370.410000 ;
      RECT 15.500000 369.590000 49.500000 370.410000 ;
      RECT 1183.500000 368.410000 1186.000000 371.590000 ;
      RECT 1169.500000 368.410000 1170.500000 369.590000 ;
      RECT 1116.500000 368.410000 1149.500000 369.590000 ;
      RECT 1107.500000 368.410000 1108.500000 369.590000 ;
      RECT 1066.500000 368.410000 1099.500000 369.590000 ;
      RECT 1057.500000 368.410000 1058.500000 369.590000 ;
      RECT 1016.500000 368.410000 1049.500000 369.590000 ;
      RECT 1007.500000 368.410000 1008.500000 369.590000 ;
      RECT 966.500000 368.410000 999.500000 369.590000 ;
      RECT 957.500000 368.410000 958.500000 369.590000 ;
      RECT 916.500000 368.410000 949.500000 369.590000 ;
      RECT 907.500000 368.410000 908.500000 369.590000 ;
      RECT 866.500000 368.410000 899.500000 369.590000 ;
      RECT 857.500000 368.410000 858.500000 369.590000 ;
      RECT 816.500000 368.410000 849.500000 369.590000 ;
      RECT 807.500000 368.410000 808.500000 369.590000 ;
      RECT 766.500000 368.410000 799.500000 369.590000 ;
      RECT 757.500000 368.410000 758.500000 369.590000 ;
      RECT 716.500000 368.410000 749.500000 369.590000 ;
      RECT 707.500000 368.410000 708.500000 369.590000 ;
      RECT 666.500000 368.410000 699.500000 369.590000 ;
      RECT 657.500000 368.410000 658.500000 369.590000 ;
      RECT 616.500000 368.410000 649.500000 369.590000 ;
      RECT 607.500000 368.410000 608.500000 369.590000 ;
      RECT 566.500000 368.410000 599.500000 369.590000 ;
      RECT 557.500000 368.410000 558.500000 369.590000 ;
      RECT 516.500000 368.410000 549.500000 369.590000 ;
      RECT 507.500000 368.410000 508.500000 369.590000 ;
      RECT 457.500000 368.410000 499.500000 370.410000 ;
      RECT 407.500000 368.410000 408.500000 369.590000 ;
      RECT 366.500000 368.410000 399.500000 369.590000 ;
      RECT 357.500000 368.410000 358.500000 369.590000 ;
      RECT 316.500000 368.410000 349.500000 369.590000 ;
      RECT 307.500000 368.410000 308.500000 369.590000 ;
      RECT 266.500000 368.410000 299.500000 369.590000 ;
      RECT 257.500000 368.410000 258.500000 369.590000 ;
      RECT 216.500000 368.410000 249.500000 369.590000 ;
      RECT 207.500000 368.410000 208.500000 369.590000 ;
      RECT 166.500000 368.410000 199.500000 369.590000 ;
      RECT 157.500000 368.410000 158.500000 369.590000 ;
      RECT 116.500000 368.410000 149.500000 369.590000 ;
      RECT 107.500000 368.410000 108.500000 369.590000 ;
      RECT 66.500000 368.410000 99.500000 369.590000 ;
      RECT 57.500000 368.410000 58.500000 369.590000 ;
      RECT 29.500000 368.410000 49.500000 369.590000 ;
      RECT 15.500000 368.410000 16.500000 369.590000 ;
      RECT 0.000000 368.410000 2.500000 371.590000 ;
      RECT 1169.500000 367.590000 1186.000000 368.410000 ;
      RECT 1116.500000 367.590000 1156.500000 368.410000 ;
      RECT 1066.500000 367.590000 1108.500000 368.410000 ;
      RECT 1016.500000 367.590000 1058.500000 368.410000 ;
      RECT 966.500000 367.590000 1008.500000 368.410000 ;
      RECT 916.500000 367.590000 958.500000 368.410000 ;
      RECT 866.500000 367.590000 908.500000 368.410000 ;
      RECT 816.500000 367.590000 858.500000 368.410000 ;
      RECT 766.500000 367.590000 808.500000 368.410000 ;
      RECT 716.500000 367.590000 758.500000 368.410000 ;
      RECT 666.500000 367.590000 708.500000 368.410000 ;
      RECT 616.500000 367.590000 658.500000 368.410000 ;
      RECT 566.500000 367.590000 608.500000 368.410000 ;
      RECT 516.500000 367.590000 558.500000 368.410000 ;
      RECT 457.500000 367.590000 508.500000 368.410000 ;
      RECT 366.500000 367.590000 408.500000 368.410000 ;
      RECT 316.500000 367.590000 358.500000 368.410000 ;
      RECT 266.500000 367.590000 308.500000 368.410000 ;
      RECT 216.500000 367.590000 258.500000 368.410000 ;
      RECT 166.500000 367.590000 208.500000 368.410000 ;
      RECT 116.500000 367.590000 158.500000 368.410000 ;
      RECT 66.500000 367.590000 108.500000 368.410000 ;
      RECT 29.500000 367.590000 58.500000 368.410000 ;
      RECT 0.000000 367.590000 16.500000 368.410000 ;
      RECT 1169.500000 366.410000 1170.500000 367.590000 ;
      RECT 1116.500000 366.410000 1149.500000 367.590000 ;
      RECT 1107.500000 366.410000 1108.500000 367.590000 ;
      RECT 1066.500000 366.410000 1099.500000 367.590000 ;
      RECT 1057.500000 366.410000 1058.500000 367.590000 ;
      RECT 1016.500000 366.410000 1049.500000 367.590000 ;
      RECT 1007.500000 366.410000 1008.500000 367.590000 ;
      RECT 966.500000 366.410000 999.500000 367.590000 ;
      RECT 957.500000 366.410000 958.500000 367.590000 ;
      RECT 916.500000 366.410000 949.500000 367.590000 ;
      RECT 907.500000 366.410000 908.500000 367.590000 ;
      RECT 866.500000 366.410000 899.500000 367.590000 ;
      RECT 857.500000 366.410000 858.500000 367.590000 ;
      RECT 816.500000 366.410000 849.500000 367.590000 ;
      RECT 807.500000 366.410000 808.500000 367.590000 ;
      RECT 766.500000 366.410000 799.500000 367.590000 ;
      RECT 757.500000 366.410000 758.500000 367.590000 ;
      RECT 716.500000 366.410000 749.500000 367.590000 ;
      RECT 707.500000 366.410000 708.500000 367.590000 ;
      RECT 666.500000 366.410000 699.500000 367.590000 ;
      RECT 657.500000 366.410000 658.500000 367.590000 ;
      RECT 616.500000 366.410000 649.500000 367.590000 ;
      RECT 607.500000 366.410000 608.500000 367.590000 ;
      RECT 566.500000 366.410000 599.500000 367.590000 ;
      RECT 557.500000 366.410000 558.500000 367.590000 ;
      RECT 516.500000 366.410000 549.500000 367.590000 ;
      RECT 507.500000 366.410000 508.500000 367.590000 ;
      RECT 416.500000 366.410000 449.500000 369.590000 ;
      RECT 407.500000 366.410000 408.500000 367.590000 ;
      RECT 366.500000 366.410000 399.500000 367.590000 ;
      RECT 357.500000 366.410000 358.500000 367.590000 ;
      RECT 316.500000 366.410000 349.500000 367.590000 ;
      RECT 307.500000 366.410000 308.500000 367.590000 ;
      RECT 266.500000 366.410000 299.500000 367.590000 ;
      RECT 257.500000 366.410000 258.500000 367.590000 ;
      RECT 216.500000 366.410000 249.500000 367.590000 ;
      RECT 207.500000 366.410000 208.500000 367.590000 ;
      RECT 166.500000 366.410000 199.500000 367.590000 ;
      RECT 157.500000 366.410000 158.500000 367.590000 ;
      RECT 116.500000 366.410000 149.500000 367.590000 ;
      RECT 107.500000 366.410000 108.500000 367.590000 ;
      RECT 66.500000 366.410000 99.500000 367.590000 ;
      RECT 57.500000 366.410000 58.500000 367.590000 ;
      RECT 29.500000 366.410000 49.500000 367.590000 ;
      RECT 15.500000 366.410000 16.500000 367.590000 ;
      RECT 1157.500000 365.590000 1170.500000 366.410000 ;
      RECT 1107.500000 365.590000 1149.500000 366.410000 ;
      RECT 1057.500000 365.590000 1099.500000 366.410000 ;
      RECT 1007.500000 365.590000 1049.500000 366.410000 ;
      RECT 957.500000 365.590000 999.500000 366.410000 ;
      RECT 907.500000 365.590000 949.500000 366.410000 ;
      RECT 857.500000 365.590000 899.500000 366.410000 ;
      RECT 807.500000 365.590000 849.500000 366.410000 ;
      RECT 757.500000 365.590000 799.500000 366.410000 ;
      RECT 707.500000 365.590000 749.500000 366.410000 ;
      RECT 657.500000 365.590000 699.500000 366.410000 ;
      RECT 607.500000 365.590000 649.500000 366.410000 ;
      RECT 557.500000 365.590000 599.500000 366.410000 ;
      RECT 507.500000 365.590000 549.500000 366.410000 ;
      RECT 407.500000 365.590000 449.500000 366.410000 ;
      RECT 357.500000 365.590000 399.500000 366.410000 ;
      RECT 307.500000 365.590000 349.500000 366.410000 ;
      RECT 257.500000 365.590000 299.500000 366.410000 ;
      RECT 207.500000 365.590000 249.500000 366.410000 ;
      RECT 157.500000 365.590000 199.500000 366.410000 ;
      RECT 107.500000 365.590000 149.500000 366.410000 ;
      RECT 57.500000 365.590000 99.500000 366.410000 ;
      RECT 15.500000 365.590000 49.500000 366.410000 ;
      RECT 457.500000 364.605000 499.500000 367.590000 ;
      RECT 416.500000 364.605000 449.500000 365.590000 ;
      RECT 1183.500000 364.410000 1186.000000 367.590000 ;
      RECT 1169.500000 364.410000 1170.500000 365.590000 ;
      RECT 1116.500000 364.410000 1149.500000 365.590000 ;
      RECT 1107.500000 364.410000 1108.500000 365.590000 ;
      RECT 1066.500000 364.410000 1099.500000 365.590000 ;
      RECT 1057.500000 364.410000 1058.500000 365.590000 ;
      RECT 1016.500000 364.410000 1049.500000 365.590000 ;
      RECT 1007.500000 364.410000 1008.500000 365.590000 ;
      RECT 966.500000 364.410000 999.500000 365.590000 ;
      RECT 957.500000 364.410000 958.500000 365.590000 ;
      RECT 916.500000 364.410000 949.500000 365.590000 ;
      RECT 907.500000 364.410000 908.500000 365.590000 ;
      RECT 866.500000 364.410000 899.500000 365.590000 ;
      RECT 857.500000 364.410000 858.500000 365.590000 ;
      RECT 816.500000 364.410000 849.500000 365.590000 ;
      RECT 807.500000 364.410000 808.500000 365.590000 ;
      RECT 766.500000 364.410000 799.500000 365.590000 ;
      RECT 757.500000 364.410000 758.500000 365.590000 ;
      RECT 716.500000 364.410000 749.500000 365.590000 ;
      RECT 707.500000 364.410000 708.500000 365.590000 ;
      RECT 666.500000 364.410000 699.500000 365.590000 ;
      RECT 657.500000 364.410000 658.500000 365.590000 ;
      RECT 616.500000 364.410000 649.500000 365.590000 ;
      RECT 607.500000 364.410000 608.500000 365.590000 ;
      RECT 566.500000 364.410000 599.500000 365.590000 ;
      RECT 557.500000 364.410000 558.500000 365.590000 ;
      RECT 516.500000 364.410000 549.500000 365.590000 ;
      RECT 507.500000 364.410000 508.500000 365.590000 ;
      RECT 416.500000 364.410000 499.500000 364.605000 ;
      RECT 407.500000 364.410000 408.500000 365.590000 ;
      RECT 366.500000 364.410000 399.500000 365.590000 ;
      RECT 357.500000 364.410000 358.500000 365.590000 ;
      RECT 316.500000 364.410000 349.500000 365.590000 ;
      RECT 307.500000 364.410000 308.500000 365.590000 ;
      RECT 266.500000 364.410000 299.500000 365.590000 ;
      RECT 257.500000 364.410000 258.500000 365.590000 ;
      RECT 216.500000 364.410000 249.500000 365.590000 ;
      RECT 207.500000 364.410000 208.500000 365.590000 ;
      RECT 166.500000 364.410000 199.500000 365.590000 ;
      RECT 157.500000 364.410000 158.500000 365.590000 ;
      RECT 116.500000 364.410000 149.500000 365.590000 ;
      RECT 107.500000 364.410000 108.500000 365.590000 ;
      RECT 66.500000 364.410000 99.500000 365.590000 ;
      RECT 57.500000 364.410000 58.500000 365.590000 ;
      RECT 29.500000 364.410000 49.500000 365.590000 ;
      RECT 15.500000 364.410000 16.500000 365.590000 ;
      RECT 0.000000 364.410000 2.500000 367.590000 ;
      RECT 1169.500000 363.590000 1186.000000 364.410000 ;
      RECT 1116.500000 363.590000 1156.500000 364.410000 ;
      RECT 1066.500000 363.590000 1108.500000 364.410000 ;
      RECT 1016.500000 363.590000 1058.500000 364.410000 ;
      RECT 966.500000 363.590000 1008.500000 364.410000 ;
      RECT 916.500000 363.590000 958.500000 364.410000 ;
      RECT 866.500000 363.590000 908.500000 364.410000 ;
      RECT 816.500000 363.590000 858.500000 364.410000 ;
      RECT 766.500000 363.590000 808.500000 364.410000 ;
      RECT 716.500000 363.590000 758.500000 364.410000 ;
      RECT 666.500000 363.590000 708.500000 364.410000 ;
      RECT 616.500000 363.590000 658.500000 364.410000 ;
      RECT 566.500000 363.590000 608.500000 364.410000 ;
      RECT 516.500000 363.590000 558.500000 364.410000 ;
      RECT 416.500000 363.590000 508.500000 364.410000 ;
      RECT 366.500000 363.590000 408.500000 364.410000 ;
      RECT 316.500000 363.590000 358.500000 364.410000 ;
      RECT 266.500000 363.590000 308.500000 364.410000 ;
      RECT 216.500000 363.590000 258.500000 364.410000 ;
      RECT 166.500000 363.590000 208.500000 364.410000 ;
      RECT 116.500000 363.590000 158.500000 364.410000 ;
      RECT 66.500000 363.590000 108.500000 364.410000 ;
      RECT 29.500000 363.590000 58.500000 364.410000 ;
      RECT 0.000000 363.590000 16.500000 364.410000 ;
      RECT 1169.500000 362.410000 1170.500000 363.590000 ;
      RECT 1116.500000 362.410000 1149.500000 363.590000 ;
      RECT 1107.500000 362.410000 1108.500000 363.590000 ;
      RECT 1066.500000 362.410000 1099.500000 363.590000 ;
      RECT 1057.500000 362.410000 1058.500000 363.590000 ;
      RECT 1016.500000 362.410000 1049.500000 363.590000 ;
      RECT 1007.500000 362.410000 1008.500000 363.590000 ;
      RECT 966.500000 362.410000 999.500000 363.590000 ;
      RECT 957.500000 362.410000 958.500000 363.590000 ;
      RECT 916.500000 362.410000 949.500000 363.590000 ;
      RECT 907.500000 362.410000 908.500000 363.590000 ;
      RECT 866.500000 362.410000 899.500000 363.590000 ;
      RECT 857.500000 362.410000 858.500000 363.590000 ;
      RECT 816.500000 362.410000 849.500000 363.590000 ;
      RECT 807.500000 362.410000 808.500000 363.590000 ;
      RECT 766.500000 362.410000 799.500000 363.590000 ;
      RECT 757.500000 362.410000 758.500000 363.590000 ;
      RECT 716.500000 362.410000 749.500000 363.590000 ;
      RECT 707.500000 362.410000 708.500000 363.590000 ;
      RECT 666.500000 362.410000 699.500000 363.590000 ;
      RECT 657.500000 362.410000 658.500000 363.590000 ;
      RECT 616.500000 362.410000 649.500000 363.590000 ;
      RECT 607.500000 362.410000 608.500000 363.590000 ;
      RECT 566.500000 362.410000 599.500000 363.590000 ;
      RECT 557.500000 362.410000 558.500000 363.590000 ;
      RECT 516.500000 362.410000 549.500000 363.590000 ;
      RECT 507.500000 362.410000 508.500000 363.590000 ;
      RECT 416.500000 362.410000 499.500000 363.590000 ;
      RECT 407.500000 362.410000 408.500000 363.590000 ;
      RECT 366.500000 362.410000 399.500000 363.590000 ;
      RECT 357.500000 362.410000 358.500000 363.590000 ;
      RECT 316.500000 362.410000 349.500000 363.590000 ;
      RECT 307.500000 362.410000 308.500000 363.590000 ;
      RECT 266.500000 362.410000 299.500000 363.590000 ;
      RECT 257.500000 362.410000 258.500000 363.590000 ;
      RECT 216.500000 362.410000 249.500000 363.590000 ;
      RECT 207.500000 362.410000 208.500000 363.590000 ;
      RECT 166.500000 362.410000 199.500000 363.590000 ;
      RECT 157.500000 362.410000 158.500000 363.590000 ;
      RECT 116.500000 362.410000 149.500000 363.590000 ;
      RECT 107.500000 362.410000 108.500000 363.590000 ;
      RECT 66.500000 362.410000 99.500000 363.590000 ;
      RECT 57.500000 362.410000 58.500000 363.590000 ;
      RECT 29.500000 362.410000 49.500000 363.590000 ;
      RECT 15.500000 362.410000 16.500000 363.590000 ;
      RECT 1157.500000 361.590000 1170.500000 362.410000 ;
      RECT 1107.500000 361.590000 1149.500000 362.410000 ;
      RECT 1057.500000 361.590000 1099.500000 362.410000 ;
      RECT 1007.500000 361.590000 1049.500000 362.410000 ;
      RECT 957.500000 361.590000 999.500000 362.410000 ;
      RECT 907.500000 361.590000 949.500000 362.410000 ;
      RECT 857.500000 361.590000 899.500000 362.410000 ;
      RECT 807.500000 361.590000 849.500000 362.410000 ;
      RECT 757.500000 361.590000 799.500000 362.410000 ;
      RECT 707.500000 361.590000 749.500000 362.410000 ;
      RECT 657.500000 361.590000 699.500000 362.410000 ;
      RECT 607.500000 361.590000 649.500000 362.410000 ;
      RECT 557.500000 361.590000 599.500000 362.410000 ;
      RECT 507.500000 361.590000 549.500000 362.410000 ;
      RECT 407.500000 361.590000 499.500000 362.410000 ;
      RECT 357.500000 361.590000 399.500000 362.410000 ;
      RECT 307.500000 361.590000 349.500000 362.410000 ;
      RECT 257.500000 361.590000 299.500000 362.410000 ;
      RECT 207.500000 361.590000 249.500000 362.410000 ;
      RECT 157.500000 361.590000 199.500000 362.410000 ;
      RECT 107.500000 361.590000 149.500000 362.410000 ;
      RECT 15.500000 361.590000 49.500000 362.410000 ;
      RECT 1183.500000 360.410000 1186.000000 363.590000 ;
      RECT 1169.500000 360.410000 1170.500000 361.590000 ;
      RECT 1116.500000 360.410000 1149.500000 361.590000 ;
      RECT 1107.500000 360.410000 1108.500000 361.590000 ;
      RECT 1066.500000 360.410000 1099.500000 361.590000 ;
      RECT 1057.500000 360.410000 1058.500000 361.590000 ;
      RECT 1016.500000 360.410000 1049.500000 361.590000 ;
      RECT 1007.500000 360.410000 1008.500000 361.590000 ;
      RECT 966.500000 360.410000 999.500000 361.590000 ;
      RECT 957.500000 360.410000 958.500000 361.590000 ;
      RECT 916.500000 360.410000 949.500000 361.590000 ;
      RECT 907.500000 360.410000 908.500000 361.590000 ;
      RECT 866.500000 360.410000 899.500000 361.590000 ;
      RECT 857.500000 360.410000 858.500000 361.590000 ;
      RECT 816.500000 360.410000 849.500000 361.590000 ;
      RECT 807.500000 360.410000 808.500000 361.590000 ;
      RECT 766.500000 360.410000 799.500000 361.590000 ;
      RECT 757.500000 360.410000 758.500000 361.590000 ;
      RECT 716.500000 360.410000 749.500000 361.590000 ;
      RECT 707.500000 360.410000 708.500000 361.590000 ;
      RECT 666.500000 360.410000 699.500000 361.590000 ;
      RECT 657.500000 360.410000 658.500000 361.590000 ;
      RECT 616.500000 360.410000 649.500000 361.590000 ;
      RECT 607.500000 360.410000 608.500000 361.590000 ;
      RECT 566.500000 360.410000 599.500000 361.590000 ;
      RECT 557.500000 360.410000 558.500000 361.590000 ;
      RECT 516.500000 360.410000 549.500000 361.590000 ;
      RECT 507.500000 360.410000 508.500000 361.590000 ;
      RECT 416.500000 360.410000 499.500000 361.590000 ;
      RECT 407.500000 360.410000 408.500000 361.590000 ;
      RECT 366.500000 360.410000 399.500000 361.590000 ;
      RECT 357.500000 360.410000 358.500000 361.590000 ;
      RECT 316.500000 360.410000 349.500000 361.590000 ;
      RECT 307.500000 360.410000 308.500000 361.590000 ;
      RECT 266.500000 360.410000 299.500000 361.590000 ;
      RECT 257.500000 360.410000 258.500000 361.590000 ;
      RECT 216.500000 360.410000 249.500000 361.590000 ;
      RECT 207.500000 360.410000 208.500000 361.590000 ;
      RECT 166.500000 360.410000 199.500000 361.590000 ;
      RECT 157.500000 360.410000 158.500000 361.590000 ;
      RECT 116.500000 360.410000 149.500000 361.590000 ;
      RECT 107.500000 360.410000 108.500000 361.590000 ;
      RECT 57.500000 360.410000 99.500000 362.410000 ;
      RECT 29.500000 360.410000 49.500000 361.590000 ;
      RECT 15.500000 360.410000 16.500000 361.590000 ;
      RECT 0.000000 360.410000 2.500000 363.590000 ;
      RECT 1169.500000 359.590000 1186.000000 360.410000 ;
      RECT 1116.500000 359.590000 1156.500000 360.410000 ;
      RECT 1066.500000 359.590000 1108.500000 360.410000 ;
      RECT 1016.500000 359.590000 1058.500000 360.410000 ;
      RECT 966.500000 359.590000 1008.500000 360.410000 ;
      RECT 916.500000 359.590000 958.500000 360.410000 ;
      RECT 866.500000 359.590000 908.500000 360.410000 ;
      RECT 816.500000 359.590000 858.500000 360.410000 ;
      RECT 766.500000 359.590000 808.500000 360.410000 ;
      RECT 716.500000 359.590000 758.500000 360.410000 ;
      RECT 666.500000 359.590000 708.500000 360.410000 ;
      RECT 616.500000 359.590000 658.500000 360.410000 ;
      RECT 566.500000 359.590000 608.500000 360.410000 ;
      RECT 516.500000 359.590000 558.500000 360.410000 ;
      RECT 416.500000 359.590000 508.500000 360.410000 ;
      RECT 366.500000 359.590000 408.500000 360.410000 ;
      RECT 316.500000 359.590000 358.500000 360.410000 ;
      RECT 266.500000 359.590000 308.500000 360.410000 ;
      RECT 216.500000 359.590000 258.500000 360.410000 ;
      RECT 166.500000 359.590000 208.500000 360.410000 ;
      RECT 116.500000 359.590000 158.500000 360.410000 ;
      RECT 29.500000 359.590000 108.500000 360.410000 ;
      RECT 0.000000 359.590000 16.500000 360.410000 ;
      RECT 1169.500000 358.410000 1170.500000 359.590000 ;
      RECT 1116.500000 358.410000 1149.500000 359.590000 ;
      RECT 1107.500000 358.410000 1108.500000 359.590000 ;
      RECT 1066.500000 358.410000 1099.500000 359.590000 ;
      RECT 1057.500000 358.410000 1058.500000 359.590000 ;
      RECT 1016.500000 358.410000 1049.500000 359.590000 ;
      RECT 1007.500000 358.410000 1008.500000 359.590000 ;
      RECT 966.500000 358.410000 999.500000 359.590000 ;
      RECT 957.500000 358.410000 958.500000 359.590000 ;
      RECT 916.500000 358.410000 949.500000 359.590000 ;
      RECT 907.500000 358.410000 908.500000 359.590000 ;
      RECT 866.500000 358.410000 899.500000 359.590000 ;
      RECT 857.500000 358.410000 858.500000 359.590000 ;
      RECT 816.500000 358.410000 849.500000 359.590000 ;
      RECT 807.500000 358.410000 808.500000 359.590000 ;
      RECT 766.500000 358.410000 799.500000 359.590000 ;
      RECT 757.500000 358.410000 758.500000 359.590000 ;
      RECT 716.500000 358.410000 749.500000 359.590000 ;
      RECT 707.500000 358.410000 708.500000 359.590000 ;
      RECT 666.500000 358.410000 699.500000 359.590000 ;
      RECT 657.500000 358.410000 658.500000 359.590000 ;
      RECT 616.500000 358.410000 649.500000 359.590000 ;
      RECT 607.500000 358.410000 608.500000 359.590000 ;
      RECT 566.500000 358.410000 599.500000 359.590000 ;
      RECT 557.500000 358.410000 558.500000 359.590000 ;
      RECT 516.500000 358.410000 549.500000 359.590000 ;
      RECT 507.500000 358.410000 508.500000 359.590000 ;
      RECT 416.500000 358.410000 499.500000 359.590000 ;
      RECT 407.500000 358.410000 408.500000 359.590000 ;
      RECT 366.500000 358.410000 399.500000 359.590000 ;
      RECT 357.500000 358.410000 358.500000 359.590000 ;
      RECT 316.500000 358.410000 349.500000 359.590000 ;
      RECT 307.500000 358.410000 308.500000 359.590000 ;
      RECT 266.500000 358.410000 299.500000 359.590000 ;
      RECT 257.500000 358.410000 258.500000 359.590000 ;
      RECT 216.500000 358.410000 249.500000 359.590000 ;
      RECT 207.500000 358.410000 208.500000 359.590000 ;
      RECT 166.500000 358.410000 199.500000 359.590000 ;
      RECT 157.500000 358.410000 158.500000 359.590000 ;
      RECT 116.500000 358.410000 149.500000 359.590000 ;
      RECT 107.500000 358.410000 108.500000 359.590000 ;
      RECT 29.500000 358.410000 99.500000 359.590000 ;
      RECT 15.500000 358.410000 16.500000 359.590000 ;
      RECT 1157.500000 357.590000 1170.500000 358.410000 ;
      RECT 1107.500000 357.590000 1149.500000 358.410000 ;
      RECT 1057.500000 357.590000 1099.500000 358.410000 ;
      RECT 1007.500000 357.590000 1049.500000 358.410000 ;
      RECT 957.500000 357.590000 999.500000 358.410000 ;
      RECT 907.500000 357.590000 949.500000 358.410000 ;
      RECT 857.500000 357.590000 899.500000 358.410000 ;
      RECT 807.500000 357.590000 849.500000 358.410000 ;
      RECT 757.500000 357.590000 799.500000 358.410000 ;
      RECT 707.500000 357.590000 749.500000 358.410000 ;
      RECT 657.500000 357.590000 699.500000 358.410000 ;
      RECT 607.500000 357.590000 649.500000 358.410000 ;
      RECT 557.500000 357.590000 599.500000 358.410000 ;
      RECT 507.500000 357.590000 549.500000 358.410000 ;
      RECT 407.500000 357.590000 499.500000 358.410000 ;
      RECT 357.500000 357.590000 399.500000 358.410000 ;
      RECT 307.500000 357.590000 349.500000 358.410000 ;
      RECT 257.500000 357.590000 299.500000 358.410000 ;
      RECT 207.500000 357.590000 249.500000 358.410000 ;
      RECT 157.500000 357.590000 199.500000 358.410000 ;
      RECT 107.500000 357.590000 149.500000 358.410000 ;
      RECT 15.500000 357.590000 99.500000 358.410000 ;
      RECT 1183.500000 356.410000 1186.000000 359.590000 ;
      RECT 1169.500000 356.410000 1170.500000 357.590000 ;
      RECT 1116.500000 356.410000 1149.500000 357.590000 ;
      RECT 1107.500000 356.410000 1108.500000 357.590000 ;
      RECT 1066.500000 356.410000 1099.500000 357.590000 ;
      RECT 1057.500000 356.410000 1058.500000 357.590000 ;
      RECT 1016.500000 356.410000 1049.500000 357.590000 ;
      RECT 1007.500000 356.410000 1008.500000 357.590000 ;
      RECT 966.500000 356.410000 999.500000 357.590000 ;
      RECT 957.500000 356.410000 958.500000 357.590000 ;
      RECT 916.500000 356.410000 949.500000 357.590000 ;
      RECT 907.500000 356.410000 908.500000 357.590000 ;
      RECT 866.500000 356.410000 899.500000 357.590000 ;
      RECT 857.500000 356.410000 858.500000 357.590000 ;
      RECT 816.500000 356.410000 849.500000 357.590000 ;
      RECT 807.500000 356.410000 808.500000 357.590000 ;
      RECT 766.500000 356.410000 799.500000 357.590000 ;
      RECT 757.500000 356.410000 758.500000 357.590000 ;
      RECT 716.500000 356.410000 749.500000 357.590000 ;
      RECT 707.500000 356.410000 708.500000 357.590000 ;
      RECT 666.500000 356.410000 699.500000 357.590000 ;
      RECT 657.500000 356.410000 658.500000 357.590000 ;
      RECT 616.500000 356.410000 649.500000 357.590000 ;
      RECT 607.500000 356.410000 608.500000 357.590000 ;
      RECT 566.500000 356.410000 599.500000 357.590000 ;
      RECT 557.500000 356.410000 558.500000 357.590000 ;
      RECT 516.500000 356.410000 549.500000 357.590000 ;
      RECT 507.500000 356.410000 508.500000 357.590000 ;
      RECT 416.500000 356.410000 499.500000 357.590000 ;
      RECT 407.500000 356.410000 408.500000 357.590000 ;
      RECT 366.500000 356.410000 399.500000 357.590000 ;
      RECT 357.500000 356.410000 358.500000 357.590000 ;
      RECT 316.500000 356.410000 349.500000 357.590000 ;
      RECT 307.500000 356.410000 308.500000 357.590000 ;
      RECT 266.500000 356.410000 299.500000 357.590000 ;
      RECT 257.500000 356.410000 258.500000 357.590000 ;
      RECT 216.500000 356.410000 249.500000 357.590000 ;
      RECT 207.500000 356.410000 208.500000 357.590000 ;
      RECT 166.500000 356.410000 199.500000 357.590000 ;
      RECT 157.500000 356.410000 158.500000 357.590000 ;
      RECT 116.500000 356.410000 149.500000 357.590000 ;
      RECT 107.500000 356.410000 108.500000 357.590000 ;
      RECT 29.500000 356.410000 99.500000 357.590000 ;
      RECT 15.500000 356.410000 16.500000 357.590000 ;
      RECT 0.000000 356.410000 2.500000 359.590000 ;
      RECT 29.500000 356.245000 108.500000 356.410000 ;
      RECT 1169.500000 355.590000 1186.000000 356.410000 ;
      RECT 1116.500000 355.590000 1156.500000 356.410000 ;
      RECT 1066.500000 355.590000 1108.500000 356.410000 ;
      RECT 1016.500000 355.590000 1058.500000 356.410000 ;
      RECT 966.500000 355.590000 1008.500000 356.410000 ;
      RECT 916.500000 355.590000 958.500000 356.410000 ;
      RECT 866.500000 355.590000 908.500000 356.410000 ;
      RECT 816.500000 355.590000 858.500000 356.410000 ;
      RECT 766.500000 355.590000 808.500000 356.410000 ;
      RECT 716.500000 355.590000 758.500000 356.410000 ;
      RECT 666.500000 355.590000 708.500000 356.410000 ;
      RECT 616.500000 355.590000 658.500000 356.410000 ;
      RECT 566.500000 355.590000 608.500000 356.410000 ;
      RECT 516.500000 355.590000 558.500000 356.410000 ;
      RECT 416.500000 355.590000 508.500000 356.410000 ;
      RECT 366.500000 355.590000 408.500000 356.410000 ;
      RECT 316.500000 355.590000 358.500000 356.410000 ;
      RECT 266.500000 355.590000 308.500000 356.410000 ;
      RECT 216.500000 355.590000 258.500000 356.410000 ;
      RECT 166.500000 355.590000 208.500000 356.410000 ;
      RECT 116.500000 355.590000 158.500000 356.410000 ;
      RECT 57.500000 355.590000 108.500000 356.245000 ;
      RECT 0.000000 355.590000 16.500000 356.410000 ;
      RECT 1169.500000 354.410000 1170.500000 355.590000 ;
      RECT 1116.500000 354.410000 1149.500000 355.590000 ;
      RECT 1107.500000 354.410000 1108.500000 355.590000 ;
      RECT 1066.500000 354.410000 1099.500000 355.590000 ;
      RECT 1057.500000 354.410000 1058.500000 355.590000 ;
      RECT 1016.500000 354.410000 1049.500000 355.590000 ;
      RECT 1007.500000 354.410000 1008.500000 355.590000 ;
      RECT 966.500000 354.410000 999.500000 355.590000 ;
      RECT 957.500000 354.410000 958.500000 355.590000 ;
      RECT 916.500000 354.410000 949.500000 355.590000 ;
      RECT 907.500000 354.410000 908.500000 355.590000 ;
      RECT 866.500000 354.410000 899.500000 355.590000 ;
      RECT 857.500000 354.410000 858.500000 355.590000 ;
      RECT 816.500000 354.410000 849.500000 355.590000 ;
      RECT 807.500000 354.410000 808.500000 355.590000 ;
      RECT 766.500000 354.410000 799.500000 355.590000 ;
      RECT 757.500000 354.410000 758.500000 355.590000 ;
      RECT 716.500000 354.410000 749.500000 355.590000 ;
      RECT 707.500000 354.410000 708.500000 355.590000 ;
      RECT 666.500000 354.410000 699.500000 355.590000 ;
      RECT 657.500000 354.410000 658.500000 355.590000 ;
      RECT 616.500000 354.410000 649.500000 355.590000 ;
      RECT 607.500000 354.410000 608.500000 355.590000 ;
      RECT 566.500000 354.410000 599.500000 355.590000 ;
      RECT 557.500000 354.410000 558.500000 355.590000 ;
      RECT 516.500000 354.410000 549.500000 355.590000 ;
      RECT 507.500000 354.410000 508.500000 355.590000 ;
      RECT 416.500000 354.410000 499.500000 355.590000 ;
      RECT 407.500000 354.410000 408.500000 355.590000 ;
      RECT 366.500000 354.410000 399.500000 355.590000 ;
      RECT 357.500000 354.410000 358.500000 355.590000 ;
      RECT 316.500000 354.410000 349.500000 355.590000 ;
      RECT 307.500000 354.410000 308.500000 355.590000 ;
      RECT 266.500000 354.410000 299.500000 355.590000 ;
      RECT 257.500000 354.410000 258.500000 355.590000 ;
      RECT 216.500000 354.410000 249.500000 355.590000 ;
      RECT 207.500000 354.410000 208.500000 355.590000 ;
      RECT 166.500000 354.410000 199.500000 355.590000 ;
      RECT 157.500000 354.410000 158.500000 355.590000 ;
      RECT 116.500000 354.410000 149.500000 355.590000 ;
      RECT 107.500000 354.410000 108.500000 355.590000 ;
      RECT 29.500000 354.410000 49.500000 356.245000 ;
      RECT 15.500000 354.410000 16.500000 355.590000 ;
      RECT 57.500000 354.245000 99.500000 355.590000 ;
      RECT 407.500000 353.730000 499.500000 354.410000 ;
      RECT 1157.500000 353.590000 1170.500000 354.410000 ;
      RECT 1107.500000 353.590000 1149.500000 354.410000 ;
      RECT 1057.500000 353.590000 1099.500000 354.410000 ;
      RECT 1007.500000 353.590000 1049.500000 354.410000 ;
      RECT 957.500000 353.590000 999.500000 354.410000 ;
      RECT 907.500000 353.590000 949.500000 354.410000 ;
      RECT 857.500000 353.590000 899.500000 354.410000 ;
      RECT 807.500000 353.590000 849.500000 354.410000 ;
      RECT 757.500000 353.590000 799.500000 354.410000 ;
      RECT 707.500000 353.590000 749.500000 354.410000 ;
      RECT 657.500000 353.590000 699.500000 354.410000 ;
      RECT 607.500000 353.590000 649.500000 354.410000 ;
      RECT 557.500000 353.590000 599.500000 354.410000 ;
      RECT 507.500000 353.590000 549.500000 354.410000 ;
      RECT 407.500000 353.590000 458.500000 353.730000 ;
      RECT 357.500000 353.590000 399.500000 354.410000 ;
      RECT 307.500000 353.590000 349.500000 354.410000 ;
      RECT 257.500000 353.590000 299.500000 354.410000 ;
      RECT 207.500000 353.590000 249.500000 354.410000 ;
      RECT 157.500000 353.590000 199.500000 354.410000 ;
      RECT 107.500000 353.590000 149.500000 354.410000 ;
      RECT 15.500000 353.590000 49.500000 354.410000 ;
      RECT 57.500000 352.945000 58.500000 354.245000 ;
      RECT 29.500000 352.945000 49.500000 353.590000 ;
      RECT 1183.500000 352.410000 1186.000000 355.590000 ;
      RECT 1169.500000 352.410000 1170.500000 353.590000 ;
      RECT 1116.500000 352.410000 1149.500000 353.590000 ;
      RECT 1107.500000 352.410000 1108.500000 353.590000 ;
      RECT 1066.500000 352.410000 1099.500000 353.590000 ;
      RECT 1057.500000 352.410000 1058.500000 353.590000 ;
      RECT 1016.500000 352.410000 1049.500000 353.590000 ;
      RECT 1007.500000 352.410000 1008.500000 353.590000 ;
      RECT 966.500000 352.410000 999.500000 353.590000 ;
      RECT 957.500000 352.410000 958.500000 353.590000 ;
      RECT 916.500000 352.410000 949.500000 353.590000 ;
      RECT 907.500000 352.410000 908.500000 353.590000 ;
      RECT 866.500000 352.410000 899.500000 353.590000 ;
      RECT 857.500000 352.410000 858.500000 353.590000 ;
      RECT 816.500000 352.410000 849.500000 353.590000 ;
      RECT 807.500000 352.410000 808.500000 353.590000 ;
      RECT 766.500000 352.410000 799.500000 353.590000 ;
      RECT 757.500000 352.410000 758.500000 353.590000 ;
      RECT 716.500000 352.410000 749.500000 353.590000 ;
      RECT 707.500000 352.410000 708.500000 353.590000 ;
      RECT 666.500000 352.410000 699.500000 353.590000 ;
      RECT 657.500000 352.410000 658.500000 353.590000 ;
      RECT 616.500000 352.410000 649.500000 353.590000 ;
      RECT 607.500000 352.410000 608.500000 353.590000 ;
      RECT 566.500000 352.410000 599.500000 353.590000 ;
      RECT 557.500000 352.410000 558.500000 353.590000 ;
      RECT 516.500000 352.410000 549.500000 353.590000 ;
      RECT 507.500000 352.410000 508.500000 353.590000 ;
      RECT 466.500000 352.410000 499.500000 353.730000 ;
      RECT 407.500000 352.410000 408.500000 353.590000 ;
      RECT 366.500000 352.410000 399.500000 353.590000 ;
      RECT 357.500000 352.410000 358.500000 353.590000 ;
      RECT 316.500000 352.410000 349.500000 353.590000 ;
      RECT 307.500000 352.410000 308.500000 353.590000 ;
      RECT 266.500000 352.410000 299.500000 353.590000 ;
      RECT 257.500000 352.410000 258.500000 353.590000 ;
      RECT 216.500000 352.410000 249.500000 353.590000 ;
      RECT 207.500000 352.410000 208.500000 353.590000 ;
      RECT 166.500000 352.410000 199.500000 353.590000 ;
      RECT 157.500000 352.410000 158.500000 353.590000 ;
      RECT 116.500000 352.410000 149.500000 353.590000 ;
      RECT 107.500000 352.410000 108.500000 353.590000 ;
      RECT 65.580000 352.410000 99.500000 354.245000 ;
      RECT 15.500000 352.410000 16.500000 353.590000 ;
      RECT 0.000000 352.410000 2.500000 355.590000 ;
      RECT 1169.500000 351.590000 1186.000000 352.410000 ;
      RECT 1116.500000 351.590000 1156.500000 352.410000 ;
      RECT 1066.500000 351.590000 1108.500000 352.410000 ;
      RECT 1016.500000 351.590000 1058.500000 352.410000 ;
      RECT 966.500000 351.590000 1008.500000 352.410000 ;
      RECT 916.500000 351.590000 958.500000 352.410000 ;
      RECT 866.500000 351.590000 908.500000 352.410000 ;
      RECT 816.500000 351.590000 858.500000 352.410000 ;
      RECT 766.500000 351.590000 808.500000 352.410000 ;
      RECT 716.500000 351.590000 758.500000 352.410000 ;
      RECT 666.500000 351.590000 708.500000 352.410000 ;
      RECT 616.500000 351.590000 658.500000 352.410000 ;
      RECT 566.500000 351.590000 608.500000 352.410000 ;
      RECT 516.500000 351.590000 558.500000 352.410000 ;
      RECT 466.500000 351.590000 508.500000 352.410000 ;
      RECT 366.500000 351.590000 408.500000 352.410000 ;
      RECT 316.500000 351.590000 358.500000 352.410000 ;
      RECT 266.500000 351.590000 308.500000 352.410000 ;
      RECT 216.500000 351.590000 258.500000 352.410000 ;
      RECT 166.500000 351.590000 208.500000 352.410000 ;
      RECT 116.500000 351.590000 158.500000 352.410000 ;
      RECT 65.580000 351.590000 108.500000 352.410000 ;
      RECT 0.000000 351.590000 16.500000 352.410000 ;
      RECT 65.580000 350.945000 99.500000 351.590000 ;
      RECT 29.500000 350.945000 58.500000 352.945000 ;
      RECT 1169.500000 350.410000 1170.500000 351.590000 ;
      RECT 1116.500000 350.410000 1149.500000 351.590000 ;
      RECT 1107.500000 350.410000 1108.500000 351.590000 ;
      RECT 1066.500000 350.410000 1099.500000 351.590000 ;
      RECT 1057.500000 350.410000 1058.500000 351.590000 ;
      RECT 1016.500000 350.410000 1049.500000 351.590000 ;
      RECT 1007.500000 350.410000 1008.500000 351.590000 ;
      RECT 966.500000 350.410000 999.500000 351.590000 ;
      RECT 957.500000 350.410000 958.500000 351.590000 ;
      RECT 916.500000 350.410000 949.500000 351.590000 ;
      RECT 907.500000 350.410000 908.500000 351.590000 ;
      RECT 866.500000 350.410000 899.500000 351.590000 ;
      RECT 857.500000 350.410000 858.500000 351.590000 ;
      RECT 816.500000 350.410000 849.500000 351.590000 ;
      RECT 807.500000 350.410000 808.500000 351.590000 ;
      RECT 766.500000 350.410000 799.500000 351.590000 ;
      RECT 757.500000 350.410000 758.500000 351.590000 ;
      RECT 716.500000 350.410000 749.500000 351.590000 ;
      RECT 707.500000 350.410000 708.500000 351.590000 ;
      RECT 666.500000 350.410000 699.500000 351.590000 ;
      RECT 657.500000 350.410000 658.500000 351.590000 ;
      RECT 616.500000 350.410000 649.500000 351.590000 ;
      RECT 607.500000 350.410000 608.500000 351.590000 ;
      RECT 566.500000 350.410000 599.500000 351.590000 ;
      RECT 557.500000 350.410000 558.500000 351.590000 ;
      RECT 516.500000 350.410000 549.500000 351.590000 ;
      RECT 507.500000 350.410000 508.500000 351.590000 ;
      RECT 416.500000 350.410000 458.500000 353.590000 ;
      RECT 407.500000 350.410000 408.500000 351.590000 ;
      RECT 366.500000 350.410000 399.500000 351.590000 ;
      RECT 357.500000 350.410000 358.500000 351.590000 ;
      RECT 316.500000 350.410000 349.500000 351.590000 ;
      RECT 307.500000 350.410000 308.500000 351.590000 ;
      RECT 266.500000 350.410000 299.500000 351.590000 ;
      RECT 257.500000 350.410000 258.500000 351.590000 ;
      RECT 216.500000 350.410000 249.500000 351.590000 ;
      RECT 207.500000 350.410000 208.500000 351.590000 ;
      RECT 166.500000 350.410000 199.500000 351.590000 ;
      RECT 157.500000 350.410000 158.500000 351.590000 ;
      RECT 116.500000 350.410000 149.500000 351.590000 ;
      RECT 107.500000 350.410000 108.500000 351.590000 ;
      RECT 29.500000 350.410000 99.500000 350.945000 ;
      RECT 15.500000 350.410000 16.500000 351.590000 ;
      RECT 466.500000 349.730000 499.500000 351.590000 ;
      RECT 407.500000 349.730000 458.500000 350.410000 ;
      RECT 1157.500000 349.590000 1170.500000 350.410000 ;
      RECT 1107.500000 349.590000 1149.500000 350.410000 ;
      RECT 1057.500000 349.590000 1099.500000 350.410000 ;
      RECT 1007.500000 349.590000 1049.500000 350.410000 ;
      RECT 957.500000 349.590000 999.500000 350.410000 ;
      RECT 907.500000 349.590000 949.500000 350.410000 ;
      RECT 857.500000 349.590000 899.500000 350.410000 ;
      RECT 807.500000 349.590000 849.500000 350.410000 ;
      RECT 757.500000 349.590000 799.500000 350.410000 ;
      RECT 707.500000 349.590000 749.500000 350.410000 ;
      RECT 657.500000 349.590000 699.500000 350.410000 ;
      RECT 607.500000 349.590000 649.500000 350.410000 ;
      RECT 557.500000 349.590000 599.500000 350.410000 ;
      RECT 507.500000 349.590000 549.500000 350.410000 ;
      RECT 407.500000 349.590000 499.500000 349.730000 ;
      RECT 357.500000 349.590000 399.500000 350.410000 ;
      RECT 307.500000 349.590000 349.500000 350.410000 ;
      RECT 257.500000 349.590000 299.500000 350.410000 ;
      RECT 207.500000 349.590000 249.500000 350.410000 ;
      RECT 157.500000 349.590000 199.500000 350.410000 ;
      RECT 107.500000 349.590000 149.500000 350.410000 ;
      RECT 15.500000 349.590000 99.500000 350.410000 ;
      RECT 1183.500000 348.410000 1186.000000 351.590000 ;
      RECT 1169.500000 348.410000 1170.500000 349.590000 ;
      RECT 1116.500000 348.410000 1149.500000 349.590000 ;
      RECT 1107.500000 348.410000 1108.500000 349.590000 ;
      RECT 1066.500000 348.410000 1099.500000 349.590000 ;
      RECT 1057.500000 348.410000 1058.500000 349.590000 ;
      RECT 1016.500000 348.410000 1049.500000 349.590000 ;
      RECT 1007.500000 348.410000 1008.500000 349.590000 ;
      RECT 966.500000 348.410000 999.500000 349.590000 ;
      RECT 957.500000 348.410000 958.500000 349.590000 ;
      RECT 916.500000 348.410000 949.500000 349.590000 ;
      RECT 907.500000 348.410000 908.500000 349.590000 ;
      RECT 866.500000 348.410000 899.500000 349.590000 ;
      RECT 857.500000 348.410000 858.500000 349.590000 ;
      RECT 816.500000 348.410000 849.500000 349.590000 ;
      RECT 807.500000 348.410000 808.500000 349.590000 ;
      RECT 766.500000 348.410000 799.500000 349.590000 ;
      RECT 757.500000 348.410000 758.500000 349.590000 ;
      RECT 716.500000 348.410000 749.500000 349.590000 ;
      RECT 707.500000 348.410000 708.500000 349.590000 ;
      RECT 666.500000 348.410000 699.500000 349.590000 ;
      RECT 657.500000 348.410000 658.500000 349.590000 ;
      RECT 616.500000 348.410000 649.500000 349.590000 ;
      RECT 607.500000 348.410000 608.500000 349.590000 ;
      RECT 566.500000 348.410000 599.500000 349.590000 ;
      RECT 557.500000 348.410000 558.500000 349.590000 ;
      RECT 516.500000 348.410000 549.500000 349.590000 ;
      RECT 507.500000 348.410000 508.500000 349.590000 ;
      RECT 466.500000 348.410000 499.500000 349.590000 ;
      RECT 407.500000 348.410000 408.500000 349.590000 ;
      RECT 366.500000 348.410000 399.500000 349.590000 ;
      RECT 357.500000 348.410000 358.500000 349.590000 ;
      RECT 316.500000 348.410000 349.500000 349.590000 ;
      RECT 307.500000 348.410000 308.500000 349.590000 ;
      RECT 266.500000 348.410000 299.500000 349.590000 ;
      RECT 257.500000 348.410000 258.500000 349.590000 ;
      RECT 216.500000 348.410000 249.500000 349.590000 ;
      RECT 207.500000 348.410000 208.500000 349.590000 ;
      RECT 166.500000 348.410000 199.500000 349.590000 ;
      RECT 157.500000 348.410000 158.500000 349.590000 ;
      RECT 116.500000 348.410000 149.500000 349.590000 ;
      RECT 107.500000 348.410000 108.500000 349.590000 ;
      RECT 66.500000 348.410000 99.500000 349.590000 ;
      RECT 15.500000 348.410000 16.500000 349.590000 ;
      RECT 0.000000 348.410000 2.500000 351.590000 ;
      RECT 1169.500000 347.590000 1186.000000 348.410000 ;
      RECT 1116.500000 347.590000 1156.500000 348.410000 ;
      RECT 1066.500000 347.590000 1108.500000 348.410000 ;
      RECT 1016.500000 347.590000 1058.500000 348.410000 ;
      RECT 966.500000 347.590000 1008.500000 348.410000 ;
      RECT 916.500000 347.590000 958.500000 348.410000 ;
      RECT 866.500000 347.590000 908.500000 348.410000 ;
      RECT 816.500000 347.590000 858.500000 348.410000 ;
      RECT 766.500000 347.590000 808.500000 348.410000 ;
      RECT 716.500000 347.590000 758.500000 348.410000 ;
      RECT 666.500000 347.590000 708.500000 348.410000 ;
      RECT 616.500000 347.590000 658.500000 348.410000 ;
      RECT 566.500000 347.590000 608.500000 348.410000 ;
      RECT 516.500000 347.590000 558.500000 348.410000 ;
      RECT 466.500000 347.590000 508.500000 348.410000 ;
      RECT 416.500000 347.590000 458.500000 349.590000 ;
      RECT 366.500000 347.590000 408.500000 348.410000 ;
      RECT 316.500000 347.590000 358.500000 348.410000 ;
      RECT 266.500000 347.590000 308.500000 348.410000 ;
      RECT 216.500000 347.590000 258.500000 348.410000 ;
      RECT 166.500000 347.590000 208.500000 348.410000 ;
      RECT 116.500000 347.590000 158.500000 348.410000 ;
      RECT 66.500000 347.590000 108.500000 348.410000 ;
      RECT 29.500000 347.590000 58.500000 349.590000 ;
      RECT 0.000000 347.590000 16.500000 348.410000 ;
      RECT 1169.500000 346.410000 1170.500000 347.590000 ;
      RECT 1116.500000 346.410000 1149.500000 347.590000 ;
      RECT 1107.500000 346.410000 1108.500000 347.590000 ;
      RECT 1066.500000 346.410000 1099.500000 347.590000 ;
      RECT 1057.500000 346.410000 1058.500000 347.590000 ;
      RECT 1016.500000 346.410000 1049.500000 347.590000 ;
      RECT 1007.500000 346.410000 1008.500000 347.590000 ;
      RECT 966.500000 346.410000 999.500000 347.590000 ;
      RECT 957.500000 346.410000 958.500000 347.590000 ;
      RECT 916.500000 346.410000 949.500000 347.590000 ;
      RECT 907.500000 346.410000 908.500000 347.590000 ;
      RECT 866.500000 346.410000 899.500000 347.590000 ;
      RECT 857.500000 346.410000 858.500000 347.590000 ;
      RECT 816.500000 346.410000 849.500000 347.590000 ;
      RECT 807.500000 346.410000 808.500000 347.590000 ;
      RECT 766.500000 346.410000 799.500000 347.590000 ;
      RECT 757.500000 346.410000 758.500000 347.590000 ;
      RECT 716.500000 346.410000 749.500000 347.590000 ;
      RECT 707.500000 346.410000 708.500000 347.590000 ;
      RECT 666.500000 346.410000 699.500000 347.590000 ;
      RECT 657.500000 346.410000 658.500000 347.590000 ;
      RECT 616.500000 346.410000 649.500000 347.590000 ;
      RECT 607.500000 346.410000 608.500000 347.590000 ;
      RECT 566.500000 346.410000 599.500000 347.590000 ;
      RECT 557.500000 346.410000 558.500000 347.590000 ;
      RECT 516.500000 346.410000 549.500000 347.590000 ;
      RECT 507.500000 346.410000 508.500000 347.590000 ;
      RECT 466.500000 346.410000 499.500000 347.590000 ;
      RECT 457.500000 346.410000 458.500000 347.590000 ;
      RECT 416.500000 346.410000 449.500000 347.590000 ;
      RECT 407.500000 346.410000 408.500000 347.590000 ;
      RECT 366.500000 346.410000 399.500000 347.590000 ;
      RECT 357.500000 346.410000 358.500000 347.590000 ;
      RECT 316.500000 346.410000 349.500000 347.590000 ;
      RECT 307.500000 346.410000 308.500000 347.590000 ;
      RECT 266.500000 346.410000 299.500000 347.590000 ;
      RECT 257.500000 346.410000 258.500000 347.590000 ;
      RECT 216.500000 346.410000 249.500000 347.590000 ;
      RECT 207.500000 346.410000 208.500000 347.590000 ;
      RECT 166.500000 346.410000 199.500000 347.590000 ;
      RECT 157.500000 346.410000 158.500000 347.590000 ;
      RECT 116.500000 346.410000 149.500000 347.590000 ;
      RECT 107.500000 346.410000 108.500000 347.590000 ;
      RECT 66.500000 346.410000 99.500000 347.590000 ;
      RECT 57.500000 346.410000 58.500000 347.590000 ;
      RECT 29.500000 346.410000 49.500000 347.590000 ;
      RECT 15.500000 346.410000 16.500000 347.590000 ;
      RECT 1157.500000 345.590000 1170.500000 346.410000 ;
      RECT 1107.500000 345.590000 1149.500000 346.410000 ;
      RECT 1057.500000 345.590000 1099.500000 346.410000 ;
      RECT 1007.500000 345.590000 1049.500000 346.410000 ;
      RECT 957.500000 345.590000 999.500000 346.410000 ;
      RECT 907.500000 345.590000 949.500000 346.410000 ;
      RECT 857.500000 345.590000 899.500000 346.410000 ;
      RECT 807.500000 345.590000 849.500000 346.410000 ;
      RECT 757.500000 345.590000 799.500000 346.410000 ;
      RECT 707.500000 345.590000 749.500000 346.410000 ;
      RECT 657.500000 345.590000 699.500000 346.410000 ;
      RECT 607.500000 345.590000 649.500000 346.410000 ;
      RECT 557.500000 345.590000 599.500000 346.410000 ;
      RECT 507.500000 345.590000 549.500000 346.410000 ;
      RECT 457.500000 345.590000 499.500000 346.410000 ;
      RECT 407.500000 345.590000 449.500000 346.410000 ;
      RECT 357.500000 345.590000 399.500000 346.410000 ;
      RECT 307.500000 345.590000 349.500000 346.410000 ;
      RECT 257.500000 345.590000 299.500000 346.410000 ;
      RECT 207.500000 345.590000 249.500000 346.410000 ;
      RECT 157.500000 345.590000 199.500000 346.410000 ;
      RECT 107.500000 345.590000 149.500000 346.410000 ;
      RECT 57.500000 345.590000 99.500000 346.410000 ;
      RECT 15.500000 345.590000 49.500000 346.410000 ;
      RECT 1183.500000 344.410000 1186.000000 347.590000 ;
      RECT 1169.500000 344.410000 1170.500000 345.590000 ;
      RECT 1116.500000 344.410000 1149.500000 345.590000 ;
      RECT 1107.500000 344.410000 1108.500000 345.590000 ;
      RECT 1066.500000 344.410000 1099.500000 345.590000 ;
      RECT 1057.500000 344.410000 1058.500000 345.590000 ;
      RECT 1016.500000 344.410000 1049.500000 345.590000 ;
      RECT 1007.500000 344.410000 1008.500000 345.590000 ;
      RECT 966.500000 344.410000 999.500000 345.590000 ;
      RECT 957.500000 344.410000 958.500000 345.590000 ;
      RECT 916.500000 344.410000 949.500000 345.590000 ;
      RECT 907.500000 344.410000 908.500000 345.590000 ;
      RECT 866.500000 344.410000 899.500000 345.590000 ;
      RECT 857.500000 344.410000 858.500000 345.590000 ;
      RECT 816.500000 344.410000 849.500000 345.590000 ;
      RECT 807.500000 344.410000 808.500000 345.590000 ;
      RECT 766.500000 344.410000 799.500000 345.590000 ;
      RECT 757.500000 344.410000 758.500000 345.590000 ;
      RECT 716.500000 344.410000 749.500000 345.590000 ;
      RECT 707.500000 344.410000 708.500000 345.590000 ;
      RECT 666.500000 344.410000 699.500000 345.590000 ;
      RECT 657.500000 344.410000 658.500000 345.590000 ;
      RECT 616.500000 344.410000 649.500000 345.590000 ;
      RECT 607.500000 344.410000 608.500000 345.590000 ;
      RECT 566.500000 344.410000 599.500000 345.590000 ;
      RECT 557.500000 344.410000 558.500000 345.590000 ;
      RECT 516.500000 344.410000 549.500000 345.590000 ;
      RECT 507.500000 344.410000 508.500000 345.590000 ;
      RECT 466.500000 344.410000 499.500000 345.590000 ;
      RECT 457.500000 344.410000 458.500000 345.590000 ;
      RECT 416.500000 344.410000 449.500000 345.590000 ;
      RECT 407.500000 344.410000 408.500000 345.590000 ;
      RECT 366.500000 344.410000 399.500000 345.590000 ;
      RECT 357.500000 344.410000 358.500000 345.590000 ;
      RECT 316.500000 344.410000 349.500000 345.590000 ;
      RECT 307.500000 344.410000 308.500000 345.590000 ;
      RECT 266.500000 344.410000 299.500000 345.590000 ;
      RECT 257.500000 344.410000 258.500000 345.590000 ;
      RECT 216.500000 344.410000 249.500000 345.590000 ;
      RECT 207.500000 344.410000 208.500000 345.590000 ;
      RECT 166.500000 344.410000 199.500000 345.590000 ;
      RECT 157.500000 344.410000 158.500000 345.590000 ;
      RECT 116.500000 344.410000 149.500000 345.590000 ;
      RECT 107.500000 344.410000 108.500000 345.590000 ;
      RECT 66.500000 344.410000 99.500000 345.590000 ;
      RECT 57.500000 344.410000 58.500000 345.590000 ;
      RECT 29.500000 344.410000 49.500000 345.590000 ;
      RECT 15.500000 344.410000 16.500000 345.590000 ;
      RECT 0.000000 344.410000 2.500000 347.590000 ;
      RECT 1169.500000 343.590000 1186.000000 344.410000 ;
      RECT 1116.500000 343.590000 1156.500000 344.410000 ;
      RECT 1066.500000 343.590000 1108.500000 344.410000 ;
      RECT 1016.500000 343.590000 1058.500000 344.410000 ;
      RECT 966.500000 343.590000 1008.500000 344.410000 ;
      RECT 916.500000 343.590000 958.500000 344.410000 ;
      RECT 866.500000 343.590000 908.500000 344.410000 ;
      RECT 816.500000 343.590000 858.500000 344.410000 ;
      RECT 766.500000 343.590000 808.500000 344.410000 ;
      RECT 716.500000 343.590000 758.500000 344.410000 ;
      RECT 666.500000 343.590000 708.500000 344.410000 ;
      RECT 616.500000 343.590000 658.500000 344.410000 ;
      RECT 566.500000 343.590000 608.500000 344.410000 ;
      RECT 516.500000 343.590000 558.500000 344.410000 ;
      RECT 466.500000 343.590000 508.500000 344.410000 ;
      RECT 416.500000 343.590000 458.500000 344.410000 ;
      RECT 366.500000 343.590000 408.500000 344.410000 ;
      RECT 316.500000 343.590000 358.500000 344.410000 ;
      RECT 266.500000 343.590000 308.500000 344.410000 ;
      RECT 216.500000 343.590000 258.500000 344.410000 ;
      RECT 166.500000 343.590000 208.500000 344.410000 ;
      RECT 116.500000 343.590000 158.500000 344.410000 ;
      RECT 66.500000 343.590000 108.500000 344.410000 ;
      RECT 29.500000 343.590000 58.500000 344.410000 ;
      RECT 0.000000 343.590000 16.500000 344.410000 ;
      RECT 1169.500000 342.410000 1170.500000 343.590000 ;
      RECT 1116.500000 342.410000 1149.500000 343.590000 ;
      RECT 1107.500000 342.410000 1108.500000 343.590000 ;
      RECT 1066.500000 342.410000 1099.500000 343.590000 ;
      RECT 1057.500000 342.410000 1058.500000 343.590000 ;
      RECT 1016.500000 342.410000 1049.500000 343.590000 ;
      RECT 1007.500000 342.410000 1008.500000 343.590000 ;
      RECT 966.500000 342.410000 999.500000 343.590000 ;
      RECT 957.500000 342.410000 958.500000 343.590000 ;
      RECT 916.500000 342.410000 949.500000 343.590000 ;
      RECT 907.500000 342.410000 908.500000 343.590000 ;
      RECT 866.500000 342.410000 899.500000 343.590000 ;
      RECT 857.500000 342.410000 858.500000 343.590000 ;
      RECT 816.500000 342.410000 849.500000 343.590000 ;
      RECT 807.500000 342.410000 808.500000 343.590000 ;
      RECT 766.500000 342.410000 799.500000 343.590000 ;
      RECT 757.500000 342.410000 758.500000 343.590000 ;
      RECT 716.500000 342.410000 749.500000 343.590000 ;
      RECT 707.500000 342.410000 708.500000 343.590000 ;
      RECT 666.500000 342.410000 699.500000 343.590000 ;
      RECT 657.500000 342.410000 658.500000 343.590000 ;
      RECT 616.500000 342.410000 649.500000 343.590000 ;
      RECT 607.500000 342.410000 608.500000 343.590000 ;
      RECT 566.500000 342.410000 599.500000 343.590000 ;
      RECT 557.500000 342.410000 558.500000 343.590000 ;
      RECT 516.500000 342.410000 549.500000 343.590000 ;
      RECT 507.500000 342.410000 508.500000 343.590000 ;
      RECT 466.500000 342.410000 499.500000 343.590000 ;
      RECT 457.500000 342.410000 458.500000 343.590000 ;
      RECT 416.500000 342.410000 449.500000 343.590000 ;
      RECT 407.500000 342.410000 408.500000 343.590000 ;
      RECT 366.500000 342.410000 399.500000 343.590000 ;
      RECT 357.500000 342.410000 358.500000 343.590000 ;
      RECT 316.500000 342.410000 349.500000 343.590000 ;
      RECT 307.500000 342.410000 308.500000 343.590000 ;
      RECT 266.500000 342.410000 299.500000 343.590000 ;
      RECT 257.500000 342.410000 258.500000 343.590000 ;
      RECT 216.500000 342.410000 249.500000 343.590000 ;
      RECT 207.500000 342.410000 208.500000 343.590000 ;
      RECT 166.500000 342.410000 199.500000 343.590000 ;
      RECT 157.500000 342.410000 158.500000 343.590000 ;
      RECT 116.500000 342.410000 149.500000 343.590000 ;
      RECT 107.500000 342.410000 108.500000 343.590000 ;
      RECT 66.500000 342.410000 99.500000 343.590000 ;
      RECT 57.500000 342.410000 58.500000 343.590000 ;
      RECT 29.500000 342.410000 49.500000 343.590000 ;
      RECT 15.500000 342.410000 16.500000 343.590000 ;
      RECT 1157.500000 341.590000 1170.500000 342.410000 ;
      RECT 1107.500000 341.590000 1149.500000 342.410000 ;
      RECT 1057.500000 341.590000 1099.500000 342.410000 ;
      RECT 1007.500000 341.590000 1049.500000 342.410000 ;
      RECT 957.500000 341.590000 999.500000 342.410000 ;
      RECT 907.500000 341.590000 949.500000 342.410000 ;
      RECT 857.500000 341.590000 899.500000 342.410000 ;
      RECT 807.500000 341.590000 849.500000 342.410000 ;
      RECT 757.500000 341.590000 799.500000 342.410000 ;
      RECT 707.500000 341.590000 749.500000 342.410000 ;
      RECT 657.500000 341.590000 699.500000 342.410000 ;
      RECT 607.500000 341.590000 649.500000 342.410000 ;
      RECT 557.500000 341.590000 599.500000 342.410000 ;
      RECT 507.500000 341.590000 549.500000 342.410000 ;
      RECT 457.500000 341.590000 499.500000 342.410000 ;
      RECT 407.500000 341.590000 449.500000 342.410000 ;
      RECT 357.500000 341.590000 399.500000 342.410000 ;
      RECT 307.500000 341.590000 349.500000 342.410000 ;
      RECT 257.500000 341.590000 299.500000 342.410000 ;
      RECT 207.500000 341.590000 249.500000 342.410000 ;
      RECT 157.500000 341.590000 199.500000 342.410000 ;
      RECT 107.500000 341.590000 149.500000 342.410000 ;
      RECT 57.500000 341.590000 99.500000 342.410000 ;
      RECT 15.500000 341.590000 49.500000 342.410000 ;
      RECT 1183.500000 340.410000 1186.000000 343.590000 ;
      RECT 1169.500000 340.410000 1170.500000 341.590000 ;
      RECT 1116.500000 340.410000 1149.500000 341.590000 ;
      RECT 1107.500000 340.410000 1108.500000 341.590000 ;
      RECT 1066.500000 340.410000 1099.500000 341.590000 ;
      RECT 1057.500000 340.410000 1058.500000 341.590000 ;
      RECT 1016.500000 340.410000 1049.500000 341.590000 ;
      RECT 1007.500000 340.410000 1008.500000 341.590000 ;
      RECT 966.500000 340.410000 999.500000 341.590000 ;
      RECT 957.500000 340.410000 958.500000 341.590000 ;
      RECT 916.500000 340.410000 949.500000 341.590000 ;
      RECT 907.500000 340.410000 908.500000 341.590000 ;
      RECT 866.500000 340.410000 899.500000 341.590000 ;
      RECT 857.500000 340.410000 858.500000 341.590000 ;
      RECT 816.500000 340.410000 849.500000 341.590000 ;
      RECT 807.500000 340.410000 808.500000 341.590000 ;
      RECT 766.500000 340.410000 799.500000 341.590000 ;
      RECT 757.500000 340.410000 758.500000 341.590000 ;
      RECT 716.500000 340.410000 749.500000 341.590000 ;
      RECT 707.500000 340.410000 708.500000 341.590000 ;
      RECT 666.500000 340.410000 699.500000 341.590000 ;
      RECT 657.500000 340.410000 658.500000 341.590000 ;
      RECT 616.500000 340.410000 649.500000 341.590000 ;
      RECT 607.500000 340.410000 608.500000 341.590000 ;
      RECT 566.500000 340.410000 599.500000 341.590000 ;
      RECT 557.500000 340.410000 558.500000 341.590000 ;
      RECT 516.500000 340.410000 549.500000 341.590000 ;
      RECT 507.500000 340.410000 508.500000 341.590000 ;
      RECT 466.500000 340.410000 499.500000 341.590000 ;
      RECT 457.500000 340.410000 458.500000 341.590000 ;
      RECT 416.500000 340.410000 449.500000 341.590000 ;
      RECT 407.500000 340.410000 408.500000 341.590000 ;
      RECT 366.500000 340.410000 399.500000 341.590000 ;
      RECT 357.500000 340.410000 358.500000 341.590000 ;
      RECT 316.500000 340.410000 349.500000 341.590000 ;
      RECT 307.500000 340.410000 308.500000 341.590000 ;
      RECT 266.500000 340.410000 299.500000 341.590000 ;
      RECT 257.500000 340.410000 258.500000 341.590000 ;
      RECT 216.500000 340.410000 249.500000 341.590000 ;
      RECT 207.500000 340.410000 208.500000 341.590000 ;
      RECT 166.500000 340.410000 199.500000 341.590000 ;
      RECT 157.500000 340.410000 158.500000 341.590000 ;
      RECT 116.500000 340.410000 149.500000 341.590000 ;
      RECT 107.500000 340.410000 108.500000 341.590000 ;
      RECT 66.500000 340.410000 99.500000 341.590000 ;
      RECT 57.500000 340.410000 58.500000 341.590000 ;
      RECT 29.500000 340.410000 49.500000 341.590000 ;
      RECT 15.500000 340.410000 16.500000 341.590000 ;
      RECT 0.000000 340.410000 2.500000 343.590000 ;
      RECT 1169.500000 339.590000 1186.000000 340.410000 ;
      RECT 1116.500000 339.590000 1156.500000 340.410000 ;
      RECT 1066.500000 339.590000 1108.500000 340.410000 ;
      RECT 1016.500000 339.590000 1058.500000 340.410000 ;
      RECT 966.500000 339.590000 1008.500000 340.410000 ;
      RECT 916.500000 339.590000 958.500000 340.410000 ;
      RECT 866.500000 339.590000 908.500000 340.410000 ;
      RECT 816.500000 339.590000 858.500000 340.410000 ;
      RECT 766.500000 339.590000 808.500000 340.410000 ;
      RECT 716.500000 339.590000 758.500000 340.410000 ;
      RECT 666.500000 339.590000 708.500000 340.410000 ;
      RECT 616.500000 339.590000 658.500000 340.410000 ;
      RECT 566.500000 339.590000 608.500000 340.410000 ;
      RECT 516.500000 339.590000 558.500000 340.410000 ;
      RECT 466.500000 339.590000 508.500000 340.410000 ;
      RECT 416.500000 339.590000 458.500000 340.410000 ;
      RECT 366.500000 339.590000 408.500000 340.410000 ;
      RECT 316.500000 339.590000 358.500000 340.410000 ;
      RECT 266.500000 339.590000 308.500000 340.410000 ;
      RECT 216.500000 339.590000 258.500000 340.410000 ;
      RECT 166.500000 339.590000 208.500000 340.410000 ;
      RECT 116.500000 339.590000 158.500000 340.410000 ;
      RECT 66.500000 339.590000 108.500000 340.410000 ;
      RECT 29.500000 339.590000 58.500000 340.410000 ;
      RECT 0.000000 339.590000 16.500000 340.410000 ;
      RECT 1169.500000 338.410000 1170.500000 339.590000 ;
      RECT 1116.500000 338.410000 1149.500000 339.590000 ;
      RECT 1107.500000 338.410000 1108.500000 339.590000 ;
      RECT 1066.500000 338.410000 1099.500000 339.590000 ;
      RECT 1057.500000 338.410000 1058.500000 339.590000 ;
      RECT 1016.500000 338.410000 1049.500000 339.590000 ;
      RECT 1007.500000 338.410000 1008.500000 339.590000 ;
      RECT 966.500000 338.410000 999.500000 339.590000 ;
      RECT 957.500000 338.410000 958.500000 339.590000 ;
      RECT 916.500000 338.410000 949.500000 339.590000 ;
      RECT 907.500000 338.410000 908.500000 339.590000 ;
      RECT 866.500000 338.410000 899.500000 339.590000 ;
      RECT 857.500000 338.410000 858.500000 339.590000 ;
      RECT 816.500000 338.410000 849.500000 339.590000 ;
      RECT 807.500000 338.410000 808.500000 339.590000 ;
      RECT 766.500000 338.410000 799.500000 339.590000 ;
      RECT 757.500000 338.410000 758.500000 339.590000 ;
      RECT 716.500000 338.410000 749.500000 339.590000 ;
      RECT 707.500000 338.410000 708.500000 339.590000 ;
      RECT 666.500000 338.410000 699.500000 339.590000 ;
      RECT 657.500000 338.410000 658.500000 339.590000 ;
      RECT 616.500000 338.410000 649.500000 339.590000 ;
      RECT 607.500000 338.410000 608.500000 339.590000 ;
      RECT 566.500000 338.410000 599.500000 339.590000 ;
      RECT 557.500000 338.410000 558.500000 339.590000 ;
      RECT 516.500000 338.410000 549.500000 339.590000 ;
      RECT 507.500000 338.410000 508.500000 339.590000 ;
      RECT 466.500000 338.410000 499.500000 339.590000 ;
      RECT 457.500000 338.410000 458.500000 339.590000 ;
      RECT 416.500000 338.410000 449.500000 339.590000 ;
      RECT 407.500000 338.410000 408.500000 339.590000 ;
      RECT 366.500000 338.410000 399.500000 339.590000 ;
      RECT 357.500000 338.410000 358.500000 339.590000 ;
      RECT 316.500000 338.410000 349.500000 339.590000 ;
      RECT 307.500000 338.410000 308.500000 339.590000 ;
      RECT 266.500000 338.410000 299.500000 339.590000 ;
      RECT 257.500000 338.410000 258.500000 339.590000 ;
      RECT 216.500000 338.410000 249.500000 339.590000 ;
      RECT 207.500000 338.410000 208.500000 339.590000 ;
      RECT 166.500000 338.410000 199.500000 339.590000 ;
      RECT 157.500000 338.410000 158.500000 339.590000 ;
      RECT 116.500000 338.410000 149.500000 339.590000 ;
      RECT 107.500000 338.410000 108.500000 339.590000 ;
      RECT 66.500000 338.410000 99.500000 339.590000 ;
      RECT 57.500000 338.410000 58.500000 339.590000 ;
      RECT 29.500000 338.410000 49.500000 339.590000 ;
      RECT 15.500000 338.410000 16.500000 339.590000 ;
      RECT 1157.500000 337.590000 1170.500000 338.410000 ;
      RECT 1107.500000 337.590000 1149.500000 338.410000 ;
      RECT 1057.500000 337.590000 1099.500000 338.410000 ;
      RECT 1007.500000 337.590000 1049.500000 338.410000 ;
      RECT 957.500000 337.590000 999.500000 338.410000 ;
      RECT 907.500000 337.590000 949.500000 338.410000 ;
      RECT 857.500000 337.590000 899.500000 338.410000 ;
      RECT 807.500000 337.590000 849.500000 338.410000 ;
      RECT 757.500000 337.590000 799.500000 338.410000 ;
      RECT 707.500000 337.590000 749.500000 338.410000 ;
      RECT 657.500000 337.590000 699.500000 338.410000 ;
      RECT 607.500000 337.590000 649.500000 338.410000 ;
      RECT 557.500000 337.590000 599.500000 338.410000 ;
      RECT 507.500000 337.590000 549.500000 338.410000 ;
      RECT 457.500000 337.590000 499.500000 338.410000 ;
      RECT 407.500000 337.590000 449.500000 338.410000 ;
      RECT 357.500000 337.590000 399.500000 338.410000 ;
      RECT 307.500000 337.590000 349.500000 338.410000 ;
      RECT 257.500000 337.590000 299.500000 338.410000 ;
      RECT 207.500000 337.590000 249.500000 338.410000 ;
      RECT 157.500000 337.590000 199.500000 338.410000 ;
      RECT 107.500000 337.590000 149.500000 338.410000 ;
      RECT 57.500000 337.590000 99.500000 338.410000 ;
      RECT 15.500000 337.590000 49.500000 338.410000 ;
      RECT 1183.500000 336.410000 1186.000000 339.590000 ;
      RECT 1169.500000 336.410000 1170.500000 337.590000 ;
      RECT 1116.500000 336.410000 1149.500000 337.590000 ;
      RECT 1107.500000 336.410000 1108.500000 337.590000 ;
      RECT 1066.500000 336.410000 1099.500000 337.590000 ;
      RECT 1057.500000 336.410000 1058.500000 337.590000 ;
      RECT 1016.500000 336.410000 1049.500000 337.590000 ;
      RECT 1007.500000 336.410000 1008.500000 337.590000 ;
      RECT 966.500000 336.410000 999.500000 337.590000 ;
      RECT 957.500000 336.410000 958.500000 337.590000 ;
      RECT 916.500000 336.410000 949.500000 337.590000 ;
      RECT 907.500000 336.410000 908.500000 337.590000 ;
      RECT 866.500000 336.410000 899.500000 337.590000 ;
      RECT 857.500000 336.410000 858.500000 337.590000 ;
      RECT 816.500000 336.410000 849.500000 337.590000 ;
      RECT 807.500000 336.410000 808.500000 337.590000 ;
      RECT 766.500000 336.410000 799.500000 337.590000 ;
      RECT 757.500000 336.410000 758.500000 337.590000 ;
      RECT 716.500000 336.410000 749.500000 337.590000 ;
      RECT 707.500000 336.410000 708.500000 337.590000 ;
      RECT 666.500000 336.410000 699.500000 337.590000 ;
      RECT 657.500000 336.410000 658.500000 337.590000 ;
      RECT 616.500000 336.410000 649.500000 337.590000 ;
      RECT 607.500000 336.410000 608.500000 337.590000 ;
      RECT 566.500000 336.410000 599.500000 337.590000 ;
      RECT 557.500000 336.410000 558.500000 337.590000 ;
      RECT 516.500000 336.410000 549.500000 337.590000 ;
      RECT 507.500000 336.410000 508.500000 337.590000 ;
      RECT 466.500000 336.410000 499.500000 337.590000 ;
      RECT 457.500000 336.410000 458.500000 337.590000 ;
      RECT 416.500000 336.410000 449.500000 337.590000 ;
      RECT 407.500000 336.410000 408.500000 337.590000 ;
      RECT 366.500000 336.410000 399.500000 337.590000 ;
      RECT 357.500000 336.410000 358.500000 337.590000 ;
      RECT 316.500000 336.410000 349.500000 337.590000 ;
      RECT 307.500000 336.410000 308.500000 337.590000 ;
      RECT 266.500000 336.410000 299.500000 337.590000 ;
      RECT 257.500000 336.410000 258.500000 337.590000 ;
      RECT 216.500000 336.410000 249.500000 337.590000 ;
      RECT 207.500000 336.410000 208.500000 337.590000 ;
      RECT 166.500000 336.410000 199.500000 337.590000 ;
      RECT 157.500000 336.410000 158.500000 337.590000 ;
      RECT 116.500000 336.410000 149.500000 337.590000 ;
      RECT 107.500000 336.410000 108.500000 337.590000 ;
      RECT 66.500000 336.410000 99.500000 337.590000 ;
      RECT 57.500000 336.410000 58.500000 337.590000 ;
      RECT 29.500000 336.410000 49.500000 337.590000 ;
      RECT 15.500000 336.410000 16.500000 337.590000 ;
      RECT 0.000000 336.410000 2.500000 339.590000 ;
      RECT 1169.500000 335.590000 1186.000000 336.410000 ;
      RECT 1116.500000 335.590000 1156.500000 336.410000 ;
      RECT 1066.500000 335.590000 1108.500000 336.410000 ;
      RECT 1016.500000 335.590000 1058.500000 336.410000 ;
      RECT 966.500000 335.590000 1008.500000 336.410000 ;
      RECT 916.500000 335.590000 958.500000 336.410000 ;
      RECT 866.500000 335.590000 908.500000 336.410000 ;
      RECT 816.500000 335.590000 858.500000 336.410000 ;
      RECT 766.500000 335.590000 808.500000 336.410000 ;
      RECT 716.500000 335.590000 758.500000 336.410000 ;
      RECT 666.500000 335.590000 708.500000 336.410000 ;
      RECT 616.500000 335.590000 658.500000 336.410000 ;
      RECT 566.500000 335.590000 608.500000 336.410000 ;
      RECT 516.500000 335.590000 558.500000 336.410000 ;
      RECT 466.500000 335.590000 508.500000 336.410000 ;
      RECT 416.500000 335.590000 458.500000 336.410000 ;
      RECT 366.500000 335.590000 408.500000 336.410000 ;
      RECT 316.500000 335.590000 358.500000 336.410000 ;
      RECT 266.500000 335.590000 308.500000 336.410000 ;
      RECT 216.500000 335.590000 258.500000 336.410000 ;
      RECT 166.500000 335.590000 208.500000 336.410000 ;
      RECT 116.500000 335.590000 158.500000 336.410000 ;
      RECT 66.500000 335.590000 108.500000 336.410000 ;
      RECT 29.500000 335.590000 58.500000 336.410000 ;
      RECT 0.000000 335.590000 16.500000 336.410000 ;
      RECT 1169.500000 334.410000 1170.500000 335.590000 ;
      RECT 1116.500000 334.410000 1149.500000 335.590000 ;
      RECT 1107.500000 334.410000 1108.500000 335.590000 ;
      RECT 1066.500000 334.410000 1099.500000 335.590000 ;
      RECT 1057.500000 334.410000 1058.500000 335.590000 ;
      RECT 1016.500000 334.410000 1049.500000 335.590000 ;
      RECT 1007.500000 334.410000 1008.500000 335.590000 ;
      RECT 966.500000 334.410000 999.500000 335.590000 ;
      RECT 957.500000 334.410000 958.500000 335.590000 ;
      RECT 916.500000 334.410000 949.500000 335.590000 ;
      RECT 907.500000 334.410000 908.500000 335.590000 ;
      RECT 866.500000 334.410000 899.500000 335.590000 ;
      RECT 857.500000 334.410000 858.500000 335.590000 ;
      RECT 816.500000 334.410000 849.500000 335.590000 ;
      RECT 807.500000 334.410000 808.500000 335.590000 ;
      RECT 766.500000 334.410000 799.500000 335.590000 ;
      RECT 757.500000 334.410000 758.500000 335.590000 ;
      RECT 716.500000 334.410000 749.500000 335.590000 ;
      RECT 707.500000 334.410000 708.500000 335.590000 ;
      RECT 666.500000 334.410000 699.500000 335.590000 ;
      RECT 657.500000 334.410000 658.500000 335.590000 ;
      RECT 616.500000 334.410000 649.500000 335.590000 ;
      RECT 607.500000 334.410000 608.500000 335.590000 ;
      RECT 566.500000 334.410000 599.500000 335.590000 ;
      RECT 557.500000 334.410000 558.500000 335.590000 ;
      RECT 516.500000 334.410000 549.500000 335.590000 ;
      RECT 507.500000 334.410000 508.500000 335.590000 ;
      RECT 466.500000 334.410000 499.500000 335.590000 ;
      RECT 457.500000 334.410000 458.500000 335.590000 ;
      RECT 416.500000 334.410000 449.500000 335.590000 ;
      RECT 407.500000 334.410000 408.500000 335.590000 ;
      RECT 366.500000 334.410000 399.500000 335.590000 ;
      RECT 357.500000 334.410000 358.500000 335.590000 ;
      RECT 316.500000 334.410000 349.500000 335.590000 ;
      RECT 307.500000 334.410000 308.500000 335.590000 ;
      RECT 266.500000 334.410000 299.500000 335.590000 ;
      RECT 257.500000 334.410000 258.500000 335.590000 ;
      RECT 216.500000 334.410000 249.500000 335.590000 ;
      RECT 207.500000 334.410000 208.500000 335.590000 ;
      RECT 166.500000 334.410000 199.500000 335.590000 ;
      RECT 157.500000 334.410000 158.500000 335.590000 ;
      RECT 116.500000 334.410000 149.500000 335.590000 ;
      RECT 107.500000 334.410000 108.500000 335.590000 ;
      RECT 66.500000 334.410000 99.500000 335.590000 ;
      RECT 57.500000 334.410000 58.500000 335.590000 ;
      RECT 29.500000 334.410000 49.500000 335.590000 ;
      RECT 15.500000 334.410000 16.500000 335.590000 ;
      RECT 1157.500000 333.590000 1170.500000 334.410000 ;
      RECT 1107.500000 333.590000 1149.500000 334.410000 ;
      RECT 1057.500000 333.590000 1099.500000 334.410000 ;
      RECT 1007.500000 333.590000 1049.500000 334.410000 ;
      RECT 957.500000 333.590000 999.500000 334.410000 ;
      RECT 907.500000 333.590000 949.500000 334.410000 ;
      RECT 857.500000 333.590000 899.500000 334.410000 ;
      RECT 807.500000 333.590000 849.500000 334.410000 ;
      RECT 757.500000 333.590000 799.500000 334.410000 ;
      RECT 707.500000 333.590000 749.500000 334.410000 ;
      RECT 657.500000 333.590000 699.500000 334.410000 ;
      RECT 607.500000 333.590000 649.500000 334.410000 ;
      RECT 557.500000 333.590000 599.500000 334.410000 ;
      RECT 507.500000 333.590000 549.500000 334.410000 ;
      RECT 457.500000 333.590000 499.500000 334.410000 ;
      RECT 407.500000 333.590000 449.500000 334.410000 ;
      RECT 357.500000 333.590000 399.500000 334.410000 ;
      RECT 307.500000 333.590000 349.500000 334.410000 ;
      RECT 257.500000 333.590000 299.500000 334.410000 ;
      RECT 207.500000 333.590000 249.500000 334.410000 ;
      RECT 157.500000 333.590000 199.500000 334.410000 ;
      RECT 107.500000 333.590000 149.500000 334.410000 ;
      RECT 57.500000 333.590000 99.500000 334.410000 ;
      RECT 15.500000 333.590000 49.500000 334.410000 ;
      RECT 1183.500000 332.410000 1186.000000 335.590000 ;
      RECT 1169.500000 332.410000 1170.500000 333.590000 ;
      RECT 1116.500000 332.410000 1149.500000 333.590000 ;
      RECT 1107.500000 332.410000 1108.500000 333.590000 ;
      RECT 1066.500000 332.410000 1099.500000 333.590000 ;
      RECT 1057.500000 332.410000 1058.500000 333.590000 ;
      RECT 1016.500000 332.410000 1049.500000 333.590000 ;
      RECT 1007.500000 332.410000 1008.500000 333.590000 ;
      RECT 966.500000 332.410000 999.500000 333.590000 ;
      RECT 957.500000 332.410000 958.500000 333.590000 ;
      RECT 916.500000 332.410000 949.500000 333.590000 ;
      RECT 907.500000 332.410000 908.500000 333.590000 ;
      RECT 866.500000 332.410000 899.500000 333.590000 ;
      RECT 857.500000 332.410000 858.500000 333.590000 ;
      RECT 816.500000 332.410000 849.500000 333.590000 ;
      RECT 807.500000 332.410000 808.500000 333.590000 ;
      RECT 766.500000 332.410000 799.500000 333.590000 ;
      RECT 757.500000 332.410000 758.500000 333.590000 ;
      RECT 716.500000 332.410000 749.500000 333.590000 ;
      RECT 707.500000 332.410000 708.500000 333.590000 ;
      RECT 666.500000 332.410000 699.500000 333.590000 ;
      RECT 657.500000 332.410000 658.500000 333.590000 ;
      RECT 616.500000 332.410000 649.500000 333.590000 ;
      RECT 607.500000 332.410000 608.500000 333.590000 ;
      RECT 566.500000 332.410000 599.500000 333.590000 ;
      RECT 557.500000 332.410000 558.500000 333.590000 ;
      RECT 516.500000 332.410000 549.500000 333.590000 ;
      RECT 507.500000 332.410000 508.500000 333.590000 ;
      RECT 466.500000 332.410000 499.500000 333.590000 ;
      RECT 457.500000 332.410000 458.500000 333.590000 ;
      RECT 416.500000 332.410000 449.500000 333.590000 ;
      RECT 407.500000 332.410000 408.500000 333.590000 ;
      RECT 366.500000 332.410000 399.500000 333.590000 ;
      RECT 357.500000 332.410000 358.500000 333.590000 ;
      RECT 316.500000 332.410000 349.500000 333.590000 ;
      RECT 307.500000 332.410000 308.500000 333.590000 ;
      RECT 266.500000 332.410000 299.500000 333.590000 ;
      RECT 257.500000 332.410000 258.500000 333.590000 ;
      RECT 216.500000 332.410000 249.500000 333.590000 ;
      RECT 207.500000 332.410000 208.500000 333.590000 ;
      RECT 166.500000 332.410000 199.500000 333.590000 ;
      RECT 157.500000 332.410000 158.500000 333.590000 ;
      RECT 116.500000 332.410000 149.500000 333.590000 ;
      RECT 107.500000 332.410000 108.500000 333.590000 ;
      RECT 66.500000 332.410000 99.500000 333.590000 ;
      RECT 57.500000 332.410000 58.500000 333.590000 ;
      RECT 29.500000 332.410000 49.500000 333.590000 ;
      RECT 15.500000 332.410000 16.500000 333.590000 ;
      RECT 0.000000 332.410000 2.500000 335.590000 ;
      RECT 1169.500000 331.590000 1186.000000 332.410000 ;
      RECT 1116.500000 331.590000 1156.500000 332.410000 ;
      RECT 1066.500000 331.590000 1108.500000 332.410000 ;
      RECT 1016.500000 331.590000 1058.500000 332.410000 ;
      RECT 966.500000 331.590000 1008.500000 332.410000 ;
      RECT 916.500000 331.590000 958.500000 332.410000 ;
      RECT 866.500000 331.590000 908.500000 332.410000 ;
      RECT 816.500000 331.590000 858.500000 332.410000 ;
      RECT 766.500000 331.590000 808.500000 332.410000 ;
      RECT 716.500000 331.590000 758.500000 332.410000 ;
      RECT 666.500000 331.590000 708.500000 332.410000 ;
      RECT 616.500000 331.590000 658.500000 332.410000 ;
      RECT 566.500000 331.590000 608.500000 332.410000 ;
      RECT 516.500000 331.590000 558.500000 332.410000 ;
      RECT 466.500000 331.590000 508.500000 332.410000 ;
      RECT 416.500000 331.590000 458.500000 332.410000 ;
      RECT 366.500000 331.590000 408.500000 332.410000 ;
      RECT 316.500000 331.590000 358.500000 332.410000 ;
      RECT 266.500000 331.590000 308.500000 332.410000 ;
      RECT 216.500000 331.590000 258.500000 332.410000 ;
      RECT 166.500000 331.590000 208.500000 332.410000 ;
      RECT 116.500000 331.590000 158.500000 332.410000 ;
      RECT 66.500000 331.590000 108.500000 332.410000 ;
      RECT 29.500000 331.590000 58.500000 332.410000 ;
      RECT 0.000000 331.590000 16.500000 332.410000 ;
      RECT 1169.500000 330.410000 1170.500000 331.590000 ;
      RECT 1116.500000 330.410000 1149.500000 331.590000 ;
      RECT 1107.500000 330.410000 1108.500000 331.590000 ;
      RECT 1066.500000 330.410000 1099.500000 331.590000 ;
      RECT 1057.500000 330.410000 1058.500000 331.590000 ;
      RECT 1016.500000 330.410000 1049.500000 331.590000 ;
      RECT 1007.500000 330.410000 1008.500000 331.590000 ;
      RECT 966.500000 330.410000 999.500000 331.590000 ;
      RECT 957.500000 330.410000 958.500000 331.590000 ;
      RECT 916.500000 330.410000 949.500000 331.590000 ;
      RECT 907.500000 330.410000 908.500000 331.590000 ;
      RECT 866.500000 330.410000 899.500000 331.590000 ;
      RECT 857.500000 330.410000 858.500000 331.590000 ;
      RECT 816.500000 330.410000 849.500000 331.590000 ;
      RECT 807.500000 330.410000 808.500000 331.590000 ;
      RECT 766.500000 330.410000 799.500000 331.590000 ;
      RECT 757.500000 330.410000 758.500000 331.590000 ;
      RECT 716.500000 330.410000 749.500000 331.590000 ;
      RECT 707.500000 330.410000 708.500000 331.590000 ;
      RECT 666.500000 330.410000 699.500000 331.590000 ;
      RECT 657.500000 330.410000 658.500000 331.590000 ;
      RECT 616.500000 330.410000 649.500000 331.590000 ;
      RECT 607.500000 330.410000 608.500000 331.590000 ;
      RECT 566.500000 330.410000 599.500000 331.590000 ;
      RECT 557.500000 330.410000 558.500000 331.590000 ;
      RECT 516.500000 330.410000 549.500000 331.590000 ;
      RECT 507.500000 330.410000 508.500000 331.590000 ;
      RECT 466.500000 330.410000 499.500000 331.590000 ;
      RECT 457.500000 330.410000 458.500000 331.590000 ;
      RECT 416.500000 330.410000 449.500000 331.590000 ;
      RECT 407.500000 330.410000 408.500000 331.590000 ;
      RECT 366.500000 330.410000 399.500000 331.590000 ;
      RECT 357.500000 330.410000 358.500000 331.590000 ;
      RECT 316.500000 330.410000 349.500000 331.590000 ;
      RECT 307.500000 330.410000 308.500000 331.590000 ;
      RECT 266.500000 330.410000 299.500000 331.590000 ;
      RECT 257.500000 330.410000 258.500000 331.590000 ;
      RECT 216.500000 330.410000 249.500000 331.590000 ;
      RECT 207.500000 330.410000 208.500000 331.590000 ;
      RECT 166.500000 330.410000 199.500000 331.590000 ;
      RECT 157.500000 330.410000 158.500000 331.590000 ;
      RECT 116.500000 330.410000 149.500000 331.590000 ;
      RECT 107.500000 330.410000 108.500000 331.590000 ;
      RECT 66.500000 330.410000 99.500000 331.590000 ;
      RECT 57.500000 330.410000 58.500000 331.590000 ;
      RECT 29.500000 330.410000 49.500000 331.590000 ;
      RECT 15.500000 330.410000 16.500000 331.590000 ;
      RECT 1157.500000 329.590000 1170.500000 330.410000 ;
      RECT 1107.500000 329.590000 1149.500000 330.410000 ;
      RECT 1057.500000 329.590000 1099.500000 330.410000 ;
      RECT 1007.500000 329.590000 1049.500000 330.410000 ;
      RECT 957.500000 329.590000 999.500000 330.410000 ;
      RECT 907.500000 329.590000 949.500000 330.410000 ;
      RECT 857.500000 329.590000 899.500000 330.410000 ;
      RECT 807.500000 329.590000 849.500000 330.410000 ;
      RECT 757.500000 329.590000 799.500000 330.410000 ;
      RECT 707.500000 329.590000 749.500000 330.410000 ;
      RECT 657.500000 329.590000 699.500000 330.410000 ;
      RECT 607.500000 329.590000 649.500000 330.410000 ;
      RECT 557.500000 329.590000 599.500000 330.410000 ;
      RECT 507.500000 329.590000 549.500000 330.410000 ;
      RECT 457.500000 329.590000 499.500000 330.410000 ;
      RECT 407.500000 329.590000 449.500000 330.410000 ;
      RECT 357.500000 329.590000 399.500000 330.410000 ;
      RECT 307.500000 329.590000 349.500000 330.410000 ;
      RECT 257.500000 329.590000 299.500000 330.410000 ;
      RECT 207.500000 329.590000 249.500000 330.410000 ;
      RECT 157.500000 329.590000 199.500000 330.410000 ;
      RECT 107.500000 329.590000 149.500000 330.410000 ;
      RECT 57.500000 329.590000 99.500000 330.410000 ;
      RECT 15.500000 329.590000 49.500000 330.410000 ;
      RECT 1183.500000 328.410000 1186.000000 331.590000 ;
      RECT 1169.500000 328.410000 1170.500000 329.590000 ;
      RECT 1116.500000 328.410000 1149.500000 329.590000 ;
      RECT 1107.500000 328.410000 1108.500000 329.590000 ;
      RECT 1066.500000 328.410000 1099.500000 329.590000 ;
      RECT 1057.500000 328.410000 1058.500000 329.590000 ;
      RECT 1016.500000 328.410000 1049.500000 329.590000 ;
      RECT 1007.500000 328.410000 1008.500000 329.590000 ;
      RECT 966.500000 328.410000 999.500000 329.590000 ;
      RECT 957.500000 328.410000 958.500000 329.590000 ;
      RECT 916.500000 328.410000 949.500000 329.590000 ;
      RECT 907.500000 328.410000 908.500000 329.590000 ;
      RECT 866.500000 328.410000 899.500000 329.590000 ;
      RECT 857.500000 328.410000 858.500000 329.590000 ;
      RECT 816.500000 328.410000 849.500000 329.590000 ;
      RECT 807.500000 328.410000 808.500000 329.590000 ;
      RECT 766.500000 328.410000 799.500000 329.590000 ;
      RECT 757.500000 328.410000 758.500000 329.590000 ;
      RECT 716.500000 328.410000 749.500000 329.590000 ;
      RECT 707.500000 328.410000 708.500000 329.590000 ;
      RECT 666.500000 328.410000 699.500000 329.590000 ;
      RECT 657.500000 328.410000 658.500000 329.590000 ;
      RECT 616.500000 328.410000 649.500000 329.590000 ;
      RECT 607.500000 328.410000 608.500000 329.590000 ;
      RECT 566.500000 328.410000 599.500000 329.590000 ;
      RECT 557.500000 328.410000 558.500000 329.590000 ;
      RECT 516.500000 328.410000 549.500000 329.590000 ;
      RECT 507.500000 328.410000 508.500000 329.590000 ;
      RECT 466.500000 328.410000 499.500000 329.590000 ;
      RECT 457.500000 328.410000 458.500000 329.590000 ;
      RECT 416.500000 328.410000 449.500000 329.590000 ;
      RECT 407.500000 328.410000 408.500000 329.590000 ;
      RECT 366.500000 328.410000 399.500000 329.590000 ;
      RECT 357.500000 328.410000 358.500000 329.590000 ;
      RECT 316.500000 328.410000 349.500000 329.590000 ;
      RECT 307.500000 328.410000 308.500000 329.590000 ;
      RECT 266.500000 328.410000 299.500000 329.590000 ;
      RECT 257.500000 328.410000 258.500000 329.590000 ;
      RECT 216.500000 328.410000 249.500000 329.590000 ;
      RECT 207.500000 328.410000 208.500000 329.590000 ;
      RECT 166.500000 328.410000 199.500000 329.590000 ;
      RECT 157.500000 328.410000 158.500000 329.590000 ;
      RECT 116.500000 328.410000 149.500000 329.590000 ;
      RECT 107.500000 328.410000 108.500000 329.590000 ;
      RECT 66.500000 328.410000 99.500000 329.590000 ;
      RECT 57.500000 328.410000 58.500000 329.590000 ;
      RECT 29.500000 328.410000 49.500000 329.590000 ;
      RECT 15.500000 328.410000 16.500000 329.590000 ;
      RECT 0.000000 328.410000 2.500000 331.590000 ;
      RECT 1169.500000 327.590000 1186.000000 328.410000 ;
      RECT 1116.500000 327.590000 1156.500000 328.410000 ;
      RECT 1066.500000 327.590000 1108.500000 328.410000 ;
      RECT 1016.500000 327.590000 1058.500000 328.410000 ;
      RECT 966.500000 327.590000 1008.500000 328.410000 ;
      RECT 916.500000 327.590000 958.500000 328.410000 ;
      RECT 866.500000 327.590000 908.500000 328.410000 ;
      RECT 816.500000 327.590000 858.500000 328.410000 ;
      RECT 766.500000 327.590000 808.500000 328.410000 ;
      RECT 716.500000 327.590000 758.500000 328.410000 ;
      RECT 666.500000 327.590000 708.500000 328.410000 ;
      RECT 616.500000 327.590000 658.500000 328.410000 ;
      RECT 566.500000 327.590000 608.500000 328.410000 ;
      RECT 516.500000 327.590000 558.500000 328.410000 ;
      RECT 466.500000 327.590000 508.500000 328.410000 ;
      RECT 416.500000 327.590000 458.500000 328.410000 ;
      RECT 366.500000 327.590000 408.500000 328.410000 ;
      RECT 316.500000 327.590000 358.500000 328.410000 ;
      RECT 266.500000 327.590000 308.500000 328.410000 ;
      RECT 216.500000 327.590000 258.500000 328.410000 ;
      RECT 166.500000 327.590000 208.500000 328.410000 ;
      RECT 116.500000 327.590000 158.500000 328.410000 ;
      RECT 66.500000 327.590000 108.500000 328.410000 ;
      RECT 29.500000 327.590000 58.500000 328.410000 ;
      RECT 0.000000 327.590000 16.500000 328.410000 ;
      RECT 1169.500000 326.410000 1170.500000 327.590000 ;
      RECT 1116.500000 326.410000 1149.500000 327.590000 ;
      RECT 1107.500000 326.410000 1108.500000 327.590000 ;
      RECT 1066.500000 326.410000 1099.500000 327.590000 ;
      RECT 1057.500000 326.410000 1058.500000 327.590000 ;
      RECT 1016.500000 326.410000 1049.500000 327.590000 ;
      RECT 1007.500000 326.410000 1008.500000 327.590000 ;
      RECT 966.500000 326.410000 999.500000 327.590000 ;
      RECT 957.500000 326.410000 958.500000 327.590000 ;
      RECT 916.500000 326.410000 949.500000 327.590000 ;
      RECT 907.500000 326.410000 908.500000 327.590000 ;
      RECT 866.500000 326.410000 899.500000 327.590000 ;
      RECT 857.500000 326.410000 858.500000 327.590000 ;
      RECT 816.500000 326.410000 849.500000 327.590000 ;
      RECT 807.500000 326.410000 808.500000 327.590000 ;
      RECT 766.500000 326.410000 799.500000 327.590000 ;
      RECT 757.500000 326.410000 758.500000 327.590000 ;
      RECT 716.500000 326.410000 749.500000 327.590000 ;
      RECT 707.500000 326.410000 708.500000 327.590000 ;
      RECT 666.500000 326.410000 699.500000 327.590000 ;
      RECT 657.500000 326.410000 658.500000 327.590000 ;
      RECT 616.500000 326.410000 649.500000 327.590000 ;
      RECT 607.500000 326.410000 608.500000 327.590000 ;
      RECT 566.500000 326.410000 599.500000 327.590000 ;
      RECT 557.500000 326.410000 558.500000 327.590000 ;
      RECT 516.500000 326.410000 549.500000 327.590000 ;
      RECT 507.500000 326.410000 508.500000 327.590000 ;
      RECT 466.500000 326.410000 499.500000 327.590000 ;
      RECT 457.500000 326.410000 458.500000 327.590000 ;
      RECT 416.500000 326.410000 449.500000 327.590000 ;
      RECT 407.500000 326.410000 408.500000 327.590000 ;
      RECT 366.500000 326.410000 399.500000 327.590000 ;
      RECT 357.500000 326.410000 358.500000 327.590000 ;
      RECT 316.500000 326.410000 349.500000 327.590000 ;
      RECT 307.500000 326.410000 308.500000 327.590000 ;
      RECT 266.500000 326.410000 299.500000 327.590000 ;
      RECT 257.500000 326.410000 258.500000 327.590000 ;
      RECT 216.500000 326.410000 249.500000 327.590000 ;
      RECT 207.500000 326.410000 208.500000 327.590000 ;
      RECT 166.500000 326.410000 199.500000 327.590000 ;
      RECT 157.500000 326.410000 158.500000 327.590000 ;
      RECT 116.500000 326.410000 149.500000 327.590000 ;
      RECT 107.500000 326.410000 108.500000 327.590000 ;
      RECT 66.500000 326.410000 99.500000 327.590000 ;
      RECT 57.500000 326.410000 58.500000 327.590000 ;
      RECT 29.500000 326.410000 49.500000 327.590000 ;
      RECT 15.500000 326.410000 16.500000 327.590000 ;
      RECT 1157.500000 325.590000 1170.500000 326.410000 ;
      RECT 1107.500000 325.590000 1149.500000 326.410000 ;
      RECT 1057.500000 325.590000 1099.500000 326.410000 ;
      RECT 1007.500000 325.590000 1049.500000 326.410000 ;
      RECT 957.500000 325.590000 999.500000 326.410000 ;
      RECT 907.500000 325.590000 949.500000 326.410000 ;
      RECT 857.500000 325.590000 899.500000 326.410000 ;
      RECT 807.500000 325.590000 849.500000 326.410000 ;
      RECT 757.500000 325.590000 799.500000 326.410000 ;
      RECT 707.500000 325.590000 749.500000 326.410000 ;
      RECT 657.500000 325.590000 699.500000 326.410000 ;
      RECT 607.500000 325.590000 649.500000 326.410000 ;
      RECT 557.500000 325.590000 599.500000 326.410000 ;
      RECT 507.500000 325.590000 549.500000 326.410000 ;
      RECT 457.500000 325.590000 499.500000 326.410000 ;
      RECT 407.500000 325.590000 449.500000 326.410000 ;
      RECT 357.500000 325.590000 399.500000 326.410000 ;
      RECT 307.500000 325.590000 349.500000 326.410000 ;
      RECT 257.500000 325.590000 299.500000 326.410000 ;
      RECT 207.500000 325.590000 249.500000 326.410000 ;
      RECT 157.500000 325.590000 199.500000 326.410000 ;
      RECT 107.500000 325.590000 149.500000 326.410000 ;
      RECT 57.500000 325.590000 99.500000 326.410000 ;
      RECT 15.500000 325.590000 49.500000 326.410000 ;
      RECT 1183.500000 324.410000 1186.000000 327.590000 ;
      RECT 1169.500000 324.410000 1170.500000 325.590000 ;
      RECT 1116.500000 324.410000 1149.500000 325.590000 ;
      RECT 1107.500000 324.410000 1108.500000 325.590000 ;
      RECT 1066.500000 324.410000 1099.500000 325.590000 ;
      RECT 1057.500000 324.410000 1058.500000 325.590000 ;
      RECT 1016.500000 324.410000 1049.500000 325.590000 ;
      RECT 1007.500000 324.410000 1008.500000 325.590000 ;
      RECT 966.500000 324.410000 999.500000 325.590000 ;
      RECT 957.500000 324.410000 958.500000 325.590000 ;
      RECT 916.500000 324.410000 949.500000 325.590000 ;
      RECT 907.500000 324.410000 908.500000 325.590000 ;
      RECT 866.500000 324.410000 899.500000 325.590000 ;
      RECT 857.500000 324.410000 858.500000 325.590000 ;
      RECT 816.500000 324.410000 849.500000 325.590000 ;
      RECT 807.500000 324.410000 808.500000 325.590000 ;
      RECT 766.500000 324.410000 799.500000 325.590000 ;
      RECT 757.500000 324.410000 758.500000 325.590000 ;
      RECT 716.500000 324.410000 749.500000 325.590000 ;
      RECT 707.500000 324.410000 708.500000 325.590000 ;
      RECT 666.500000 324.410000 699.500000 325.590000 ;
      RECT 657.500000 324.410000 658.500000 325.590000 ;
      RECT 616.500000 324.410000 649.500000 325.590000 ;
      RECT 607.500000 324.410000 608.500000 325.590000 ;
      RECT 566.500000 324.410000 599.500000 325.590000 ;
      RECT 557.500000 324.410000 558.500000 325.590000 ;
      RECT 516.500000 324.410000 549.500000 325.590000 ;
      RECT 507.500000 324.410000 508.500000 325.590000 ;
      RECT 466.500000 324.410000 499.500000 325.590000 ;
      RECT 457.500000 324.410000 458.500000 325.590000 ;
      RECT 416.500000 324.410000 449.500000 325.590000 ;
      RECT 407.500000 324.410000 408.500000 325.590000 ;
      RECT 366.500000 324.410000 399.500000 325.590000 ;
      RECT 357.500000 324.410000 358.500000 325.590000 ;
      RECT 316.500000 324.410000 349.500000 325.590000 ;
      RECT 307.500000 324.410000 308.500000 325.590000 ;
      RECT 266.500000 324.410000 299.500000 325.590000 ;
      RECT 257.500000 324.410000 258.500000 325.590000 ;
      RECT 216.500000 324.410000 249.500000 325.590000 ;
      RECT 207.500000 324.410000 208.500000 325.590000 ;
      RECT 166.500000 324.410000 199.500000 325.590000 ;
      RECT 157.500000 324.410000 158.500000 325.590000 ;
      RECT 116.500000 324.410000 149.500000 325.590000 ;
      RECT 107.500000 324.410000 108.500000 325.590000 ;
      RECT 66.500000 324.410000 99.500000 325.590000 ;
      RECT 57.500000 324.410000 58.500000 325.590000 ;
      RECT 29.500000 324.410000 49.500000 325.590000 ;
      RECT 15.500000 324.410000 16.500000 325.590000 ;
      RECT 0.000000 324.410000 2.500000 327.590000 ;
      RECT 1169.500000 323.590000 1186.000000 324.410000 ;
      RECT 1116.500000 323.590000 1156.500000 324.410000 ;
      RECT 1066.500000 323.590000 1108.500000 324.410000 ;
      RECT 1016.500000 323.590000 1058.500000 324.410000 ;
      RECT 966.500000 323.590000 1008.500000 324.410000 ;
      RECT 916.500000 323.590000 958.500000 324.410000 ;
      RECT 866.500000 323.590000 908.500000 324.410000 ;
      RECT 816.500000 323.590000 858.500000 324.410000 ;
      RECT 766.500000 323.590000 808.500000 324.410000 ;
      RECT 716.500000 323.590000 758.500000 324.410000 ;
      RECT 666.500000 323.590000 708.500000 324.410000 ;
      RECT 616.500000 323.590000 658.500000 324.410000 ;
      RECT 566.500000 323.590000 608.500000 324.410000 ;
      RECT 516.500000 323.590000 558.500000 324.410000 ;
      RECT 466.500000 323.590000 508.500000 324.410000 ;
      RECT 416.500000 323.590000 458.500000 324.410000 ;
      RECT 366.500000 323.590000 408.500000 324.410000 ;
      RECT 316.500000 323.590000 358.500000 324.410000 ;
      RECT 266.500000 323.590000 308.500000 324.410000 ;
      RECT 216.500000 323.590000 258.500000 324.410000 ;
      RECT 166.500000 323.590000 208.500000 324.410000 ;
      RECT 116.500000 323.590000 158.500000 324.410000 ;
      RECT 66.500000 323.590000 108.500000 324.410000 ;
      RECT 29.500000 323.590000 58.500000 324.410000 ;
      RECT 0.000000 323.590000 16.500000 324.410000 ;
      RECT 1169.500000 322.410000 1170.500000 323.590000 ;
      RECT 1116.500000 322.410000 1149.500000 323.590000 ;
      RECT 1107.500000 322.410000 1108.500000 323.590000 ;
      RECT 1066.500000 322.410000 1099.500000 323.590000 ;
      RECT 1057.500000 322.410000 1058.500000 323.590000 ;
      RECT 1016.500000 322.410000 1049.500000 323.590000 ;
      RECT 1007.500000 322.410000 1008.500000 323.590000 ;
      RECT 966.500000 322.410000 999.500000 323.590000 ;
      RECT 957.500000 322.410000 958.500000 323.590000 ;
      RECT 916.500000 322.410000 949.500000 323.590000 ;
      RECT 907.500000 322.410000 908.500000 323.590000 ;
      RECT 866.500000 322.410000 899.500000 323.590000 ;
      RECT 857.500000 322.410000 858.500000 323.590000 ;
      RECT 816.500000 322.410000 849.500000 323.590000 ;
      RECT 807.500000 322.410000 808.500000 323.590000 ;
      RECT 766.500000 322.410000 799.500000 323.590000 ;
      RECT 757.500000 322.410000 758.500000 323.590000 ;
      RECT 716.500000 322.410000 749.500000 323.590000 ;
      RECT 707.500000 322.410000 708.500000 323.590000 ;
      RECT 666.500000 322.410000 699.500000 323.590000 ;
      RECT 657.500000 322.410000 658.500000 323.590000 ;
      RECT 616.500000 322.410000 649.500000 323.590000 ;
      RECT 607.500000 322.410000 608.500000 323.590000 ;
      RECT 566.500000 322.410000 599.500000 323.590000 ;
      RECT 557.500000 322.410000 558.500000 323.590000 ;
      RECT 516.500000 322.410000 549.500000 323.590000 ;
      RECT 507.500000 322.410000 508.500000 323.590000 ;
      RECT 466.500000 322.410000 499.500000 323.590000 ;
      RECT 457.500000 322.410000 458.500000 323.590000 ;
      RECT 416.500000 322.410000 449.500000 323.590000 ;
      RECT 407.500000 322.410000 408.500000 323.590000 ;
      RECT 366.500000 322.410000 399.500000 323.590000 ;
      RECT 357.500000 322.410000 358.500000 323.590000 ;
      RECT 316.500000 322.410000 349.500000 323.590000 ;
      RECT 307.500000 322.410000 308.500000 323.590000 ;
      RECT 266.500000 322.410000 299.500000 323.590000 ;
      RECT 257.500000 322.410000 258.500000 323.590000 ;
      RECT 216.500000 322.410000 249.500000 323.590000 ;
      RECT 207.500000 322.410000 208.500000 323.590000 ;
      RECT 166.500000 322.410000 199.500000 323.590000 ;
      RECT 157.500000 322.410000 158.500000 323.590000 ;
      RECT 116.500000 322.410000 149.500000 323.590000 ;
      RECT 107.500000 322.410000 108.500000 323.590000 ;
      RECT 66.500000 322.410000 99.500000 323.590000 ;
      RECT 57.500000 322.410000 58.500000 323.590000 ;
      RECT 29.500000 322.410000 49.500000 323.590000 ;
      RECT 15.500000 322.410000 16.500000 323.590000 ;
      RECT 1157.500000 321.590000 1170.500000 322.410000 ;
      RECT 1107.500000 321.590000 1149.500000 322.410000 ;
      RECT 1057.500000 321.590000 1099.500000 322.410000 ;
      RECT 1007.500000 321.590000 1049.500000 322.410000 ;
      RECT 957.500000 321.590000 999.500000 322.410000 ;
      RECT 907.500000 321.590000 949.500000 322.410000 ;
      RECT 857.500000 321.590000 899.500000 322.410000 ;
      RECT 807.500000 321.590000 849.500000 322.410000 ;
      RECT 757.500000 321.590000 799.500000 322.410000 ;
      RECT 707.500000 321.590000 749.500000 322.410000 ;
      RECT 657.500000 321.590000 699.500000 322.410000 ;
      RECT 607.500000 321.590000 649.500000 322.410000 ;
      RECT 557.500000 321.590000 599.500000 322.410000 ;
      RECT 507.500000 321.590000 549.500000 322.410000 ;
      RECT 457.500000 321.590000 499.500000 322.410000 ;
      RECT 407.500000 321.590000 449.500000 322.410000 ;
      RECT 357.500000 321.590000 399.500000 322.410000 ;
      RECT 307.500000 321.590000 349.500000 322.410000 ;
      RECT 257.500000 321.590000 299.500000 322.410000 ;
      RECT 207.500000 321.590000 249.500000 322.410000 ;
      RECT 157.500000 321.590000 199.500000 322.410000 ;
      RECT 107.500000 321.590000 149.500000 322.410000 ;
      RECT 57.500000 321.590000 99.500000 322.410000 ;
      RECT 15.500000 321.590000 49.500000 322.410000 ;
      RECT 1183.500000 320.410000 1186.000000 323.590000 ;
      RECT 1169.500000 320.410000 1170.500000 321.590000 ;
      RECT 1116.500000 320.410000 1149.500000 321.590000 ;
      RECT 1107.500000 320.410000 1108.500000 321.590000 ;
      RECT 1066.500000 320.410000 1099.500000 321.590000 ;
      RECT 1057.500000 320.410000 1058.500000 321.590000 ;
      RECT 1016.500000 320.410000 1049.500000 321.590000 ;
      RECT 1007.500000 320.410000 1008.500000 321.590000 ;
      RECT 966.500000 320.410000 999.500000 321.590000 ;
      RECT 957.500000 320.410000 958.500000 321.590000 ;
      RECT 916.500000 320.410000 949.500000 321.590000 ;
      RECT 907.500000 320.410000 908.500000 321.590000 ;
      RECT 866.500000 320.410000 899.500000 321.590000 ;
      RECT 857.500000 320.410000 858.500000 321.590000 ;
      RECT 816.500000 320.410000 849.500000 321.590000 ;
      RECT 807.500000 320.410000 808.500000 321.590000 ;
      RECT 766.500000 320.410000 799.500000 321.590000 ;
      RECT 757.500000 320.410000 758.500000 321.590000 ;
      RECT 716.500000 320.410000 749.500000 321.590000 ;
      RECT 707.500000 320.410000 708.500000 321.590000 ;
      RECT 666.500000 320.410000 699.500000 321.590000 ;
      RECT 657.500000 320.410000 658.500000 321.590000 ;
      RECT 616.500000 320.410000 649.500000 321.590000 ;
      RECT 607.500000 320.410000 608.500000 321.590000 ;
      RECT 566.500000 320.410000 599.500000 321.590000 ;
      RECT 557.500000 320.410000 558.500000 321.590000 ;
      RECT 516.500000 320.410000 549.500000 321.590000 ;
      RECT 507.500000 320.410000 508.500000 321.590000 ;
      RECT 466.500000 320.410000 499.500000 321.590000 ;
      RECT 457.500000 320.410000 458.500000 321.590000 ;
      RECT 416.500000 320.410000 449.500000 321.590000 ;
      RECT 407.500000 320.410000 408.500000 321.590000 ;
      RECT 366.500000 320.410000 399.500000 321.590000 ;
      RECT 357.500000 320.410000 358.500000 321.590000 ;
      RECT 316.500000 320.410000 349.500000 321.590000 ;
      RECT 307.500000 320.410000 308.500000 321.590000 ;
      RECT 266.500000 320.410000 299.500000 321.590000 ;
      RECT 257.500000 320.410000 258.500000 321.590000 ;
      RECT 216.500000 320.410000 249.500000 321.590000 ;
      RECT 207.500000 320.410000 208.500000 321.590000 ;
      RECT 166.500000 320.410000 199.500000 321.590000 ;
      RECT 157.500000 320.410000 158.500000 321.590000 ;
      RECT 116.500000 320.410000 149.500000 321.590000 ;
      RECT 107.500000 320.410000 108.500000 321.590000 ;
      RECT 66.500000 320.410000 99.500000 321.590000 ;
      RECT 57.500000 320.410000 58.500000 321.590000 ;
      RECT 29.500000 320.410000 49.500000 321.590000 ;
      RECT 15.500000 320.410000 16.500000 321.590000 ;
      RECT 0.000000 320.410000 2.500000 323.590000 ;
      RECT 1169.500000 319.590000 1186.000000 320.410000 ;
      RECT 1116.500000 319.590000 1156.500000 320.410000 ;
      RECT 1066.500000 319.590000 1108.500000 320.410000 ;
      RECT 1016.500000 319.590000 1058.500000 320.410000 ;
      RECT 966.500000 319.590000 1008.500000 320.410000 ;
      RECT 916.500000 319.590000 958.500000 320.410000 ;
      RECT 866.500000 319.590000 908.500000 320.410000 ;
      RECT 816.500000 319.590000 858.500000 320.410000 ;
      RECT 766.500000 319.590000 808.500000 320.410000 ;
      RECT 716.500000 319.590000 758.500000 320.410000 ;
      RECT 666.500000 319.590000 708.500000 320.410000 ;
      RECT 616.500000 319.590000 658.500000 320.410000 ;
      RECT 566.500000 319.590000 608.500000 320.410000 ;
      RECT 516.500000 319.590000 558.500000 320.410000 ;
      RECT 466.500000 319.590000 508.500000 320.410000 ;
      RECT 366.500000 319.590000 408.500000 320.410000 ;
      RECT 316.500000 319.590000 358.500000 320.410000 ;
      RECT 266.500000 319.590000 308.500000 320.410000 ;
      RECT 216.500000 319.590000 258.500000 320.410000 ;
      RECT 166.500000 319.590000 208.500000 320.410000 ;
      RECT 116.500000 319.590000 158.500000 320.410000 ;
      RECT 66.500000 319.590000 108.500000 320.410000 ;
      RECT 29.500000 319.590000 58.500000 320.410000 ;
      RECT 0.000000 319.590000 16.500000 320.410000 ;
      RECT 416.500000 318.605000 458.500000 320.410000 ;
      RECT 1169.500000 318.410000 1170.500000 319.590000 ;
      RECT 1116.500000 318.410000 1149.500000 319.590000 ;
      RECT 1107.500000 318.410000 1108.500000 319.590000 ;
      RECT 1066.500000 318.410000 1099.500000 319.590000 ;
      RECT 1057.500000 318.410000 1058.500000 319.590000 ;
      RECT 1016.500000 318.410000 1049.500000 319.590000 ;
      RECT 1007.500000 318.410000 1008.500000 319.590000 ;
      RECT 966.500000 318.410000 999.500000 319.590000 ;
      RECT 957.500000 318.410000 958.500000 319.590000 ;
      RECT 916.500000 318.410000 949.500000 319.590000 ;
      RECT 907.500000 318.410000 908.500000 319.590000 ;
      RECT 866.500000 318.410000 899.500000 319.590000 ;
      RECT 857.500000 318.410000 858.500000 319.590000 ;
      RECT 816.500000 318.410000 849.500000 319.590000 ;
      RECT 807.500000 318.410000 808.500000 319.590000 ;
      RECT 766.500000 318.410000 799.500000 319.590000 ;
      RECT 757.500000 318.410000 758.500000 319.590000 ;
      RECT 716.500000 318.410000 749.500000 319.590000 ;
      RECT 707.500000 318.410000 708.500000 319.590000 ;
      RECT 666.500000 318.410000 699.500000 319.590000 ;
      RECT 657.500000 318.410000 658.500000 319.590000 ;
      RECT 616.500000 318.410000 649.500000 319.590000 ;
      RECT 607.500000 318.410000 608.500000 319.590000 ;
      RECT 566.500000 318.410000 599.500000 319.590000 ;
      RECT 557.500000 318.410000 558.500000 319.590000 ;
      RECT 516.500000 318.410000 549.500000 319.590000 ;
      RECT 507.500000 318.410000 508.500000 319.590000 ;
      RECT 466.500000 318.410000 499.500000 319.590000 ;
      RECT 457.500000 318.410000 458.500000 318.605000 ;
      RECT 416.500000 318.410000 449.500000 318.605000 ;
      RECT 407.500000 318.410000 408.500000 319.590000 ;
      RECT 366.500000 318.410000 399.500000 319.590000 ;
      RECT 357.500000 318.410000 358.500000 319.590000 ;
      RECT 316.500000 318.410000 349.500000 319.590000 ;
      RECT 307.500000 318.410000 308.500000 319.590000 ;
      RECT 266.500000 318.410000 299.500000 319.590000 ;
      RECT 257.500000 318.410000 258.500000 319.590000 ;
      RECT 216.500000 318.410000 249.500000 319.590000 ;
      RECT 207.500000 318.410000 208.500000 319.590000 ;
      RECT 166.500000 318.410000 199.500000 319.590000 ;
      RECT 157.500000 318.410000 158.500000 319.590000 ;
      RECT 116.500000 318.410000 149.500000 319.590000 ;
      RECT 107.500000 318.410000 108.500000 319.590000 ;
      RECT 66.500000 318.410000 99.500000 319.590000 ;
      RECT 57.500000 318.410000 58.500000 319.590000 ;
      RECT 29.500000 318.410000 49.500000 319.590000 ;
      RECT 15.500000 318.410000 16.500000 319.590000 ;
      RECT 1157.500000 317.590000 1170.500000 318.410000 ;
      RECT 1107.500000 317.590000 1149.500000 318.410000 ;
      RECT 1057.500000 317.590000 1099.500000 318.410000 ;
      RECT 1007.500000 317.590000 1049.500000 318.410000 ;
      RECT 957.500000 317.590000 999.500000 318.410000 ;
      RECT 907.500000 317.590000 949.500000 318.410000 ;
      RECT 857.500000 317.590000 899.500000 318.410000 ;
      RECT 807.500000 317.590000 849.500000 318.410000 ;
      RECT 757.500000 317.590000 799.500000 318.410000 ;
      RECT 707.500000 317.590000 749.500000 318.410000 ;
      RECT 657.500000 317.590000 699.500000 318.410000 ;
      RECT 607.500000 317.590000 649.500000 318.410000 ;
      RECT 557.500000 317.590000 599.500000 318.410000 ;
      RECT 507.500000 317.590000 549.500000 318.410000 ;
      RECT 407.500000 317.590000 449.500000 318.410000 ;
      RECT 357.500000 317.590000 399.500000 318.410000 ;
      RECT 307.500000 317.590000 349.500000 318.410000 ;
      RECT 257.500000 317.590000 299.500000 318.410000 ;
      RECT 207.500000 317.590000 249.500000 318.410000 ;
      RECT 157.500000 317.590000 199.500000 318.410000 ;
      RECT 107.500000 317.590000 149.500000 318.410000 ;
      RECT 57.500000 317.590000 99.500000 318.410000 ;
      RECT 15.500000 317.590000 49.500000 318.410000 ;
      RECT 1183.500000 316.410000 1186.000000 319.590000 ;
      RECT 1169.500000 316.410000 1170.500000 317.590000 ;
      RECT 1116.500000 316.410000 1149.500000 317.590000 ;
      RECT 1107.500000 316.410000 1108.500000 317.590000 ;
      RECT 1066.500000 316.410000 1099.500000 317.590000 ;
      RECT 1057.500000 316.410000 1058.500000 317.590000 ;
      RECT 1016.500000 316.410000 1049.500000 317.590000 ;
      RECT 1007.500000 316.410000 1008.500000 317.590000 ;
      RECT 966.500000 316.410000 999.500000 317.590000 ;
      RECT 957.500000 316.410000 958.500000 317.590000 ;
      RECT 916.500000 316.410000 949.500000 317.590000 ;
      RECT 907.500000 316.410000 908.500000 317.590000 ;
      RECT 866.500000 316.410000 899.500000 317.590000 ;
      RECT 857.500000 316.410000 858.500000 317.590000 ;
      RECT 816.500000 316.410000 849.500000 317.590000 ;
      RECT 807.500000 316.410000 808.500000 317.590000 ;
      RECT 766.500000 316.410000 799.500000 317.590000 ;
      RECT 757.500000 316.410000 758.500000 317.590000 ;
      RECT 716.500000 316.410000 749.500000 317.590000 ;
      RECT 707.500000 316.410000 708.500000 317.590000 ;
      RECT 666.500000 316.410000 699.500000 317.590000 ;
      RECT 657.500000 316.410000 658.500000 317.590000 ;
      RECT 616.500000 316.410000 649.500000 317.590000 ;
      RECT 607.500000 316.410000 608.500000 317.590000 ;
      RECT 566.500000 316.410000 599.500000 317.590000 ;
      RECT 557.500000 316.410000 558.500000 317.590000 ;
      RECT 516.500000 316.410000 549.500000 317.590000 ;
      RECT 507.500000 316.410000 508.500000 317.590000 ;
      RECT 457.500000 316.410000 499.500000 318.410000 ;
      RECT 407.500000 316.410000 408.500000 317.590000 ;
      RECT 366.500000 316.410000 399.500000 317.590000 ;
      RECT 357.500000 316.410000 358.500000 317.590000 ;
      RECT 316.500000 316.410000 349.500000 317.590000 ;
      RECT 307.500000 316.410000 308.500000 317.590000 ;
      RECT 266.500000 316.410000 299.500000 317.590000 ;
      RECT 257.500000 316.410000 258.500000 317.590000 ;
      RECT 216.500000 316.410000 249.500000 317.590000 ;
      RECT 207.500000 316.410000 208.500000 317.590000 ;
      RECT 166.500000 316.410000 199.500000 317.590000 ;
      RECT 157.500000 316.410000 158.500000 317.590000 ;
      RECT 116.500000 316.410000 149.500000 317.590000 ;
      RECT 107.500000 316.410000 108.500000 317.590000 ;
      RECT 66.500000 316.410000 99.500000 317.590000 ;
      RECT 57.500000 316.410000 58.500000 317.590000 ;
      RECT 29.500000 316.410000 49.500000 317.590000 ;
      RECT 15.500000 316.410000 16.500000 317.590000 ;
      RECT 0.000000 316.410000 2.500000 319.590000 ;
      RECT 1169.500000 315.590000 1186.000000 316.410000 ;
      RECT 1116.500000 315.590000 1156.500000 316.410000 ;
      RECT 1066.500000 315.590000 1108.500000 316.410000 ;
      RECT 1016.500000 315.590000 1058.500000 316.410000 ;
      RECT 966.500000 315.590000 1008.500000 316.410000 ;
      RECT 916.500000 315.590000 958.500000 316.410000 ;
      RECT 866.500000 315.590000 908.500000 316.410000 ;
      RECT 816.500000 315.590000 858.500000 316.410000 ;
      RECT 766.500000 315.590000 808.500000 316.410000 ;
      RECT 716.500000 315.590000 758.500000 316.410000 ;
      RECT 666.500000 315.590000 708.500000 316.410000 ;
      RECT 616.500000 315.590000 658.500000 316.410000 ;
      RECT 566.500000 315.590000 608.500000 316.410000 ;
      RECT 516.500000 315.590000 558.500000 316.410000 ;
      RECT 457.500000 315.590000 508.500000 316.410000 ;
      RECT 366.500000 315.590000 408.500000 316.410000 ;
      RECT 316.500000 315.590000 358.500000 316.410000 ;
      RECT 266.500000 315.590000 308.500000 316.410000 ;
      RECT 216.500000 315.590000 258.500000 316.410000 ;
      RECT 166.500000 315.590000 208.500000 316.410000 ;
      RECT 116.500000 315.590000 158.500000 316.410000 ;
      RECT 66.500000 315.590000 108.500000 316.410000 ;
      RECT 29.500000 315.590000 58.500000 316.410000 ;
      RECT 0.000000 315.590000 16.500000 316.410000 ;
      RECT 457.500000 314.605000 499.500000 315.590000 ;
      RECT 416.500000 314.605000 449.500000 317.590000 ;
      RECT 1169.500000 314.410000 1170.500000 315.590000 ;
      RECT 1116.500000 314.410000 1149.500000 315.590000 ;
      RECT 1107.500000 314.410000 1108.500000 315.590000 ;
      RECT 1066.500000 314.410000 1099.500000 315.590000 ;
      RECT 1057.500000 314.410000 1058.500000 315.590000 ;
      RECT 1016.500000 314.410000 1049.500000 315.590000 ;
      RECT 1007.500000 314.410000 1008.500000 315.590000 ;
      RECT 966.500000 314.410000 999.500000 315.590000 ;
      RECT 957.500000 314.410000 958.500000 315.590000 ;
      RECT 916.500000 314.410000 949.500000 315.590000 ;
      RECT 907.500000 314.410000 908.500000 315.590000 ;
      RECT 866.500000 314.410000 899.500000 315.590000 ;
      RECT 857.500000 314.410000 858.500000 315.590000 ;
      RECT 816.500000 314.410000 849.500000 315.590000 ;
      RECT 807.500000 314.410000 808.500000 315.590000 ;
      RECT 766.500000 314.410000 799.500000 315.590000 ;
      RECT 757.500000 314.410000 758.500000 315.590000 ;
      RECT 716.500000 314.410000 749.500000 315.590000 ;
      RECT 707.500000 314.410000 708.500000 315.590000 ;
      RECT 666.500000 314.410000 699.500000 315.590000 ;
      RECT 657.500000 314.410000 658.500000 315.590000 ;
      RECT 616.500000 314.410000 649.500000 315.590000 ;
      RECT 607.500000 314.410000 608.500000 315.590000 ;
      RECT 566.500000 314.410000 599.500000 315.590000 ;
      RECT 557.500000 314.410000 558.500000 315.590000 ;
      RECT 516.500000 314.410000 549.500000 315.590000 ;
      RECT 507.500000 314.410000 508.500000 315.590000 ;
      RECT 416.500000 314.410000 499.500000 314.605000 ;
      RECT 407.500000 314.410000 408.500000 315.590000 ;
      RECT 366.500000 314.410000 399.500000 315.590000 ;
      RECT 357.500000 314.410000 358.500000 315.590000 ;
      RECT 316.500000 314.410000 349.500000 315.590000 ;
      RECT 307.500000 314.410000 308.500000 315.590000 ;
      RECT 266.500000 314.410000 299.500000 315.590000 ;
      RECT 257.500000 314.410000 258.500000 315.590000 ;
      RECT 216.500000 314.410000 249.500000 315.590000 ;
      RECT 207.500000 314.410000 208.500000 315.590000 ;
      RECT 166.500000 314.410000 199.500000 315.590000 ;
      RECT 157.500000 314.410000 158.500000 315.590000 ;
      RECT 116.500000 314.410000 149.500000 315.590000 ;
      RECT 107.500000 314.410000 108.500000 315.590000 ;
      RECT 66.500000 314.410000 99.500000 315.590000 ;
      RECT 57.500000 314.410000 58.500000 315.590000 ;
      RECT 29.500000 314.410000 49.500000 315.590000 ;
      RECT 15.500000 314.410000 16.500000 315.590000 ;
      RECT 1157.500000 313.590000 1170.500000 314.410000 ;
      RECT 1107.500000 313.590000 1149.500000 314.410000 ;
      RECT 1057.500000 313.590000 1099.500000 314.410000 ;
      RECT 1007.500000 313.590000 1049.500000 314.410000 ;
      RECT 957.500000 313.590000 999.500000 314.410000 ;
      RECT 907.500000 313.590000 949.500000 314.410000 ;
      RECT 857.500000 313.590000 899.500000 314.410000 ;
      RECT 807.500000 313.590000 849.500000 314.410000 ;
      RECT 757.500000 313.590000 799.500000 314.410000 ;
      RECT 707.500000 313.590000 749.500000 314.410000 ;
      RECT 657.500000 313.590000 699.500000 314.410000 ;
      RECT 607.500000 313.590000 649.500000 314.410000 ;
      RECT 557.500000 313.590000 599.500000 314.410000 ;
      RECT 507.500000 313.590000 549.500000 314.410000 ;
      RECT 407.500000 313.590000 499.500000 314.410000 ;
      RECT 357.500000 313.590000 399.500000 314.410000 ;
      RECT 307.500000 313.590000 349.500000 314.410000 ;
      RECT 257.500000 313.590000 299.500000 314.410000 ;
      RECT 207.500000 313.590000 249.500000 314.410000 ;
      RECT 157.500000 313.590000 199.500000 314.410000 ;
      RECT 107.500000 313.590000 149.500000 314.410000 ;
      RECT 57.500000 313.590000 99.500000 314.410000 ;
      RECT 15.500000 313.590000 49.500000 314.410000 ;
      RECT 1183.500000 312.410000 1186.000000 315.590000 ;
      RECT 1169.500000 312.410000 1170.500000 313.590000 ;
      RECT 1116.500000 312.410000 1149.500000 313.590000 ;
      RECT 1107.500000 312.410000 1108.500000 313.590000 ;
      RECT 1066.500000 312.410000 1099.500000 313.590000 ;
      RECT 1057.500000 312.410000 1058.500000 313.590000 ;
      RECT 1016.500000 312.410000 1049.500000 313.590000 ;
      RECT 1007.500000 312.410000 1008.500000 313.590000 ;
      RECT 966.500000 312.410000 999.500000 313.590000 ;
      RECT 957.500000 312.410000 958.500000 313.590000 ;
      RECT 916.500000 312.410000 949.500000 313.590000 ;
      RECT 907.500000 312.410000 908.500000 313.590000 ;
      RECT 866.500000 312.410000 899.500000 313.590000 ;
      RECT 857.500000 312.410000 858.500000 313.590000 ;
      RECT 816.500000 312.410000 849.500000 313.590000 ;
      RECT 807.500000 312.410000 808.500000 313.590000 ;
      RECT 766.500000 312.410000 799.500000 313.590000 ;
      RECT 757.500000 312.410000 758.500000 313.590000 ;
      RECT 716.500000 312.410000 749.500000 313.590000 ;
      RECT 707.500000 312.410000 708.500000 313.590000 ;
      RECT 666.500000 312.410000 699.500000 313.590000 ;
      RECT 657.500000 312.410000 658.500000 313.590000 ;
      RECT 616.500000 312.410000 649.500000 313.590000 ;
      RECT 607.500000 312.410000 608.500000 313.590000 ;
      RECT 566.500000 312.410000 599.500000 313.590000 ;
      RECT 557.500000 312.410000 558.500000 313.590000 ;
      RECT 516.500000 312.410000 549.500000 313.590000 ;
      RECT 507.500000 312.410000 508.500000 313.590000 ;
      RECT 416.500000 312.410000 499.500000 313.590000 ;
      RECT 407.500000 312.410000 408.500000 313.590000 ;
      RECT 366.500000 312.410000 399.500000 313.590000 ;
      RECT 357.500000 312.410000 358.500000 313.590000 ;
      RECT 316.500000 312.410000 349.500000 313.590000 ;
      RECT 307.500000 312.410000 308.500000 313.590000 ;
      RECT 266.500000 312.410000 299.500000 313.590000 ;
      RECT 257.500000 312.410000 258.500000 313.590000 ;
      RECT 216.500000 312.410000 249.500000 313.590000 ;
      RECT 207.500000 312.410000 208.500000 313.590000 ;
      RECT 166.500000 312.410000 199.500000 313.590000 ;
      RECT 157.500000 312.410000 158.500000 313.590000 ;
      RECT 116.500000 312.410000 149.500000 313.590000 ;
      RECT 107.500000 312.410000 108.500000 313.590000 ;
      RECT 66.500000 312.410000 99.500000 313.590000 ;
      RECT 57.500000 312.410000 58.500000 313.590000 ;
      RECT 29.500000 312.410000 49.500000 313.590000 ;
      RECT 15.500000 312.410000 16.500000 313.590000 ;
      RECT 0.000000 312.410000 2.500000 315.590000 ;
      RECT 1169.500000 311.590000 1186.000000 312.410000 ;
      RECT 1116.500000 311.590000 1156.500000 312.410000 ;
      RECT 1066.500000 311.590000 1108.500000 312.410000 ;
      RECT 1016.500000 311.590000 1058.500000 312.410000 ;
      RECT 966.500000 311.590000 1008.500000 312.410000 ;
      RECT 916.500000 311.590000 958.500000 312.410000 ;
      RECT 866.500000 311.590000 908.500000 312.410000 ;
      RECT 816.500000 311.590000 858.500000 312.410000 ;
      RECT 766.500000 311.590000 808.500000 312.410000 ;
      RECT 716.500000 311.590000 758.500000 312.410000 ;
      RECT 666.500000 311.590000 708.500000 312.410000 ;
      RECT 616.500000 311.590000 658.500000 312.410000 ;
      RECT 566.500000 311.590000 608.500000 312.410000 ;
      RECT 516.500000 311.590000 558.500000 312.410000 ;
      RECT 416.500000 311.590000 508.500000 312.410000 ;
      RECT 366.500000 311.590000 408.500000 312.410000 ;
      RECT 316.500000 311.590000 358.500000 312.410000 ;
      RECT 266.500000 311.590000 308.500000 312.410000 ;
      RECT 216.500000 311.590000 258.500000 312.410000 ;
      RECT 166.500000 311.590000 208.500000 312.410000 ;
      RECT 116.500000 311.590000 158.500000 312.410000 ;
      RECT 66.500000 311.590000 108.500000 312.410000 ;
      RECT 29.500000 311.590000 58.500000 312.410000 ;
      RECT 0.000000 311.590000 16.500000 312.410000 ;
      RECT 1169.500000 310.410000 1170.500000 311.590000 ;
      RECT 1116.500000 310.410000 1149.500000 311.590000 ;
      RECT 1107.500000 310.410000 1108.500000 311.590000 ;
      RECT 1066.500000 310.410000 1099.500000 311.590000 ;
      RECT 1057.500000 310.410000 1058.500000 311.590000 ;
      RECT 1016.500000 310.410000 1049.500000 311.590000 ;
      RECT 1007.500000 310.410000 1008.500000 311.590000 ;
      RECT 966.500000 310.410000 999.500000 311.590000 ;
      RECT 957.500000 310.410000 958.500000 311.590000 ;
      RECT 916.500000 310.410000 949.500000 311.590000 ;
      RECT 907.500000 310.410000 908.500000 311.590000 ;
      RECT 866.500000 310.410000 899.500000 311.590000 ;
      RECT 857.500000 310.410000 858.500000 311.590000 ;
      RECT 816.500000 310.410000 849.500000 311.590000 ;
      RECT 807.500000 310.410000 808.500000 311.590000 ;
      RECT 766.500000 310.410000 799.500000 311.590000 ;
      RECT 757.500000 310.410000 758.500000 311.590000 ;
      RECT 716.500000 310.410000 749.500000 311.590000 ;
      RECT 707.500000 310.410000 708.500000 311.590000 ;
      RECT 666.500000 310.410000 699.500000 311.590000 ;
      RECT 657.500000 310.410000 658.500000 311.590000 ;
      RECT 616.500000 310.410000 649.500000 311.590000 ;
      RECT 607.500000 310.410000 608.500000 311.590000 ;
      RECT 566.500000 310.410000 599.500000 311.590000 ;
      RECT 557.500000 310.410000 558.500000 311.590000 ;
      RECT 516.500000 310.410000 549.500000 311.590000 ;
      RECT 507.500000 310.410000 508.500000 311.590000 ;
      RECT 416.500000 310.410000 499.500000 311.590000 ;
      RECT 407.500000 310.410000 408.500000 311.590000 ;
      RECT 366.500000 310.410000 399.500000 311.590000 ;
      RECT 357.500000 310.410000 358.500000 311.590000 ;
      RECT 316.500000 310.410000 349.500000 311.590000 ;
      RECT 307.500000 310.410000 308.500000 311.590000 ;
      RECT 266.500000 310.410000 299.500000 311.590000 ;
      RECT 257.500000 310.410000 258.500000 311.590000 ;
      RECT 216.500000 310.410000 249.500000 311.590000 ;
      RECT 207.500000 310.410000 208.500000 311.590000 ;
      RECT 166.500000 310.410000 199.500000 311.590000 ;
      RECT 157.500000 310.410000 158.500000 311.590000 ;
      RECT 116.500000 310.410000 149.500000 311.590000 ;
      RECT 107.500000 310.410000 108.500000 311.590000 ;
      RECT 66.500000 310.410000 99.500000 311.590000 ;
      RECT 57.500000 310.410000 58.500000 311.590000 ;
      RECT 29.500000 310.410000 49.500000 311.590000 ;
      RECT 15.500000 310.410000 16.500000 311.590000 ;
      RECT 1157.500000 309.590000 1170.500000 310.410000 ;
      RECT 1107.500000 309.590000 1149.500000 310.410000 ;
      RECT 1057.500000 309.590000 1099.500000 310.410000 ;
      RECT 1007.500000 309.590000 1049.500000 310.410000 ;
      RECT 957.500000 309.590000 999.500000 310.410000 ;
      RECT 907.500000 309.590000 949.500000 310.410000 ;
      RECT 857.500000 309.590000 899.500000 310.410000 ;
      RECT 807.500000 309.590000 849.500000 310.410000 ;
      RECT 757.500000 309.590000 799.500000 310.410000 ;
      RECT 707.500000 309.590000 749.500000 310.410000 ;
      RECT 657.500000 309.590000 699.500000 310.410000 ;
      RECT 607.500000 309.590000 649.500000 310.410000 ;
      RECT 557.500000 309.590000 599.500000 310.410000 ;
      RECT 507.500000 309.590000 549.500000 310.410000 ;
      RECT 407.500000 309.590000 499.500000 310.410000 ;
      RECT 357.500000 309.590000 399.500000 310.410000 ;
      RECT 307.500000 309.590000 349.500000 310.410000 ;
      RECT 257.500000 309.590000 299.500000 310.410000 ;
      RECT 207.500000 309.590000 249.500000 310.410000 ;
      RECT 157.500000 309.590000 199.500000 310.410000 ;
      RECT 107.500000 309.590000 149.500000 310.410000 ;
      RECT 57.500000 309.590000 99.500000 310.410000 ;
      RECT 15.500000 309.590000 49.500000 310.410000 ;
      RECT 1183.500000 308.410000 1186.000000 311.590000 ;
      RECT 1169.500000 308.410000 1170.500000 309.590000 ;
      RECT 1116.500000 308.410000 1149.500000 309.590000 ;
      RECT 1107.500000 308.410000 1108.500000 309.590000 ;
      RECT 1066.500000 308.410000 1099.500000 309.590000 ;
      RECT 1057.500000 308.410000 1058.500000 309.590000 ;
      RECT 1016.500000 308.410000 1049.500000 309.590000 ;
      RECT 1007.500000 308.410000 1008.500000 309.590000 ;
      RECT 966.500000 308.410000 999.500000 309.590000 ;
      RECT 957.500000 308.410000 958.500000 309.590000 ;
      RECT 916.500000 308.410000 949.500000 309.590000 ;
      RECT 907.500000 308.410000 908.500000 309.590000 ;
      RECT 866.500000 308.410000 899.500000 309.590000 ;
      RECT 857.500000 308.410000 858.500000 309.590000 ;
      RECT 816.500000 308.410000 849.500000 309.590000 ;
      RECT 807.500000 308.410000 808.500000 309.590000 ;
      RECT 766.500000 308.410000 799.500000 309.590000 ;
      RECT 757.500000 308.410000 758.500000 309.590000 ;
      RECT 716.500000 308.410000 749.500000 309.590000 ;
      RECT 707.500000 308.410000 708.500000 309.590000 ;
      RECT 666.500000 308.410000 699.500000 309.590000 ;
      RECT 657.500000 308.410000 658.500000 309.590000 ;
      RECT 616.500000 308.410000 649.500000 309.590000 ;
      RECT 607.500000 308.410000 608.500000 309.590000 ;
      RECT 566.500000 308.410000 599.500000 309.590000 ;
      RECT 557.500000 308.410000 558.500000 309.590000 ;
      RECT 516.500000 308.410000 549.500000 309.590000 ;
      RECT 507.500000 308.410000 508.500000 309.590000 ;
      RECT 416.500000 308.410000 499.500000 309.590000 ;
      RECT 407.500000 308.410000 408.500000 309.590000 ;
      RECT 366.500000 308.410000 399.500000 309.590000 ;
      RECT 357.500000 308.410000 358.500000 309.590000 ;
      RECT 316.500000 308.410000 349.500000 309.590000 ;
      RECT 307.500000 308.410000 308.500000 309.590000 ;
      RECT 266.500000 308.410000 299.500000 309.590000 ;
      RECT 257.500000 308.410000 258.500000 309.590000 ;
      RECT 216.500000 308.410000 249.500000 309.590000 ;
      RECT 207.500000 308.410000 208.500000 309.590000 ;
      RECT 166.500000 308.410000 199.500000 309.590000 ;
      RECT 157.500000 308.410000 158.500000 309.590000 ;
      RECT 116.500000 308.410000 149.500000 309.590000 ;
      RECT 107.500000 308.410000 108.500000 309.590000 ;
      RECT 66.500000 308.410000 99.500000 309.590000 ;
      RECT 57.500000 308.410000 58.500000 309.590000 ;
      RECT 29.500000 308.410000 49.500000 309.590000 ;
      RECT 15.500000 308.410000 16.500000 309.590000 ;
      RECT 0.000000 308.410000 2.500000 311.590000 ;
      RECT 1169.500000 307.590000 1186.000000 308.410000 ;
      RECT 1116.500000 307.590000 1156.500000 308.410000 ;
      RECT 1066.500000 307.590000 1108.500000 308.410000 ;
      RECT 1016.500000 307.590000 1058.500000 308.410000 ;
      RECT 966.500000 307.590000 1008.500000 308.410000 ;
      RECT 916.500000 307.590000 958.500000 308.410000 ;
      RECT 866.500000 307.590000 908.500000 308.410000 ;
      RECT 816.500000 307.590000 858.500000 308.410000 ;
      RECT 766.500000 307.590000 808.500000 308.410000 ;
      RECT 716.500000 307.590000 758.500000 308.410000 ;
      RECT 666.500000 307.590000 708.500000 308.410000 ;
      RECT 616.500000 307.590000 658.500000 308.410000 ;
      RECT 566.500000 307.590000 608.500000 308.410000 ;
      RECT 516.500000 307.590000 558.500000 308.410000 ;
      RECT 416.500000 307.590000 508.500000 308.410000 ;
      RECT 366.500000 307.590000 408.500000 308.410000 ;
      RECT 316.500000 307.590000 358.500000 308.410000 ;
      RECT 266.500000 307.590000 308.500000 308.410000 ;
      RECT 216.500000 307.590000 258.500000 308.410000 ;
      RECT 166.500000 307.590000 208.500000 308.410000 ;
      RECT 116.500000 307.590000 158.500000 308.410000 ;
      RECT 66.500000 307.590000 108.500000 308.410000 ;
      RECT 29.500000 307.590000 58.500000 308.410000 ;
      RECT 0.000000 307.590000 16.500000 308.410000 ;
      RECT 1169.500000 306.410000 1170.500000 307.590000 ;
      RECT 1116.500000 306.410000 1149.500000 307.590000 ;
      RECT 1107.500000 306.410000 1108.500000 307.590000 ;
      RECT 1066.500000 306.410000 1099.500000 307.590000 ;
      RECT 1057.500000 306.410000 1058.500000 307.590000 ;
      RECT 1016.500000 306.410000 1049.500000 307.590000 ;
      RECT 1007.500000 306.410000 1008.500000 307.590000 ;
      RECT 966.500000 306.410000 999.500000 307.590000 ;
      RECT 957.500000 306.410000 958.500000 307.590000 ;
      RECT 916.500000 306.410000 949.500000 307.590000 ;
      RECT 907.500000 306.410000 908.500000 307.590000 ;
      RECT 866.500000 306.410000 899.500000 307.590000 ;
      RECT 857.500000 306.410000 858.500000 307.590000 ;
      RECT 816.500000 306.410000 849.500000 307.590000 ;
      RECT 807.500000 306.410000 808.500000 307.590000 ;
      RECT 766.500000 306.410000 799.500000 307.590000 ;
      RECT 757.500000 306.410000 758.500000 307.590000 ;
      RECT 716.500000 306.410000 749.500000 307.590000 ;
      RECT 707.500000 306.410000 708.500000 307.590000 ;
      RECT 666.500000 306.410000 699.500000 307.590000 ;
      RECT 657.500000 306.410000 658.500000 307.590000 ;
      RECT 616.500000 306.410000 649.500000 307.590000 ;
      RECT 607.500000 306.410000 608.500000 307.590000 ;
      RECT 566.500000 306.410000 599.500000 307.590000 ;
      RECT 557.500000 306.410000 558.500000 307.590000 ;
      RECT 516.500000 306.410000 549.500000 307.590000 ;
      RECT 507.500000 306.410000 508.500000 307.590000 ;
      RECT 416.500000 306.410000 499.500000 307.590000 ;
      RECT 407.500000 306.410000 408.500000 307.590000 ;
      RECT 366.500000 306.410000 399.500000 307.590000 ;
      RECT 357.500000 306.410000 358.500000 307.590000 ;
      RECT 316.500000 306.410000 349.500000 307.590000 ;
      RECT 307.500000 306.410000 308.500000 307.590000 ;
      RECT 266.500000 306.410000 299.500000 307.590000 ;
      RECT 257.500000 306.410000 258.500000 307.590000 ;
      RECT 216.500000 306.410000 249.500000 307.590000 ;
      RECT 207.500000 306.410000 208.500000 307.590000 ;
      RECT 166.500000 306.410000 199.500000 307.590000 ;
      RECT 157.500000 306.410000 158.500000 307.590000 ;
      RECT 116.500000 306.410000 149.500000 307.590000 ;
      RECT 107.500000 306.410000 108.500000 307.590000 ;
      RECT 66.500000 306.410000 99.500000 307.590000 ;
      RECT 57.500000 306.410000 58.500000 307.590000 ;
      RECT 29.500000 306.410000 49.500000 307.590000 ;
      RECT 15.500000 306.410000 16.500000 307.590000 ;
      RECT 1157.500000 305.590000 1170.500000 306.410000 ;
      RECT 1107.500000 305.590000 1149.500000 306.410000 ;
      RECT 1057.500000 305.590000 1099.500000 306.410000 ;
      RECT 1007.500000 305.590000 1049.500000 306.410000 ;
      RECT 957.500000 305.590000 999.500000 306.410000 ;
      RECT 907.500000 305.590000 949.500000 306.410000 ;
      RECT 857.500000 305.590000 899.500000 306.410000 ;
      RECT 807.500000 305.590000 849.500000 306.410000 ;
      RECT 757.500000 305.590000 799.500000 306.410000 ;
      RECT 707.500000 305.590000 749.500000 306.410000 ;
      RECT 657.500000 305.590000 699.500000 306.410000 ;
      RECT 607.500000 305.590000 649.500000 306.410000 ;
      RECT 557.500000 305.590000 599.500000 306.410000 ;
      RECT 507.500000 305.590000 549.500000 306.410000 ;
      RECT 407.500000 305.590000 499.500000 306.410000 ;
      RECT 357.500000 305.590000 399.500000 306.410000 ;
      RECT 307.500000 305.590000 349.500000 306.410000 ;
      RECT 257.500000 305.590000 299.500000 306.410000 ;
      RECT 207.500000 305.590000 249.500000 306.410000 ;
      RECT 157.500000 305.590000 199.500000 306.410000 ;
      RECT 107.500000 305.590000 149.500000 306.410000 ;
      RECT 57.500000 305.590000 99.500000 306.410000 ;
      RECT 15.500000 305.590000 49.500000 306.410000 ;
      RECT 1183.500000 304.410000 1186.000000 307.590000 ;
      RECT 1169.500000 304.410000 1170.500000 305.590000 ;
      RECT 1116.500000 304.410000 1149.500000 305.590000 ;
      RECT 1107.500000 304.410000 1108.500000 305.590000 ;
      RECT 1066.500000 304.410000 1099.500000 305.590000 ;
      RECT 1057.500000 304.410000 1058.500000 305.590000 ;
      RECT 1016.500000 304.410000 1049.500000 305.590000 ;
      RECT 1007.500000 304.410000 1008.500000 305.590000 ;
      RECT 966.500000 304.410000 999.500000 305.590000 ;
      RECT 957.500000 304.410000 958.500000 305.590000 ;
      RECT 916.500000 304.410000 949.500000 305.590000 ;
      RECT 907.500000 304.410000 908.500000 305.590000 ;
      RECT 866.500000 304.410000 899.500000 305.590000 ;
      RECT 857.500000 304.410000 858.500000 305.590000 ;
      RECT 816.500000 304.410000 849.500000 305.590000 ;
      RECT 807.500000 304.410000 808.500000 305.590000 ;
      RECT 766.500000 304.410000 799.500000 305.590000 ;
      RECT 757.500000 304.410000 758.500000 305.590000 ;
      RECT 716.500000 304.410000 749.500000 305.590000 ;
      RECT 707.500000 304.410000 708.500000 305.590000 ;
      RECT 666.500000 304.410000 699.500000 305.590000 ;
      RECT 657.500000 304.410000 658.500000 305.590000 ;
      RECT 616.500000 304.410000 649.500000 305.590000 ;
      RECT 607.500000 304.410000 608.500000 305.590000 ;
      RECT 566.500000 304.410000 599.500000 305.590000 ;
      RECT 557.500000 304.410000 558.500000 305.590000 ;
      RECT 516.500000 304.410000 549.500000 305.590000 ;
      RECT 507.500000 304.410000 508.500000 305.590000 ;
      RECT 416.500000 304.410000 499.500000 305.590000 ;
      RECT 407.500000 304.410000 408.500000 305.590000 ;
      RECT 366.500000 304.410000 399.500000 305.590000 ;
      RECT 357.500000 304.410000 358.500000 305.590000 ;
      RECT 316.500000 304.410000 349.500000 305.590000 ;
      RECT 307.500000 304.410000 308.500000 305.590000 ;
      RECT 266.500000 304.410000 299.500000 305.590000 ;
      RECT 257.500000 304.410000 258.500000 305.590000 ;
      RECT 216.500000 304.410000 249.500000 305.590000 ;
      RECT 207.500000 304.410000 208.500000 305.590000 ;
      RECT 166.500000 304.410000 199.500000 305.590000 ;
      RECT 157.500000 304.410000 158.500000 305.590000 ;
      RECT 116.500000 304.410000 149.500000 305.590000 ;
      RECT 107.500000 304.410000 108.500000 305.590000 ;
      RECT 66.500000 304.410000 99.500000 305.590000 ;
      RECT 57.500000 304.410000 58.500000 305.590000 ;
      RECT 29.500000 304.410000 49.500000 305.590000 ;
      RECT 15.500000 304.410000 16.500000 305.590000 ;
      RECT 0.000000 304.410000 2.500000 307.590000 ;
      RECT 416.500000 303.730000 508.500000 304.410000 ;
      RECT 1169.500000 303.590000 1186.000000 304.410000 ;
      RECT 1116.500000 303.590000 1156.500000 304.410000 ;
      RECT 1066.500000 303.590000 1108.500000 304.410000 ;
      RECT 1016.500000 303.590000 1058.500000 304.410000 ;
      RECT 966.500000 303.590000 1008.500000 304.410000 ;
      RECT 916.500000 303.590000 958.500000 304.410000 ;
      RECT 866.500000 303.590000 908.500000 304.410000 ;
      RECT 816.500000 303.590000 858.500000 304.410000 ;
      RECT 766.500000 303.590000 808.500000 304.410000 ;
      RECT 716.500000 303.590000 758.500000 304.410000 ;
      RECT 666.500000 303.590000 708.500000 304.410000 ;
      RECT 616.500000 303.590000 658.500000 304.410000 ;
      RECT 566.500000 303.590000 608.500000 304.410000 ;
      RECT 516.500000 303.590000 558.500000 304.410000 ;
      RECT 466.500000 303.590000 508.500000 303.730000 ;
      RECT 366.500000 303.590000 408.500000 304.410000 ;
      RECT 316.500000 303.590000 358.500000 304.410000 ;
      RECT 266.500000 303.590000 308.500000 304.410000 ;
      RECT 216.500000 303.590000 258.500000 304.410000 ;
      RECT 166.500000 303.590000 208.500000 304.410000 ;
      RECT 116.500000 303.590000 158.500000 304.410000 ;
      RECT 66.500000 303.590000 108.500000 304.410000 ;
      RECT 29.500000 303.590000 58.500000 304.410000 ;
      RECT 0.000000 303.590000 16.500000 304.410000 ;
      RECT 1169.500000 302.410000 1170.500000 303.590000 ;
      RECT 1116.500000 302.410000 1149.500000 303.590000 ;
      RECT 1107.500000 302.410000 1108.500000 303.590000 ;
      RECT 1066.500000 302.410000 1099.500000 303.590000 ;
      RECT 1057.500000 302.410000 1058.500000 303.590000 ;
      RECT 1016.500000 302.410000 1049.500000 303.590000 ;
      RECT 1007.500000 302.410000 1008.500000 303.590000 ;
      RECT 966.500000 302.410000 999.500000 303.590000 ;
      RECT 957.500000 302.410000 958.500000 303.590000 ;
      RECT 916.500000 302.410000 949.500000 303.590000 ;
      RECT 907.500000 302.410000 908.500000 303.590000 ;
      RECT 866.500000 302.410000 899.500000 303.590000 ;
      RECT 857.500000 302.410000 858.500000 303.590000 ;
      RECT 816.500000 302.410000 849.500000 303.590000 ;
      RECT 807.500000 302.410000 808.500000 303.590000 ;
      RECT 766.500000 302.410000 799.500000 303.590000 ;
      RECT 757.500000 302.410000 758.500000 303.590000 ;
      RECT 716.500000 302.410000 749.500000 303.590000 ;
      RECT 707.500000 302.410000 708.500000 303.590000 ;
      RECT 666.500000 302.410000 699.500000 303.590000 ;
      RECT 657.500000 302.410000 658.500000 303.590000 ;
      RECT 616.500000 302.410000 649.500000 303.590000 ;
      RECT 607.500000 302.410000 608.500000 303.590000 ;
      RECT 566.500000 302.410000 599.500000 303.590000 ;
      RECT 557.500000 302.410000 558.500000 303.590000 ;
      RECT 516.500000 302.410000 549.500000 303.590000 ;
      RECT 507.500000 302.410000 508.500000 303.590000 ;
      RECT 416.500000 302.410000 458.500000 303.730000 ;
      RECT 407.500000 302.410000 408.500000 303.590000 ;
      RECT 366.500000 302.410000 399.500000 303.590000 ;
      RECT 357.500000 302.410000 358.500000 303.590000 ;
      RECT 316.500000 302.410000 349.500000 303.590000 ;
      RECT 307.500000 302.410000 308.500000 303.590000 ;
      RECT 266.500000 302.410000 299.500000 303.590000 ;
      RECT 257.500000 302.410000 258.500000 303.590000 ;
      RECT 216.500000 302.410000 249.500000 303.590000 ;
      RECT 207.500000 302.410000 208.500000 303.590000 ;
      RECT 166.500000 302.410000 199.500000 303.590000 ;
      RECT 157.500000 302.410000 158.500000 303.590000 ;
      RECT 116.500000 302.410000 149.500000 303.590000 ;
      RECT 107.500000 302.410000 108.500000 303.590000 ;
      RECT 66.500000 302.410000 99.500000 303.590000 ;
      RECT 57.500000 302.410000 58.500000 303.590000 ;
      RECT 29.500000 302.410000 49.500000 303.590000 ;
      RECT 15.500000 302.410000 16.500000 303.590000 ;
      RECT 1157.500000 301.590000 1170.500000 302.410000 ;
      RECT 1107.500000 301.590000 1149.500000 302.410000 ;
      RECT 1057.500000 301.590000 1099.500000 302.410000 ;
      RECT 1007.500000 301.590000 1049.500000 302.410000 ;
      RECT 957.500000 301.590000 999.500000 302.410000 ;
      RECT 907.500000 301.590000 949.500000 302.410000 ;
      RECT 857.500000 301.590000 899.500000 302.410000 ;
      RECT 807.500000 301.590000 849.500000 302.410000 ;
      RECT 757.500000 301.590000 799.500000 302.410000 ;
      RECT 707.500000 301.590000 749.500000 302.410000 ;
      RECT 657.500000 301.590000 699.500000 302.410000 ;
      RECT 607.500000 301.590000 649.500000 302.410000 ;
      RECT 557.500000 301.590000 599.500000 302.410000 ;
      RECT 507.500000 301.590000 549.500000 302.410000 ;
      RECT 407.500000 301.590000 458.500000 302.410000 ;
      RECT 357.500000 301.590000 399.500000 302.410000 ;
      RECT 307.500000 301.590000 349.500000 302.410000 ;
      RECT 257.500000 301.590000 299.500000 302.410000 ;
      RECT 207.500000 301.590000 249.500000 302.410000 ;
      RECT 157.500000 301.590000 199.500000 302.410000 ;
      RECT 107.500000 301.590000 149.500000 302.410000 ;
      RECT 57.500000 301.590000 99.500000 302.410000 ;
      RECT 15.500000 301.590000 49.500000 302.410000 ;
      RECT 1183.500000 300.410000 1186.000000 303.590000 ;
      RECT 1169.500000 300.410000 1170.500000 301.590000 ;
      RECT 1116.500000 300.410000 1149.500000 301.590000 ;
      RECT 1107.500000 300.410000 1108.500000 301.590000 ;
      RECT 1066.500000 300.410000 1099.500000 301.590000 ;
      RECT 1057.500000 300.410000 1058.500000 301.590000 ;
      RECT 1016.500000 300.410000 1049.500000 301.590000 ;
      RECT 1007.500000 300.410000 1008.500000 301.590000 ;
      RECT 966.500000 300.410000 999.500000 301.590000 ;
      RECT 957.500000 300.410000 958.500000 301.590000 ;
      RECT 916.500000 300.410000 949.500000 301.590000 ;
      RECT 907.500000 300.410000 908.500000 301.590000 ;
      RECT 866.500000 300.410000 899.500000 301.590000 ;
      RECT 857.500000 300.410000 858.500000 301.590000 ;
      RECT 816.500000 300.410000 849.500000 301.590000 ;
      RECT 807.500000 300.410000 808.500000 301.590000 ;
      RECT 766.500000 300.410000 799.500000 301.590000 ;
      RECT 757.500000 300.410000 758.500000 301.590000 ;
      RECT 716.500000 300.410000 749.500000 301.590000 ;
      RECT 707.500000 300.410000 708.500000 301.590000 ;
      RECT 666.500000 300.410000 699.500000 301.590000 ;
      RECT 657.500000 300.410000 658.500000 301.590000 ;
      RECT 616.500000 300.410000 649.500000 301.590000 ;
      RECT 607.500000 300.410000 608.500000 301.590000 ;
      RECT 566.500000 300.410000 599.500000 301.590000 ;
      RECT 557.500000 300.410000 558.500000 301.590000 ;
      RECT 516.500000 300.410000 549.500000 301.590000 ;
      RECT 507.500000 300.410000 508.500000 301.590000 ;
      RECT 466.500000 300.410000 499.500000 303.590000 ;
      RECT 407.500000 300.410000 408.500000 301.590000 ;
      RECT 366.500000 300.410000 399.500000 301.590000 ;
      RECT 357.500000 300.410000 358.500000 301.590000 ;
      RECT 316.500000 300.410000 349.500000 301.590000 ;
      RECT 307.500000 300.410000 308.500000 301.590000 ;
      RECT 266.500000 300.410000 299.500000 301.590000 ;
      RECT 257.500000 300.410000 258.500000 301.590000 ;
      RECT 216.500000 300.410000 249.500000 301.590000 ;
      RECT 207.500000 300.410000 208.500000 301.590000 ;
      RECT 166.500000 300.410000 199.500000 301.590000 ;
      RECT 157.500000 300.410000 158.500000 301.590000 ;
      RECT 116.500000 300.410000 149.500000 301.590000 ;
      RECT 107.500000 300.410000 108.500000 301.590000 ;
      RECT 66.500000 300.410000 99.500000 301.590000 ;
      RECT 57.500000 300.410000 58.500000 301.590000 ;
      RECT 29.500000 300.410000 49.500000 301.590000 ;
      RECT 15.500000 300.410000 16.500000 301.590000 ;
      RECT 0.000000 300.410000 2.500000 303.590000 ;
      RECT 466.500000 299.730000 508.500000 300.410000 ;
      RECT 416.500000 299.730000 458.500000 301.590000 ;
      RECT 1169.500000 299.590000 1186.000000 300.410000 ;
      RECT 1116.500000 299.590000 1156.500000 300.410000 ;
      RECT 1066.500000 299.590000 1108.500000 300.410000 ;
      RECT 1016.500000 299.590000 1058.500000 300.410000 ;
      RECT 966.500000 299.590000 1008.500000 300.410000 ;
      RECT 916.500000 299.590000 958.500000 300.410000 ;
      RECT 866.500000 299.590000 908.500000 300.410000 ;
      RECT 816.500000 299.590000 858.500000 300.410000 ;
      RECT 766.500000 299.590000 808.500000 300.410000 ;
      RECT 716.500000 299.590000 758.500000 300.410000 ;
      RECT 666.500000 299.590000 708.500000 300.410000 ;
      RECT 616.500000 299.590000 658.500000 300.410000 ;
      RECT 566.500000 299.590000 608.500000 300.410000 ;
      RECT 516.500000 299.590000 558.500000 300.410000 ;
      RECT 416.500000 299.590000 508.500000 299.730000 ;
      RECT 366.500000 299.590000 408.500000 300.410000 ;
      RECT 316.500000 299.590000 358.500000 300.410000 ;
      RECT 266.500000 299.590000 308.500000 300.410000 ;
      RECT 216.500000 299.590000 258.500000 300.410000 ;
      RECT 166.500000 299.590000 208.500000 300.410000 ;
      RECT 116.500000 299.590000 158.500000 300.410000 ;
      RECT 66.500000 299.590000 108.500000 300.410000 ;
      RECT 29.500000 299.590000 58.500000 300.410000 ;
      RECT 0.000000 299.590000 16.500000 300.410000 ;
      RECT 1169.500000 298.410000 1170.500000 299.590000 ;
      RECT 1116.500000 298.410000 1149.500000 299.590000 ;
      RECT 1107.500000 298.410000 1108.500000 299.590000 ;
      RECT 1066.500000 298.410000 1099.500000 299.590000 ;
      RECT 1057.500000 298.410000 1058.500000 299.590000 ;
      RECT 1016.500000 298.410000 1049.500000 299.590000 ;
      RECT 1007.500000 298.410000 1008.500000 299.590000 ;
      RECT 966.500000 298.410000 999.500000 299.590000 ;
      RECT 957.500000 298.410000 958.500000 299.590000 ;
      RECT 916.500000 298.410000 949.500000 299.590000 ;
      RECT 907.500000 298.410000 908.500000 299.590000 ;
      RECT 866.500000 298.410000 899.500000 299.590000 ;
      RECT 857.500000 298.410000 858.500000 299.590000 ;
      RECT 816.500000 298.410000 849.500000 299.590000 ;
      RECT 807.500000 298.410000 808.500000 299.590000 ;
      RECT 766.500000 298.410000 799.500000 299.590000 ;
      RECT 757.500000 298.410000 758.500000 299.590000 ;
      RECT 716.500000 298.410000 749.500000 299.590000 ;
      RECT 707.500000 298.410000 708.500000 299.590000 ;
      RECT 666.500000 298.410000 699.500000 299.590000 ;
      RECT 657.500000 298.410000 658.500000 299.590000 ;
      RECT 616.500000 298.410000 649.500000 299.590000 ;
      RECT 607.500000 298.410000 608.500000 299.590000 ;
      RECT 566.500000 298.410000 599.500000 299.590000 ;
      RECT 557.500000 298.410000 558.500000 299.590000 ;
      RECT 516.500000 298.410000 549.500000 299.590000 ;
      RECT 507.500000 298.410000 508.500000 299.590000 ;
      RECT 416.500000 298.410000 449.500000 299.590000 ;
      RECT 407.500000 298.410000 408.500000 299.590000 ;
      RECT 366.500000 298.410000 399.500000 299.590000 ;
      RECT 357.500000 298.410000 358.500000 299.590000 ;
      RECT 316.500000 298.410000 349.500000 299.590000 ;
      RECT 307.500000 298.410000 308.500000 299.590000 ;
      RECT 266.500000 298.410000 299.500000 299.590000 ;
      RECT 257.500000 298.410000 258.500000 299.590000 ;
      RECT 216.500000 298.410000 249.500000 299.590000 ;
      RECT 207.500000 298.410000 208.500000 299.590000 ;
      RECT 166.500000 298.410000 199.500000 299.590000 ;
      RECT 157.500000 298.410000 158.500000 299.590000 ;
      RECT 116.500000 298.410000 149.500000 299.590000 ;
      RECT 107.500000 298.410000 108.500000 299.590000 ;
      RECT 66.500000 298.410000 99.500000 299.590000 ;
      RECT 57.500000 298.410000 58.500000 299.590000 ;
      RECT 29.500000 298.410000 49.500000 299.590000 ;
      RECT 15.500000 298.410000 16.500000 299.590000 ;
      RECT 1157.500000 297.590000 1170.500000 298.410000 ;
      RECT 1107.500000 297.590000 1149.500000 298.410000 ;
      RECT 1057.500000 297.590000 1099.500000 298.410000 ;
      RECT 1007.500000 297.590000 1049.500000 298.410000 ;
      RECT 957.500000 297.590000 999.500000 298.410000 ;
      RECT 907.500000 297.590000 949.500000 298.410000 ;
      RECT 857.500000 297.590000 899.500000 298.410000 ;
      RECT 807.500000 297.590000 849.500000 298.410000 ;
      RECT 757.500000 297.590000 799.500000 298.410000 ;
      RECT 707.500000 297.590000 749.500000 298.410000 ;
      RECT 657.500000 297.590000 699.500000 298.410000 ;
      RECT 607.500000 297.590000 649.500000 298.410000 ;
      RECT 557.500000 297.590000 599.500000 298.410000 ;
      RECT 507.500000 297.590000 549.500000 298.410000 ;
      RECT 457.500000 297.590000 499.500000 299.590000 ;
      RECT 407.500000 297.590000 449.500000 298.410000 ;
      RECT 357.500000 297.590000 399.500000 298.410000 ;
      RECT 307.500000 297.590000 349.500000 298.410000 ;
      RECT 257.500000 297.590000 299.500000 298.410000 ;
      RECT 207.500000 297.590000 249.500000 298.410000 ;
      RECT 157.500000 297.590000 199.500000 298.410000 ;
      RECT 107.500000 297.590000 149.500000 298.410000 ;
      RECT 57.500000 297.590000 99.500000 298.410000 ;
      RECT 15.500000 297.590000 49.500000 298.410000 ;
      RECT 1183.500000 296.410000 1186.000000 299.590000 ;
      RECT 1169.500000 296.410000 1170.500000 297.590000 ;
      RECT 1116.500000 296.410000 1149.500000 297.590000 ;
      RECT 1107.500000 296.410000 1108.500000 297.590000 ;
      RECT 1066.500000 296.410000 1099.500000 297.590000 ;
      RECT 1057.500000 296.410000 1058.500000 297.590000 ;
      RECT 1016.500000 296.410000 1049.500000 297.590000 ;
      RECT 1007.500000 296.410000 1008.500000 297.590000 ;
      RECT 966.500000 296.410000 999.500000 297.590000 ;
      RECT 957.500000 296.410000 958.500000 297.590000 ;
      RECT 916.500000 296.410000 949.500000 297.590000 ;
      RECT 907.500000 296.410000 908.500000 297.590000 ;
      RECT 866.500000 296.410000 899.500000 297.590000 ;
      RECT 857.500000 296.410000 858.500000 297.590000 ;
      RECT 816.500000 296.410000 849.500000 297.590000 ;
      RECT 807.500000 296.410000 808.500000 297.590000 ;
      RECT 766.500000 296.410000 799.500000 297.590000 ;
      RECT 757.500000 296.410000 758.500000 297.590000 ;
      RECT 716.500000 296.410000 749.500000 297.590000 ;
      RECT 707.500000 296.410000 708.500000 297.590000 ;
      RECT 666.500000 296.410000 699.500000 297.590000 ;
      RECT 657.500000 296.410000 658.500000 297.590000 ;
      RECT 616.500000 296.410000 649.500000 297.590000 ;
      RECT 607.500000 296.410000 608.500000 297.590000 ;
      RECT 566.500000 296.410000 599.500000 297.590000 ;
      RECT 557.500000 296.410000 558.500000 297.590000 ;
      RECT 516.500000 296.410000 549.500000 297.590000 ;
      RECT 507.500000 296.410000 508.500000 297.590000 ;
      RECT 466.500000 296.410000 499.500000 297.590000 ;
      RECT 457.500000 296.410000 458.500000 297.590000 ;
      RECT 416.500000 296.410000 449.500000 297.590000 ;
      RECT 407.500000 296.410000 408.500000 297.590000 ;
      RECT 366.500000 296.410000 399.500000 297.590000 ;
      RECT 357.500000 296.410000 358.500000 297.590000 ;
      RECT 316.500000 296.410000 349.500000 297.590000 ;
      RECT 307.500000 296.410000 308.500000 297.590000 ;
      RECT 266.500000 296.410000 299.500000 297.590000 ;
      RECT 257.500000 296.410000 258.500000 297.590000 ;
      RECT 216.500000 296.410000 249.500000 297.590000 ;
      RECT 207.500000 296.410000 208.500000 297.590000 ;
      RECT 166.500000 296.410000 199.500000 297.590000 ;
      RECT 157.500000 296.410000 158.500000 297.590000 ;
      RECT 116.500000 296.410000 149.500000 297.590000 ;
      RECT 107.500000 296.410000 108.500000 297.590000 ;
      RECT 66.500000 296.410000 99.500000 297.590000 ;
      RECT 57.500000 296.410000 58.500000 297.590000 ;
      RECT 29.500000 296.410000 49.500000 297.590000 ;
      RECT 15.500000 296.410000 16.500000 297.590000 ;
      RECT 0.000000 296.410000 2.500000 299.590000 ;
      RECT 1169.500000 295.590000 1186.000000 296.410000 ;
      RECT 1116.500000 295.590000 1156.500000 296.410000 ;
      RECT 1066.500000 295.590000 1108.500000 296.410000 ;
      RECT 1016.500000 295.590000 1058.500000 296.410000 ;
      RECT 966.500000 295.590000 1008.500000 296.410000 ;
      RECT 916.500000 295.590000 958.500000 296.410000 ;
      RECT 866.500000 295.590000 908.500000 296.410000 ;
      RECT 816.500000 295.590000 858.500000 296.410000 ;
      RECT 766.500000 295.590000 808.500000 296.410000 ;
      RECT 716.500000 295.590000 758.500000 296.410000 ;
      RECT 666.500000 295.590000 708.500000 296.410000 ;
      RECT 616.500000 295.590000 658.500000 296.410000 ;
      RECT 566.500000 295.590000 608.500000 296.410000 ;
      RECT 516.500000 295.590000 558.500000 296.410000 ;
      RECT 466.500000 295.590000 508.500000 296.410000 ;
      RECT 416.500000 295.590000 458.500000 296.410000 ;
      RECT 366.500000 295.590000 408.500000 296.410000 ;
      RECT 316.500000 295.590000 358.500000 296.410000 ;
      RECT 266.500000 295.590000 308.500000 296.410000 ;
      RECT 216.500000 295.590000 258.500000 296.410000 ;
      RECT 166.500000 295.590000 208.500000 296.410000 ;
      RECT 116.500000 295.590000 158.500000 296.410000 ;
      RECT 66.500000 295.590000 108.500000 296.410000 ;
      RECT 29.500000 295.590000 58.500000 296.410000 ;
      RECT 0.000000 295.590000 16.500000 296.410000 ;
      RECT 1169.500000 294.410000 1170.500000 295.590000 ;
      RECT 1116.500000 294.410000 1149.500000 295.590000 ;
      RECT 1107.500000 294.410000 1108.500000 295.590000 ;
      RECT 1066.500000 294.410000 1099.500000 295.590000 ;
      RECT 1057.500000 294.410000 1058.500000 295.590000 ;
      RECT 1016.500000 294.410000 1049.500000 295.590000 ;
      RECT 1007.500000 294.410000 1008.500000 295.590000 ;
      RECT 966.500000 294.410000 999.500000 295.590000 ;
      RECT 957.500000 294.410000 958.500000 295.590000 ;
      RECT 916.500000 294.410000 949.500000 295.590000 ;
      RECT 907.500000 294.410000 908.500000 295.590000 ;
      RECT 866.500000 294.410000 899.500000 295.590000 ;
      RECT 857.500000 294.410000 858.500000 295.590000 ;
      RECT 816.500000 294.410000 849.500000 295.590000 ;
      RECT 807.500000 294.410000 808.500000 295.590000 ;
      RECT 766.500000 294.410000 799.500000 295.590000 ;
      RECT 757.500000 294.410000 758.500000 295.590000 ;
      RECT 716.500000 294.410000 749.500000 295.590000 ;
      RECT 707.500000 294.410000 708.500000 295.590000 ;
      RECT 666.500000 294.410000 699.500000 295.590000 ;
      RECT 657.500000 294.410000 658.500000 295.590000 ;
      RECT 616.500000 294.410000 649.500000 295.590000 ;
      RECT 607.500000 294.410000 608.500000 295.590000 ;
      RECT 566.500000 294.410000 599.500000 295.590000 ;
      RECT 557.500000 294.410000 558.500000 295.590000 ;
      RECT 516.500000 294.410000 549.500000 295.590000 ;
      RECT 507.500000 294.410000 508.500000 295.590000 ;
      RECT 466.500000 294.410000 499.500000 295.590000 ;
      RECT 457.500000 294.410000 458.500000 295.590000 ;
      RECT 416.500000 294.410000 449.500000 295.590000 ;
      RECT 407.500000 294.410000 408.500000 295.590000 ;
      RECT 366.500000 294.410000 399.500000 295.590000 ;
      RECT 357.500000 294.410000 358.500000 295.590000 ;
      RECT 316.500000 294.410000 349.500000 295.590000 ;
      RECT 307.500000 294.410000 308.500000 295.590000 ;
      RECT 266.500000 294.410000 299.500000 295.590000 ;
      RECT 257.500000 294.410000 258.500000 295.590000 ;
      RECT 216.500000 294.410000 249.500000 295.590000 ;
      RECT 207.500000 294.410000 208.500000 295.590000 ;
      RECT 166.500000 294.410000 199.500000 295.590000 ;
      RECT 157.500000 294.410000 158.500000 295.590000 ;
      RECT 116.500000 294.410000 149.500000 295.590000 ;
      RECT 107.500000 294.410000 108.500000 295.590000 ;
      RECT 66.500000 294.410000 99.500000 295.590000 ;
      RECT 57.500000 294.410000 58.500000 295.590000 ;
      RECT 29.500000 294.410000 49.500000 295.590000 ;
      RECT 15.500000 294.410000 16.500000 295.590000 ;
      RECT 1157.500000 293.590000 1170.500000 294.410000 ;
      RECT 1107.500000 293.590000 1149.500000 294.410000 ;
      RECT 1057.500000 293.590000 1099.500000 294.410000 ;
      RECT 1007.500000 293.590000 1049.500000 294.410000 ;
      RECT 957.500000 293.590000 999.500000 294.410000 ;
      RECT 907.500000 293.590000 949.500000 294.410000 ;
      RECT 857.500000 293.590000 899.500000 294.410000 ;
      RECT 807.500000 293.590000 849.500000 294.410000 ;
      RECT 757.500000 293.590000 799.500000 294.410000 ;
      RECT 707.500000 293.590000 749.500000 294.410000 ;
      RECT 657.500000 293.590000 699.500000 294.410000 ;
      RECT 607.500000 293.590000 649.500000 294.410000 ;
      RECT 557.500000 293.590000 599.500000 294.410000 ;
      RECT 507.500000 293.590000 549.500000 294.410000 ;
      RECT 457.500000 293.590000 499.500000 294.410000 ;
      RECT 407.500000 293.590000 449.500000 294.410000 ;
      RECT 357.500000 293.590000 399.500000 294.410000 ;
      RECT 307.500000 293.590000 349.500000 294.410000 ;
      RECT 257.500000 293.590000 299.500000 294.410000 ;
      RECT 207.500000 293.590000 249.500000 294.410000 ;
      RECT 157.500000 293.590000 199.500000 294.410000 ;
      RECT 107.500000 293.590000 149.500000 294.410000 ;
      RECT 57.500000 293.590000 99.500000 294.410000 ;
      RECT 15.500000 293.590000 49.500000 294.410000 ;
      RECT 1183.500000 292.410000 1186.000000 295.590000 ;
      RECT 1169.500000 292.410000 1170.500000 293.590000 ;
      RECT 1116.500000 292.410000 1149.500000 293.590000 ;
      RECT 1107.500000 292.410000 1108.500000 293.590000 ;
      RECT 1066.500000 292.410000 1099.500000 293.590000 ;
      RECT 1057.500000 292.410000 1058.500000 293.590000 ;
      RECT 1016.500000 292.410000 1049.500000 293.590000 ;
      RECT 1007.500000 292.410000 1008.500000 293.590000 ;
      RECT 966.500000 292.410000 999.500000 293.590000 ;
      RECT 957.500000 292.410000 958.500000 293.590000 ;
      RECT 916.500000 292.410000 949.500000 293.590000 ;
      RECT 907.500000 292.410000 908.500000 293.590000 ;
      RECT 866.500000 292.410000 899.500000 293.590000 ;
      RECT 857.500000 292.410000 858.500000 293.590000 ;
      RECT 816.500000 292.410000 849.500000 293.590000 ;
      RECT 807.500000 292.410000 808.500000 293.590000 ;
      RECT 766.500000 292.410000 799.500000 293.590000 ;
      RECT 757.500000 292.410000 758.500000 293.590000 ;
      RECT 716.500000 292.410000 749.500000 293.590000 ;
      RECT 707.500000 292.410000 708.500000 293.590000 ;
      RECT 666.500000 292.410000 699.500000 293.590000 ;
      RECT 657.500000 292.410000 658.500000 293.590000 ;
      RECT 616.500000 292.410000 649.500000 293.590000 ;
      RECT 607.500000 292.410000 608.500000 293.590000 ;
      RECT 566.500000 292.410000 599.500000 293.590000 ;
      RECT 557.500000 292.410000 558.500000 293.590000 ;
      RECT 516.500000 292.410000 549.500000 293.590000 ;
      RECT 507.500000 292.410000 508.500000 293.590000 ;
      RECT 466.500000 292.410000 499.500000 293.590000 ;
      RECT 457.500000 292.410000 458.500000 293.590000 ;
      RECT 416.500000 292.410000 449.500000 293.590000 ;
      RECT 407.500000 292.410000 408.500000 293.590000 ;
      RECT 366.500000 292.410000 399.500000 293.590000 ;
      RECT 357.500000 292.410000 358.500000 293.590000 ;
      RECT 316.500000 292.410000 349.500000 293.590000 ;
      RECT 307.500000 292.410000 308.500000 293.590000 ;
      RECT 266.500000 292.410000 299.500000 293.590000 ;
      RECT 257.500000 292.410000 258.500000 293.590000 ;
      RECT 216.500000 292.410000 249.500000 293.590000 ;
      RECT 207.500000 292.410000 208.500000 293.590000 ;
      RECT 166.500000 292.410000 199.500000 293.590000 ;
      RECT 157.500000 292.410000 158.500000 293.590000 ;
      RECT 116.500000 292.410000 149.500000 293.590000 ;
      RECT 107.500000 292.410000 108.500000 293.590000 ;
      RECT 66.500000 292.410000 99.500000 293.590000 ;
      RECT 57.500000 292.410000 58.500000 293.590000 ;
      RECT 29.500000 292.410000 49.500000 293.590000 ;
      RECT 15.500000 292.410000 16.500000 293.590000 ;
      RECT 0.000000 292.410000 2.500000 295.590000 ;
      RECT 1169.500000 291.590000 1186.000000 292.410000 ;
      RECT 1116.500000 291.590000 1156.500000 292.410000 ;
      RECT 1066.500000 291.590000 1108.500000 292.410000 ;
      RECT 1016.500000 291.590000 1058.500000 292.410000 ;
      RECT 966.500000 291.590000 1008.500000 292.410000 ;
      RECT 916.500000 291.590000 958.500000 292.410000 ;
      RECT 866.500000 291.590000 908.500000 292.410000 ;
      RECT 816.500000 291.590000 858.500000 292.410000 ;
      RECT 766.500000 291.590000 808.500000 292.410000 ;
      RECT 716.500000 291.590000 758.500000 292.410000 ;
      RECT 666.500000 291.590000 708.500000 292.410000 ;
      RECT 616.500000 291.590000 658.500000 292.410000 ;
      RECT 566.500000 291.590000 608.500000 292.410000 ;
      RECT 516.500000 291.590000 558.500000 292.410000 ;
      RECT 466.500000 291.590000 508.500000 292.410000 ;
      RECT 416.500000 291.590000 458.500000 292.410000 ;
      RECT 366.500000 291.590000 408.500000 292.410000 ;
      RECT 316.500000 291.590000 358.500000 292.410000 ;
      RECT 266.500000 291.590000 308.500000 292.410000 ;
      RECT 216.500000 291.590000 258.500000 292.410000 ;
      RECT 166.500000 291.590000 208.500000 292.410000 ;
      RECT 116.500000 291.590000 158.500000 292.410000 ;
      RECT 66.500000 291.590000 108.500000 292.410000 ;
      RECT 29.500000 291.590000 58.500000 292.410000 ;
      RECT 0.000000 291.590000 16.500000 292.410000 ;
      RECT 1169.500000 290.410000 1170.500000 291.590000 ;
      RECT 1116.500000 290.410000 1149.500000 291.590000 ;
      RECT 1107.500000 290.410000 1108.500000 291.590000 ;
      RECT 1066.500000 290.410000 1099.500000 291.590000 ;
      RECT 1057.500000 290.410000 1058.500000 291.590000 ;
      RECT 1016.500000 290.410000 1049.500000 291.590000 ;
      RECT 1007.500000 290.410000 1008.500000 291.590000 ;
      RECT 966.500000 290.410000 999.500000 291.590000 ;
      RECT 957.500000 290.410000 958.500000 291.590000 ;
      RECT 916.500000 290.410000 949.500000 291.590000 ;
      RECT 907.500000 290.410000 908.500000 291.590000 ;
      RECT 866.500000 290.410000 899.500000 291.590000 ;
      RECT 857.500000 290.410000 858.500000 291.590000 ;
      RECT 816.500000 290.410000 849.500000 291.590000 ;
      RECT 807.500000 290.410000 808.500000 291.590000 ;
      RECT 766.500000 290.410000 799.500000 291.590000 ;
      RECT 757.500000 290.410000 758.500000 291.590000 ;
      RECT 716.500000 290.410000 749.500000 291.590000 ;
      RECT 707.500000 290.410000 708.500000 291.590000 ;
      RECT 666.500000 290.410000 699.500000 291.590000 ;
      RECT 657.500000 290.410000 658.500000 291.590000 ;
      RECT 616.500000 290.410000 649.500000 291.590000 ;
      RECT 607.500000 290.410000 608.500000 291.590000 ;
      RECT 566.500000 290.410000 599.500000 291.590000 ;
      RECT 557.500000 290.410000 558.500000 291.590000 ;
      RECT 516.500000 290.410000 549.500000 291.590000 ;
      RECT 507.500000 290.410000 508.500000 291.590000 ;
      RECT 466.500000 290.410000 499.500000 291.590000 ;
      RECT 457.500000 290.410000 458.500000 291.590000 ;
      RECT 416.500000 290.410000 449.500000 291.590000 ;
      RECT 407.500000 290.410000 408.500000 291.590000 ;
      RECT 366.500000 290.410000 399.500000 291.590000 ;
      RECT 357.500000 290.410000 358.500000 291.590000 ;
      RECT 316.500000 290.410000 349.500000 291.590000 ;
      RECT 307.500000 290.410000 308.500000 291.590000 ;
      RECT 266.500000 290.410000 299.500000 291.590000 ;
      RECT 257.500000 290.410000 258.500000 291.590000 ;
      RECT 216.500000 290.410000 249.500000 291.590000 ;
      RECT 207.500000 290.410000 208.500000 291.590000 ;
      RECT 166.500000 290.410000 199.500000 291.590000 ;
      RECT 157.500000 290.410000 158.500000 291.590000 ;
      RECT 116.500000 290.410000 149.500000 291.590000 ;
      RECT 107.500000 290.410000 108.500000 291.590000 ;
      RECT 66.500000 290.410000 99.500000 291.590000 ;
      RECT 57.500000 290.410000 58.500000 291.590000 ;
      RECT 29.500000 290.410000 49.500000 291.590000 ;
      RECT 15.500000 290.410000 16.500000 291.590000 ;
      RECT 1157.500000 289.590000 1170.500000 290.410000 ;
      RECT 1107.500000 289.590000 1149.500000 290.410000 ;
      RECT 1057.500000 289.590000 1099.500000 290.410000 ;
      RECT 1007.500000 289.590000 1049.500000 290.410000 ;
      RECT 957.500000 289.590000 999.500000 290.410000 ;
      RECT 907.500000 289.590000 949.500000 290.410000 ;
      RECT 857.500000 289.590000 899.500000 290.410000 ;
      RECT 807.500000 289.590000 849.500000 290.410000 ;
      RECT 757.500000 289.590000 799.500000 290.410000 ;
      RECT 707.500000 289.590000 749.500000 290.410000 ;
      RECT 657.500000 289.590000 699.500000 290.410000 ;
      RECT 607.500000 289.590000 649.500000 290.410000 ;
      RECT 557.500000 289.590000 599.500000 290.410000 ;
      RECT 507.500000 289.590000 549.500000 290.410000 ;
      RECT 457.500000 289.590000 499.500000 290.410000 ;
      RECT 407.500000 289.590000 449.500000 290.410000 ;
      RECT 357.500000 289.590000 399.500000 290.410000 ;
      RECT 307.500000 289.590000 349.500000 290.410000 ;
      RECT 257.500000 289.590000 299.500000 290.410000 ;
      RECT 207.500000 289.590000 249.500000 290.410000 ;
      RECT 157.500000 289.590000 199.500000 290.410000 ;
      RECT 107.500000 289.590000 149.500000 290.410000 ;
      RECT 57.500000 289.590000 99.500000 290.410000 ;
      RECT 15.500000 289.590000 49.500000 290.410000 ;
      RECT 1183.500000 288.410000 1186.000000 291.590000 ;
      RECT 1169.500000 288.410000 1170.500000 289.590000 ;
      RECT 1116.500000 288.410000 1149.500000 289.590000 ;
      RECT 1107.500000 288.410000 1108.500000 289.590000 ;
      RECT 1066.500000 288.410000 1099.500000 289.590000 ;
      RECT 1057.500000 288.410000 1058.500000 289.590000 ;
      RECT 1016.500000 288.410000 1049.500000 289.590000 ;
      RECT 1007.500000 288.410000 1008.500000 289.590000 ;
      RECT 966.500000 288.410000 999.500000 289.590000 ;
      RECT 957.500000 288.410000 958.500000 289.590000 ;
      RECT 916.500000 288.410000 949.500000 289.590000 ;
      RECT 907.500000 288.410000 908.500000 289.590000 ;
      RECT 866.500000 288.410000 899.500000 289.590000 ;
      RECT 857.500000 288.410000 858.500000 289.590000 ;
      RECT 816.500000 288.410000 849.500000 289.590000 ;
      RECT 807.500000 288.410000 808.500000 289.590000 ;
      RECT 766.500000 288.410000 799.500000 289.590000 ;
      RECT 757.500000 288.410000 758.500000 289.590000 ;
      RECT 716.500000 288.410000 749.500000 289.590000 ;
      RECT 707.500000 288.410000 708.500000 289.590000 ;
      RECT 666.500000 288.410000 699.500000 289.590000 ;
      RECT 657.500000 288.410000 658.500000 289.590000 ;
      RECT 616.500000 288.410000 649.500000 289.590000 ;
      RECT 607.500000 288.410000 608.500000 289.590000 ;
      RECT 566.500000 288.410000 599.500000 289.590000 ;
      RECT 557.500000 288.410000 558.500000 289.590000 ;
      RECT 516.500000 288.410000 549.500000 289.590000 ;
      RECT 507.500000 288.410000 508.500000 289.590000 ;
      RECT 466.500000 288.410000 499.500000 289.590000 ;
      RECT 457.500000 288.410000 458.500000 289.590000 ;
      RECT 416.500000 288.410000 449.500000 289.590000 ;
      RECT 407.500000 288.410000 408.500000 289.590000 ;
      RECT 366.500000 288.410000 399.500000 289.590000 ;
      RECT 357.500000 288.410000 358.500000 289.590000 ;
      RECT 316.500000 288.410000 349.500000 289.590000 ;
      RECT 307.500000 288.410000 308.500000 289.590000 ;
      RECT 266.500000 288.410000 299.500000 289.590000 ;
      RECT 257.500000 288.410000 258.500000 289.590000 ;
      RECT 216.500000 288.410000 249.500000 289.590000 ;
      RECT 207.500000 288.410000 208.500000 289.590000 ;
      RECT 166.500000 288.410000 199.500000 289.590000 ;
      RECT 157.500000 288.410000 158.500000 289.590000 ;
      RECT 116.500000 288.410000 149.500000 289.590000 ;
      RECT 107.500000 288.410000 108.500000 289.590000 ;
      RECT 66.500000 288.410000 99.500000 289.590000 ;
      RECT 57.500000 288.410000 58.500000 289.590000 ;
      RECT 29.500000 288.410000 49.500000 289.590000 ;
      RECT 15.500000 288.410000 16.500000 289.590000 ;
      RECT 0.000000 288.410000 2.500000 291.590000 ;
      RECT 1169.500000 287.590000 1186.000000 288.410000 ;
      RECT 1116.500000 287.590000 1156.500000 288.410000 ;
      RECT 1066.500000 287.590000 1108.500000 288.410000 ;
      RECT 1016.500000 287.590000 1058.500000 288.410000 ;
      RECT 966.500000 287.590000 1008.500000 288.410000 ;
      RECT 916.500000 287.590000 958.500000 288.410000 ;
      RECT 866.500000 287.590000 908.500000 288.410000 ;
      RECT 816.500000 287.590000 858.500000 288.410000 ;
      RECT 766.500000 287.590000 808.500000 288.410000 ;
      RECT 716.500000 287.590000 758.500000 288.410000 ;
      RECT 666.500000 287.590000 708.500000 288.410000 ;
      RECT 616.500000 287.590000 658.500000 288.410000 ;
      RECT 566.500000 287.590000 608.500000 288.410000 ;
      RECT 516.500000 287.590000 558.500000 288.410000 ;
      RECT 466.500000 287.590000 508.500000 288.410000 ;
      RECT 416.500000 287.590000 458.500000 288.410000 ;
      RECT 366.500000 287.590000 408.500000 288.410000 ;
      RECT 316.500000 287.590000 358.500000 288.410000 ;
      RECT 266.500000 287.590000 308.500000 288.410000 ;
      RECT 216.500000 287.590000 258.500000 288.410000 ;
      RECT 166.500000 287.590000 208.500000 288.410000 ;
      RECT 116.500000 287.590000 158.500000 288.410000 ;
      RECT 66.500000 287.590000 108.500000 288.410000 ;
      RECT 29.500000 287.590000 58.500000 288.410000 ;
      RECT 0.000000 287.590000 16.500000 288.410000 ;
      RECT 1169.500000 286.410000 1170.500000 287.590000 ;
      RECT 1116.500000 286.410000 1149.500000 287.590000 ;
      RECT 1107.500000 286.410000 1108.500000 287.590000 ;
      RECT 1066.500000 286.410000 1099.500000 287.590000 ;
      RECT 1057.500000 286.410000 1058.500000 287.590000 ;
      RECT 1016.500000 286.410000 1049.500000 287.590000 ;
      RECT 1007.500000 286.410000 1008.500000 287.590000 ;
      RECT 966.500000 286.410000 999.500000 287.590000 ;
      RECT 957.500000 286.410000 958.500000 287.590000 ;
      RECT 916.500000 286.410000 949.500000 287.590000 ;
      RECT 907.500000 286.410000 908.500000 287.590000 ;
      RECT 866.500000 286.410000 899.500000 287.590000 ;
      RECT 857.500000 286.410000 858.500000 287.590000 ;
      RECT 816.500000 286.410000 849.500000 287.590000 ;
      RECT 807.500000 286.410000 808.500000 287.590000 ;
      RECT 766.500000 286.410000 799.500000 287.590000 ;
      RECT 757.500000 286.410000 758.500000 287.590000 ;
      RECT 716.500000 286.410000 749.500000 287.590000 ;
      RECT 707.500000 286.410000 708.500000 287.590000 ;
      RECT 666.500000 286.410000 699.500000 287.590000 ;
      RECT 657.500000 286.410000 658.500000 287.590000 ;
      RECT 616.500000 286.410000 649.500000 287.590000 ;
      RECT 607.500000 286.410000 608.500000 287.590000 ;
      RECT 566.500000 286.410000 599.500000 287.590000 ;
      RECT 557.500000 286.410000 558.500000 287.590000 ;
      RECT 516.500000 286.410000 549.500000 287.590000 ;
      RECT 507.500000 286.410000 508.500000 287.590000 ;
      RECT 466.500000 286.410000 499.500000 287.590000 ;
      RECT 457.500000 286.410000 458.500000 287.590000 ;
      RECT 416.500000 286.410000 449.500000 287.590000 ;
      RECT 407.500000 286.410000 408.500000 287.590000 ;
      RECT 366.500000 286.410000 399.500000 287.590000 ;
      RECT 357.500000 286.410000 358.500000 287.590000 ;
      RECT 316.500000 286.410000 349.500000 287.590000 ;
      RECT 307.500000 286.410000 308.500000 287.590000 ;
      RECT 266.500000 286.410000 299.500000 287.590000 ;
      RECT 257.500000 286.410000 258.500000 287.590000 ;
      RECT 216.500000 286.410000 249.500000 287.590000 ;
      RECT 207.500000 286.410000 208.500000 287.590000 ;
      RECT 166.500000 286.410000 199.500000 287.590000 ;
      RECT 157.500000 286.410000 158.500000 287.590000 ;
      RECT 116.500000 286.410000 149.500000 287.590000 ;
      RECT 107.500000 286.410000 108.500000 287.590000 ;
      RECT 66.500000 286.410000 99.500000 287.590000 ;
      RECT 57.500000 286.410000 58.500000 287.590000 ;
      RECT 29.500000 286.410000 49.500000 287.590000 ;
      RECT 15.500000 286.410000 16.500000 287.590000 ;
      RECT 1157.500000 285.590000 1170.500000 286.410000 ;
      RECT 1107.500000 285.590000 1149.500000 286.410000 ;
      RECT 1057.500000 285.590000 1099.500000 286.410000 ;
      RECT 1007.500000 285.590000 1049.500000 286.410000 ;
      RECT 957.500000 285.590000 999.500000 286.410000 ;
      RECT 907.500000 285.590000 949.500000 286.410000 ;
      RECT 857.500000 285.590000 899.500000 286.410000 ;
      RECT 807.500000 285.590000 849.500000 286.410000 ;
      RECT 757.500000 285.590000 799.500000 286.410000 ;
      RECT 707.500000 285.590000 749.500000 286.410000 ;
      RECT 657.500000 285.590000 699.500000 286.410000 ;
      RECT 607.500000 285.590000 649.500000 286.410000 ;
      RECT 557.500000 285.590000 599.500000 286.410000 ;
      RECT 507.500000 285.590000 549.500000 286.410000 ;
      RECT 457.500000 285.590000 499.500000 286.410000 ;
      RECT 407.500000 285.590000 449.500000 286.410000 ;
      RECT 357.500000 285.590000 399.500000 286.410000 ;
      RECT 307.500000 285.590000 349.500000 286.410000 ;
      RECT 257.500000 285.590000 299.500000 286.410000 ;
      RECT 207.500000 285.590000 249.500000 286.410000 ;
      RECT 157.500000 285.590000 199.500000 286.410000 ;
      RECT 107.500000 285.590000 149.500000 286.410000 ;
      RECT 57.500000 285.590000 99.500000 286.410000 ;
      RECT 15.500000 285.590000 49.500000 286.410000 ;
      RECT 1183.500000 284.410000 1186.000000 287.590000 ;
      RECT 1169.500000 284.410000 1170.500000 285.590000 ;
      RECT 1116.500000 284.410000 1149.500000 285.590000 ;
      RECT 1107.500000 284.410000 1108.500000 285.590000 ;
      RECT 1066.500000 284.410000 1099.500000 285.590000 ;
      RECT 1057.500000 284.410000 1058.500000 285.590000 ;
      RECT 1016.500000 284.410000 1049.500000 285.590000 ;
      RECT 1007.500000 284.410000 1008.500000 285.590000 ;
      RECT 966.500000 284.410000 999.500000 285.590000 ;
      RECT 957.500000 284.410000 958.500000 285.590000 ;
      RECT 916.500000 284.410000 949.500000 285.590000 ;
      RECT 907.500000 284.410000 908.500000 285.590000 ;
      RECT 866.500000 284.410000 899.500000 285.590000 ;
      RECT 857.500000 284.410000 858.500000 285.590000 ;
      RECT 816.500000 284.410000 849.500000 285.590000 ;
      RECT 807.500000 284.410000 808.500000 285.590000 ;
      RECT 766.500000 284.410000 799.500000 285.590000 ;
      RECT 757.500000 284.410000 758.500000 285.590000 ;
      RECT 716.500000 284.410000 749.500000 285.590000 ;
      RECT 707.500000 284.410000 708.500000 285.590000 ;
      RECT 666.500000 284.410000 699.500000 285.590000 ;
      RECT 657.500000 284.410000 658.500000 285.590000 ;
      RECT 616.500000 284.410000 649.500000 285.590000 ;
      RECT 607.500000 284.410000 608.500000 285.590000 ;
      RECT 566.500000 284.410000 599.500000 285.590000 ;
      RECT 557.500000 284.410000 558.500000 285.590000 ;
      RECT 516.500000 284.410000 549.500000 285.590000 ;
      RECT 507.500000 284.410000 508.500000 285.590000 ;
      RECT 466.500000 284.410000 499.500000 285.590000 ;
      RECT 457.500000 284.410000 458.500000 285.590000 ;
      RECT 416.500000 284.410000 449.500000 285.590000 ;
      RECT 407.500000 284.410000 408.500000 285.590000 ;
      RECT 366.500000 284.410000 399.500000 285.590000 ;
      RECT 357.500000 284.410000 358.500000 285.590000 ;
      RECT 316.500000 284.410000 349.500000 285.590000 ;
      RECT 307.500000 284.410000 308.500000 285.590000 ;
      RECT 266.500000 284.410000 299.500000 285.590000 ;
      RECT 257.500000 284.410000 258.500000 285.590000 ;
      RECT 216.500000 284.410000 249.500000 285.590000 ;
      RECT 207.500000 284.410000 208.500000 285.590000 ;
      RECT 166.500000 284.410000 199.500000 285.590000 ;
      RECT 157.500000 284.410000 158.500000 285.590000 ;
      RECT 116.500000 284.410000 149.500000 285.590000 ;
      RECT 107.500000 284.410000 108.500000 285.590000 ;
      RECT 66.500000 284.410000 99.500000 285.590000 ;
      RECT 57.500000 284.410000 58.500000 285.590000 ;
      RECT 29.500000 284.410000 49.500000 285.590000 ;
      RECT 15.500000 284.410000 16.500000 285.590000 ;
      RECT 0.000000 284.410000 2.500000 287.590000 ;
      RECT 1169.500000 283.590000 1186.000000 284.410000 ;
      RECT 1116.500000 283.590000 1156.500000 284.410000 ;
      RECT 1066.500000 283.590000 1108.500000 284.410000 ;
      RECT 1016.500000 283.590000 1058.500000 284.410000 ;
      RECT 966.500000 283.590000 1008.500000 284.410000 ;
      RECT 916.500000 283.590000 958.500000 284.410000 ;
      RECT 866.500000 283.590000 908.500000 284.410000 ;
      RECT 816.500000 283.590000 858.500000 284.410000 ;
      RECT 766.500000 283.590000 808.500000 284.410000 ;
      RECT 716.500000 283.590000 758.500000 284.410000 ;
      RECT 666.500000 283.590000 708.500000 284.410000 ;
      RECT 616.500000 283.590000 658.500000 284.410000 ;
      RECT 566.500000 283.590000 608.500000 284.410000 ;
      RECT 516.500000 283.590000 558.500000 284.410000 ;
      RECT 466.500000 283.590000 508.500000 284.410000 ;
      RECT 416.500000 283.590000 458.500000 284.410000 ;
      RECT 366.500000 283.590000 408.500000 284.410000 ;
      RECT 316.500000 283.590000 358.500000 284.410000 ;
      RECT 266.500000 283.590000 308.500000 284.410000 ;
      RECT 216.500000 283.590000 258.500000 284.410000 ;
      RECT 166.500000 283.590000 208.500000 284.410000 ;
      RECT 116.500000 283.590000 158.500000 284.410000 ;
      RECT 66.500000 283.590000 108.500000 284.410000 ;
      RECT 29.500000 283.590000 58.500000 284.410000 ;
      RECT 0.000000 283.590000 16.500000 284.410000 ;
      RECT 1169.500000 282.410000 1170.500000 283.590000 ;
      RECT 1116.500000 282.410000 1149.500000 283.590000 ;
      RECT 1107.500000 282.410000 1108.500000 283.590000 ;
      RECT 1066.500000 282.410000 1099.500000 283.590000 ;
      RECT 1057.500000 282.410000 1058.500000 283.590000 ;
      RECT 1016.500000 282.410000 1049.500000 283.590000 ;
      RECT 1007.500000 282.410000 1008.500000 283.590000 ;
      RECT 966.500000 282.410000 999.500000 283.590000 ;
      RECT 957.500000 282.410000 958.500000 283.590000 ;
      RECT 916.500000 282.410000 949.500000 283.590000 ;
      RECT 907.500000 282.410000 908.500000 283.590000 ;
      RECT 866.500000 282.410000 899.500000 283.590000 ;
      RECT 857.500000 282.410000 858.500000 283.590000 ;
      RECT 816.500000 282.410000 849.500000 283.590000 ;
      RECT 807.500000 282.410000 808.500000 283.590000 ;
      RECT 766.500000 282.410000 799.500000 283.590000 ;
      RECT 757.500000 282.410000 758.500000 283.590000 ;
      RECT 716.500000 282.410000 749.500000 283.590000 ;
      RECT 707.500000 282.410000 708.500000 283.590000 ;
      RECT 666.500000 282.410000 699.500000 283.590000 ;
      RECT 657.500000 282.410000 658.500000 283.590000 ;
      RECT 616.500000 282.410000 649.500000 283.590000 ;
      RECT 607.500000 282.410000 608.500000 283.590000 ;
      RECT 566.500000 282.410000 599.500000 283.590000 ;
      RECT 557.500000 282.410000 558.500000 283.590000 ;
      RECT 516.500000 282.410000 549.500000 283.590000 ;
      RECT 507.500000 282.410000 508.500000 283.590000 ;
      RECT 466.500000 282.410000 499.500000 283.590000 ;
      RECT 457.500000 282.410000 458.500000 283.590000 ;
      RECT 416.500000 282.410000 449.500000 283.590000 ;
      RECT 407.500000 282.410000 408.500000 283.590000 ;
      RECT 366.500000 282.410000 399.500000 283.590000 ;
      RECT 357.500000 282.410000 358.500000 283.590000 ;
      RECT 316.500000 282.410000 349.500000 283.590000 ;
      RECT 307.500000 282.410000 308.500000 283.590000 ;
      RECT 266.500000 282.410000 299.500000 283.590000 ;
      RECT 257.500000 282.410000 258.500000 283.590000 ;
      RECT 216.500000 282.410000 249.500000 283.590000 ;
      RECT 207.500000 282.410000 208.500000 283.590000 ;
      RECT 166.500000 282.410000 199.500000 283.590000 ;
      RECT 157.500000 282.410000 158.500000 283.590000 ;
      RECT 116.500000 282.410000 149.500000 283.590000 ;
      RECT 107.500000 282.410000 108.500000 283.590000 ;
      RECT 66.500000 282.410000 99.500000 283.590000 ;
      RECT 57.500000 282.410000 58.500000 283.590000 ;
      RECT 29.500000 282.410000 49.500000 283.590000 ;
      RECT 15.500000 282.410000 16.500000 283.590000 ;
      RECT 1157.500000 281.590000 1170.500000 282.410000 ;
      RECT 1107.500000 281.590000 1149.500000 282.410000 ;
      RECT 1057.500000 281.590000 1099.500000 282.410000 ;
      RECT 1007.500000 281.590000 1049.500000 282.410000 ;
      RECT 957.500000 281.590000 999.500000 282.410000 ;
      RECT 907.500000 281.590000 949.500000 282.410000 ;
      RECT 857.500000 281.590000 899.500000 282.410000 ;
      RECT 807.500000 281.590000 849.500000 282.410000 ;
      RECT 757.500000 281.590000 799.500000 282.410000 ;
      RECT 707.500000 281.590000 749.500000 282.410000 ;
      RECT 657.500000 281.590000 699.500000 282.410000 ;
      RECT 607.500000 281.590000 649.500000 282.410000 ;
      RECT 557.500000 281.590000 599.500000 282.410000 ;
      RECT 507.500000 281.590000 549.500000 282.410000 ;
      RECT 457.500000 281.590000 499.500000 282.410000 ;
      RECT 407.500000 281.590000 449.500000 282.410000 ;
      RECT 357.500000 281.590000 399.500000 282.410000 ;
      RECT 307.500000 281.590000 349.500000 282.410000 ;
      RECT 257.500000 281.590000 299.500000 282.410000 ;
      RECT 207.500000 281.590000 249.500000 282.410000 ;
      RECT 157.500000 281.590000 199.500000 282.410000 ;
      RECT 107.500000 281.590000 149.500000 282.410000 ;
      RECT 57.500000 281.590000 99.500000 282.410000 ;
      RECT 15.500000 281.590000 49.500000 282.410000 ;
      RECT 1183.500000 280.410000 1186.000000 283.590000 ;
      RECT 1169.500000 280.410000 1170.500000 281.590000 ;
      RECT 1116.500000 280.410000 1149.500000 281.590000 ;
      RECT 1107.500000 280.410000 1108.500000 281.590000 ;
      RECT 1066.500000 280.410000 1099.500000 281.590000 ;
      RECT 1057.500000 280.410000 1058.500000 281.590000 ;
      RECT 1016.500000 280.410000 1049.500000 281.590000 ;
      RECT 1007.500000 280.410000 1008.500000 281.590000 ;
      RECT 966.500000 280.410000 999.500000 281.590000 ;
      RECT 957.500000 280.410000 958.500000 281.590000 ;
      RECT 916.500000 280.410000 949.500000 281.590000 ;
      RECT 907.500000 280.410000 908.500000 281.590000 ;
      RECT 866.500000 280.410000 899.500000 281.590000 ;
      RECT 857.500000 280.410000 858.500000 281.590000 ;
      RECT 816.500000 280.410000 849.500000 281.590000 ;
      RECT 807.500000 280.410000 808.500000 281.590000 ;
      RECT 766.500000 280.410000 799.500000 281.590000 ;
      RECT 757.500000 280.410000 758.500000 281.590000 ;
      RECT 716.500000 280.410000 749.500000 281.590000 ;
      RECT 707.500000 280.410000 708.500000 281.590000 ;
      RECT 666.500000 280.410000 699.500000 281.590000 ;
      RECT 657.500000 280.410000 658.500000 281.590000 ;
      RECT 616.500000 280.410000 649.500000 281.590000 ;
      RECT 607.500000 280.410000 608.500000 281.590000 ;
      RECT 566.500000 280.410000 599.500000 281.590000 ;
      RECT 557.500000 280.410000 558.500000 281.590000 ;
      RECT 516.500000 280.410000 549.500000 281.590000 ;
      RECT 507.500000 280.410000 508.500000 281.590000 ;
      RECT 466.500000 280.410000 499.500000 281.590000 ;
      RECT 457.500000 280.410000 458.500000 281.590000 ;
      RECT 416.500000 280.410000 449.500000 281.590000 ;
      RECT 407.500000 280.410000 408.500000 281.590000 ;
      RECT 366.500000 280.410000 399.500000 281.590000 ;
      RECT 357.500000 280.410000 358.500000 281.590000 ;
      RECT 316.500000 280.410000 349.500000 281.590000 ;
      RECT 307.500000 280.410000 308.500000 281.590000 ;
      RECT 266.500000 280.410000 299.500000 281.590000 ;
      RECT 257.500000 280.410000 258.500000 281.590000 ;
      RECT 216.500000 280.410000 249.500000 281.590000 ;
      RECT 207.500000 280.410000 208.500000 281.590000 ;
      RECT 166.500000 280.410000 199.500000 281.590000 ;
      RECT 157.500000 280.410000 158.500000 281.590000 ;
      RECT 116.500000 280.410000 149.500000 281.590000 ;
      RECT 107.500000 280.410000 108.500000 281.590000 ;
      RECT 66.500000 280.410000 99.500000 281.590000 ;
      RECT 57.500000 280.410000 58.500000 281.590000 ;
      RECT 29.500000 280.410000 49.500000 281.590000 ;
      RECT 15.500000 280.410000 16.500000 281.590000 ;
      RECT 0.000000 280.410000 2.500000 283.590000 ;
      RECT 1169.500000 279.590000 1186.000000 280.410000 ;
      RECT 1116.500000 279.590000 1156.500000 280.410000 ;
      RECT 1066.500000 279.590000 1108.500000 280.410000 ;
      RECT 1016.500000 279.590000 1058.500000 280.410000 ;
      RECT 966.500000 279.590000 1008.500000 280.410000 ;
      RECT 916.500000 279.590000 958.500000 280.410000 ;
      RECT 866.500000 279.590000 908.500000 280.410000 ;
      RECT 816.500000 279.590000 858.500000 280.410000 ;
      RECT 766.500000 279.590000 808.500000 280.410000 ;
      RECT 716.500000 279.590000 758.500000 280.410000 ;
      RECT 666.500000 279.590000 708.500000 280.410000 ;
      RECT 616.500000 279.590000 658.500000 280.410000 ;
      RECT 566.500000 279.590000 608.500000 280.410000 ;
      RECT 516.500000 279.590000 558.500000 280.410000 ;
      RECT 466.500000 279.590000 508.500000 280.410000 ;
      RECT 416.500000 279.590000 458.500000 280.410000 ;
      RECT 366.500000 279.590000 408.500000 280.410000 ;
      RECT 316.500000 279.590000 358.500000 280.410000 ;
      RECT 266.500000 279.590000 308.500000 280.410000 ;
      RECT 216.500000 279.590000 258.500000 280.410000 ;
      RECT 166.500000 279.590000 208.500000 280.410000 ;
      RECT 116.500000 279.590000 158.500000 280.410000 ;
      RECT 66.500000 279.590000 108.500000 280.410000 ;
      RECT 29.500000 279.590000 58.500000 280.410000 ;
      RECT 0.000000 279.590000 16.500000 280.410000 ;
      RECT 1169.500000 278.410000 1170.500000 279.590000 ;
      RECT 1116.500000 278.410000 1149.500000 279.590000 ;
      RECT 1107.500000 278.410000 1108.500000 279.590000 ;
      RECT 1066.500000 278.410000 1099.500000 279.590000 ;
      RECT 1057.500000 278.410000 1058.500000 279.590000 ;
      RECT 1016.500000 278.410000 1049.500000 279.590000 ;
      RECT 1007.500000 278.410000 1008.500000 279.590000 ;
      RECT 966.500000 278.410000 999.500000 279.590000 ;
      RECT 957.500000 278.410000 958.500000 279.590000 ;
      RECT 916.500000 278.410000 949.500000 279.590000 ;
      RECT 907.500000 278.410000 908.500000 279.590000 ;
      RECT 866.500000 278.410000 899.500000 279.590000 ;
      RECT 857.500000 278.410000 858.500000 279.590000 ;
      RECT 816.500000 278.410000 849.500000 279.590000 ;
      RECT 807.500000 278.410000 808.500000 279.590000 ;
      RECT 766.500000 278.410000 799.500000 279.590000 ;
      RECT 757.500000 278.410000 758.500000 279.590000 ;
      RECT 716.500000 278.410000 749.500000 279.590000 ;
      RECT 707.500000 278.410000 708.500000 279.590000 ;
      RECT 666.500000 278.410000 699.500000 279.590000 ;
      RECT 657.500000 278.410000 658.500000 279.590000 ;
      RECT 616.500000 278.410000 649.500000 279.590000 ;
      RECT 607.500000 278.410000 608.500000 279.590000 ;
      RECT 566.500000 278.410000 599.500000 279.590000 ;
      RECT 557.500000 278.410000 558.500000 279.590000 ;
      RECT 516.500000 278.410000 549.500000 279.590000 ;
      RECT 507.500000 278.410000 508.500000 279.590000 ;
      RECT 466.500000 278.410000 499.500000 279.590000 ;
      RECT 457.500000 278.410000 458.500000 279.590000 ;
      RECT 416.500000 278.410000 449.500000 279.590000 ;
      RECT 407.500000 278.410000 408.500000 279.590000 ;
      RECT 366.500000 278.410000 399.500000 279.590000 ;
      RECT 357.500000 278.410000 358.500000 279.590000 ;
      RECT 316.500000 278.410000 349.500000 279.590000 ;
      RECT 307.500000 278.410000 308.500000 279.590000 ;
      RECT 266.500000 278.410000 299.500000 279.590000 ;
      RECT 257.500000 278.410000 258.500000 279.590000 ;
      RECT 216.500000 278.410000 249.500000 279.590000 ;
      RECT 207.500000 278.410000 208.500000 279.590000 ;
      RECT 166.500000 278.410000 199.500000 279.590000 ;
      RECT 157.500000 278.410000 158.500000 279.590000 ;
      RECT 116.500000 278.410000 149.500000 279.590000 ;
      RECT 107.500000 278.410000 108.500000 279.590000 ;
      RECT 66.500000 278.410000 99.500000 279.590000 ;
      RECT 57.500000 278.410000 58.500000 279.590000 ;
      RECT 29.500000 278.410000 49.500000 279.590000 ;
      RECT 15.500000 278.410000 16.500000 279.590000 ;
      RECT 1157.500000 277.590000 1170.500000 278.410000 ;
      RECT 1107.500000 277.590000 1149.500000 278.410000 ;
      RECT 1057.500000 277.590000 1099.500000 278.410000 ;
      RECT 1007.500000 277.590000 1049.500000 278.410000 ;
      RECT 957.500000 277.590000 999.500000 278.410000 ;
      RECT 907.500000 277.590000 949.500000 278.410000 ;
      RECT 857.500000 277.590000 899.500000 278.410000 ;
      RECT 807.500000 277.590000 849.500000 278.410000 ;
      RECT 757.500000 277.590000 799.500000 278.410000 ;
      RECT 707.500000 277.590000 749.500000 278.410000 ;
      RECT 657.500000 277.590000 699.500000 278.410000 ;
      RECT 607.500000 277.590000 649.500000 278.410000 ;
      RECT 557.500000 277.590000 599.500000 278.410000 ;
      RECT 507.500000 277.590000 549.500000 278.410000 ;
      RECT 457.500000 277.590000 499.500000 278.410000 ;
      RECT 407.500000 277.590000 449.500000 278.410000 ;
      RECT 357.500000 277.590000 399.500000 278.410000 ;
      RECT 307.500000 277.590000 349.500000 278.410000 ;
      RECT 257.500000 277.590000 299.500000 278.410000 ;
      RECT 207.500000 277.590000 249.500000 278.410000 ;
      RECT 157.500000 277.590000 199.500000 278.410000 ;
      RECT 107.500000 277.590000 149.500000 278.410000 ;
      RECT 57.500000 277.590000 99.500000 278.410000 ;
      RECT 15.500000 277.590000 49.500000 278.410000 ;
      RECT 1183.500000 276.410000 1186.000000 279.590000 ;
      RECT 1169.500000 276.410000 1170.500000 277.590000 ;
      RECT 1116.500000 276.410000 1149.500000 277.590000 ;
      RECT 1107.500000 276.410000 1108.500000 277.590000 ;
      RECT 1066.500000 276.410000 1099.500000 277.590000 ;
      RECT 1057.500000 276.410000 1058.500000 277.590000 ;
      RECT 1016.500000 276.410000 1049.500000 277.590000 ;
      RECT 1007.500000 276.410000 1008.500000 277.590000 ;
      RECT 966.500000 276.410000 999.500000 277.590000 ;
      RECT 957.500000 276.410000 958.500000 277.590000 ;
      RECT 916.500000 276.410000 949.500000 277.590000 ;
      RECT 907.500000 276.410000 908.500000 277.590000 ;
      RECT 866.500000 276.410000 899.500000 277.590000 ;
      RECT 857.500000 276.410000 858.500000 277.590000 ;
      RECT 816.500000 276.410000 849.500000 277.590000 ;
      RECT 807.500000 276.410000 808.500000 277.590000 ;
      RECT 766.500000 276.410000 799.500000 277.590000 ;
      RECT 757.500000 276.410000 758.500000 277.590000 ;
      RECT 716.500000 276.410000 749.500000 277.590000 ;
      RECT 707.500000 276.410000 708.500000 277.590000 ;
      RECT 666.500000 276.410000 699.500000 277.590000 ;
      RECT 657.500000 276.410000 658.500000 277.590000 ;
      RECT 616.500000 276.410000 649.500000 277.590000 ;
      RECT 607.500000 276.410000 608.500000 277.590000 ;
      RECT 566.500000 276.410000 599.500000 277.590000 ;
      RECT 557.500000 276.410000 558.500000 277.590000 ;
      RECT 516.500000 276.410000 549.500000 277.590000 ;
      RECT 507.500000 276.410000 508.500000 277.590000 ;
      RECT 466.500000 276.410000 499.500000 277.590000 ;
      RECT 457.500000 276.410000 458.500000 277.590000 ;
      RECT 416.500000 276.410000 449.500000 277.590000 ;
      RECT 407.500000 276.410000 408.500000 277.590000 ;
      RECT 366.500000 276.410000 399.500000 277.590000 ;
      RECT 357.500000 276.410000 358.500000 277.590000 ;
      RECT 316.500000 276.410000 349.500000 277.590000 ;
      RECT 307.500000 276.410000 308.500000 277.590000 ;
      RECT 266.500000 276.410000 299.500000 277.590000 ;
      RECT 257.500000 276.410000 258.500000 277.590000 ;
      RECT 216.500000 276.410000 249.500000 277.590000 ;
      RECT 207.500000 276.410000 208.500000 277.590000 ;
      RECT 166.500000 276.410000 199.500000 277.590000 ;
      RECT 157.500000 276.410000 158.500000 277.590000 ;
      RECT 116.500000 276.410000 149.500000 277.590000 ;
      RECT 107.500000 276.410000 108.500000 277.590000 ;
      RECT 66.500000 276.410000 99.500000 277.590000 ;
      RECT 57.500000 276.410000 58.500000 277.590000 ;
      RECT 29.500000 276.410000 49.500000 277.590000 ;
      RECT 15.500000 276.410000 16.500000 277.590000 ;
      RECT 0.000000 276.410000 2.500000 279.590000 ;
      RECT 1169.500000 275.590000 1186.000000 276.410000 ;
      RECT 1116.500000 275.590000 1156.500000 276.410000 ;
      RECT 1066.500000 275.590000 1108.500000 276.410000 ;
      RECT 1016.500000 275.590000 1058.500000 276.410000 ;
      RECT 966.500000 275.590000 1008.500000 276.410000 ;
      RECT 916.500000 275.590000 958.500000 276.410000 ;
      RECT 866.500000 275.590000 908.500000 276.410000 ;
      RECT 816.500000 275.590000 858.500000 276.410000 ;
      RECT 766.500000 275.590000 808.500000 276.410000 ;
      RECT 716.500000 275.590000 758.500000 276.410000 ;
      RECT 666.500000 275.590000 708.500000 276.410000 ;
      RECT 616.500000 275.590000 658.500000 276.410000 ;
      RECT 566.500000 275.590000 608.500000 276.410000 ;
      RECT 516.500000 275.590000 558.500000 276.410000 ;
      RECT 466.500000 275.590000 508.500000 276.410000 ;
      RECT 416.500000 275.590000 458.500000 276.410000 ;
      RECT 366.500000 275.590000 408.500000 276.410000 ;
      RECT 316.500000 275.590000 358.500000 276.410000 ;
      RECT 266.500000 275.590000 308.500000 276.410000 ;
      RECT 216.500000 275.590000 258.500000 276.410000 ;
      RECT 166.500000 275.590000 208.500000 276.410000 ;
      RECT 116.500000 275.590000 158.500000 276.410000 ;
      RECT 66.500000 275.590000 108.500000 276.410000 ;
      RECT 29.500000 275.590000 58.500000 276.410000 ;
      RECT 0.000000 275.590000 16.500000 276.410000 ;
      RECT 1169.500000 274.410000 1170.500000 275.590000 ;
      RECT 1116.500000 274.410000 1149.500000 275.590000 ;
      RECT 1107.500000 274.410000 1108.500000 275.590000 ;
      RECT 1066.500000 274.410000 1099.500000 275.590000 ;
      RECT 1057.500000 274.410000 1058.500000 275.590000 ;
      RECT 1016.500000 274.410000 1049.500000 275.590000 ;
      RECT 1007.500000 274.410000 1008.500000 275.590000 ;
      RECT 966.500000 274.410000 999.500000 275.590000 ;
      RECT 957.500000 274.410000 958.500000 275.590000 ;
      RECT 916.500000 274.410000 949.500000 275.590000 ;
      RECT 907.500000 274.410000 908.500000 275.590000 ;
      RECT 866.500000 274.410000 899.500000 275.590000 ;
      RECT 857.500000 274.410000 858.500000 275.590000 ;
      RECT 816.500000 274.410000 849.500000 275.590000 ;
      RECT 807.500000 274.410000 808.500000 275.590000 ;
      RECT 766.500000 274.410000 799.500000 275.590000 ;
      RECT 757.500000 274.410000 758.500000 275.590000 ;
      RECT 716.500000 274.410000 749.500000 275.590000 ;
      RECT 707.500000 274.410000 708.500000 275.590000 ;
      RECT 666.500000 274.410000 699.500000 275.590000 ;
      RECT 657.500000 274.410000 658.500000 275.590000 ;
      RECT 616.500000 274.410000 649.500000 275.590000 ;
      RECT 607.500000 274.410000 608.500000 275.590000 ;
      RECT 566.500000 274.410000 599.500000 275.590000 ;
      RECT 557.500000 274.410000 558.500000 275.590000 ;
      RECT 516.500000 274.410000 549.500000 275.590000 ;
      RECT 507.500000 274.410000 508.500000 275.590000 ;
      RECT 466.500000 274.410000 499.500000 275.590000 ;
      RECT 457.500000 274.410000 458.500000 275.590000 ;
      RECT 416.500000 274.410000 449.500000 275.590000 ;
      RECT 407.500000 274.410000 408.500000 275.590000 ;
      RECT 366.500000 274.410000 399.500000 275.590000 ;
      RECT 357.500000 274.410000 358.500000 275.590000 ;
      RECT 316.500000 274.410000 349.500000 275.590000 ;
      RECT 307.500000 274.410000 308.500000 275.590000 ;
      RECT 266.500000 274.410000 299.500000 275.590000 ;
      RECT 257.500000 274.410000 258.500000 275.590000 ;
      RECT 216.500000 274.410000 249.500000 275.590000 ;
      RECT 207.500000 274.410000 208.500000 275.590000 ;
      RECT 166.500000 274.410000 199.500000 275.590000 ;
      RECT 157.500000 274.410000 158.500000 275.590000 ;
      RECT 116.500000 274.410000 149.500000 275.590000 ;
      RECT 107.500000 274.410000 108.500000 275.590000 ;
      RECT 66.500000 274.410000 99.500000 275.590000 ;
      RECT 57.500000 274.410000 58.500000 275.590000 ;
      RECT 29.500000 274.410000 49.500000 275.590000 ;
      RECT 15.500000 274.410000 16.500000 275.590000 ;
      RECT 1157.500000 273.590000 1170.500000 274.410000 ;
      RECT 1107.500000 273.590000 1149.500000 274.410000 ;
      RECT 1057.500000 273.590000 1099.500000 274.410000 ;
      RECT 1007.500000 273.590000 1049.500000 274.410000 ;
      RECT 957.500000 273.590000 999.500000 274.410000 ;
      RECT 907.500000 273.590000 949.500000 274.410000 ;
      RECT 857.500000 273.590000 899.500000 274.410000 ;
      RECT 807.500000 273.590000 849.500000 274.410000 ;
      RECT 757.500000 273.590000 799.500000 274.410000 ;
      RECT 707.500000 273.590000 749.500000 274.410000 ;
      RECT 657.500000 273.590000 699.500000 274.410000 ;
      RECT 607.500000 273.590000 649.500000 274.410000 ;
      RECT 557.500000 273.590000 599.500000 274.410000 ;
      RECT 507.500000 273.590000 549.500000 274.410000 ;
      RECT 457.500000 273.590000 499.500000 274.410000 ;
      RECT 407.500000 273.590000 449.500000 274.410000 ;
      RECT 357.500000 273.590000 399.500000 274.410000 ;
      RECT 307.500000 273.590000 349.500000 274.410000 ;
      RECT 257.500000 273.590000 299.500000 274.410000 ;
      RECT 207.500000 273.590000 249.500000 274.410000 ;
      RECT 157.500000 273.590000 199.500000 274.410000 ;
      RECT 107.500000 273.590000 149.500000 274.410000 ;
      RECT 57.500000 273.590000 99.500000 274.410000 ;
      RECT 15.500000 273.590000 49.500000 274.410000 ;
      RECT 1183.500000 272.410000 1186.000000 275.590000 ;
      RECT 1169.500000 272.410000 1170.500000 273.590000 ;
      RECT 1116.500000 272.410000 1149.500000 273.590000 ;
      RECT 1107.500000 272.410000 1108.500000 273.590000 ;
      RECT 1066.500000 272.410000 1099.500000 273.590000 ;
      RECT 1057.500000 272.410000 1058.500000 273.590000 ;
      RECT 1016.500000 272.410000 1049.500000 273.590000 ;
      RECT 1007.500000 272.410000 1008.500000 273.590000 ;
      RECT 966.500000 272.410000 999.500000 273.590000 ;
      RECT 957.500000 272.410000 958.500000 273.590000 ;
      RECT 916.500000 272.410000 949.500000 273.590000 ;
      RECT 907.500000 272.410000 908.500000 273.590000 ;
      RECT 866.500000 272.410000 899.500000 273.590000 ;
      RECT 857.500000 272.410000 858.500000 273.590000 ;
      RECT 816.500000 272.410000 849.500000 273.590000 ;
      RECT 807.500000 272.410000 808.500000 273.590000 ;
      RECT 766.500000 272.410000 799.500000 273.590000 ;
      RECT 757.500000 272.410000 758.500000 273.590000 ;
      RECT 716.500000 272.410000 749.500000 273.590000 ;
      RECT 707.500000 272.410000 708.500000 273.590000 ;
      RECT 666.500000 272.410000 699.500000 273.590000 ;
      RECT 657.500000 272.410000 658.500000 273.590000 ;
      RECT 616.500000 272.410000 649.500000 273.590000 ;
      RECT 607.500000 272.410000 608.500000 273.590000 ;
      RECT 566.500000 272.410000 599.500000 273.590000 ;
      RECT 557.500000 272.410000 558.500000 273.590000 ;
      RECT 516.500000 272.410000 549.500000 273.590000 ;
      RECT 507.500000 272.410000 508.500000 273.590000 ;
      RECT 466.500000 272.410000 499.500000 273.590000 ;
      RECT 457.500000 272.410000 458.500000 273.590000 ;
      RECT 416.500000 272.410000 449.500000 273.590000 ;
      RECT 407.500000 272.410000 408.500000 273.590000 ;
      RECT 366.500000 272.410000 399.500000 273.590000 ;
      RECT 357.500000 272.410000 358.500000 273.590000 ;
      RECT 316.500000 272.410000 349.500000 273.590000 ;
      RECT 307.500000 272.410000 308.500000 273.590000 ;
      RECT 266.500000 272.410000 299.500000 273.590000 ;
      RECT 257.500000 272.410000 258.500000 273.590000 ;
      RECT 216.500000 272.410000 249.500000 273.590000 ;
      RECT 207.500000 272.410000 208.500000 273.590000 ;
      RECT 166.500000 272.410000 199.500000 273.590000 ;
      RECT 157.500000 272.410000 158.500000 273.590000 ;
      RECT 116.500000 272.410000 149.500000 273.590000 ;
      RECT 107.500000 272.410000 108.500000 273.590000 ;
      RECT 66.500000 272.410000 99.500000 273.590000 ;
      RECT 57.500000 272.410000 58.500000 273.590000 ;
      RECT 29.500000 272.410000 49.500000 273.590000 ;
      RECT 15.500000 272.410000 16.500000 273.590000 ;
      RECT 0.000000 272.410000 2.500000 275.590000 ;
      RECT 1169.500000 271.590000 1186.000000 272.410000 ;
      RECT 1116.500000 271.590000 1156.500000 272.410000 ;
      RECT 1066.500000 271.590000 1108.500000 272.410000 ;
      RECT 1016.500000 271.590000 1058.500000 272.410000 ;
      RECT 966.500000 271.590000 1008.500000 272.410000 ;
      RECT 916.500000 271.590000 958.500000 272.410000 ;
      RECT 866.500000 271.590000 908.500000 272.410000 ;
      RECT 816.500000 271.590000 858.500000 272.410000 ;
      RECT 766.500000 271.590000 808.500000 272.410000 ;
      RECT 716.500000 271.590000 758.500000 272.410000 ;
      RECT 666.500000 271.590000 708.500000 272.410000 ;
      RECT 616.500000 271.590000 658.500000 272.410000 ;
      RECT 566.500000 271.590000 608.500000 272.410000 ;
      RECT 516.500000 271.590000 558.500000 272.410000 ;
      RECT 466.500000 271.590000 508.500000 272.410000 ;
      RECT 416.500000 271.590000 458.500000 272.410000 ;
      RECT 366.500000 271.590000 408.500000 272.410000 ;
      RECT 316.500000 271.590000 358.500000 272.410000 ;
      RECT 266.500000 271.590000 308.500000 272.410000 ;
      RECT 216.500000 271.590000 258.500000 272.410000 ;
      RECT 166.500000 271.590000 208.500000 272.410000 ;
      RECT 116.500000 271.590000 158.500000 272.410000 ;
      RECT 66.500000 271.590000 108.500000 272.410000 ;
      RECT 29.500000 271.590000 58.500000 272.410000 ;
      RECT 0.000000 271.590000 16.500000 272.410000 ;
      RECT 1169.500000 270.410000 1170.500000 271.590000 ;
      RECT 1116.500000 270.410000 1149.500000 271.590000 ;
      RECT 1107.500000 270.410000 1108.500000 271.590000 ;
      RECT 1066.500000 270.410000 1099.500000 271.590000 ;
      RECT 1057.500000 270.410000 1058.500000 271.590000 ;
      RECT 1016.500000 270.410000 1049.500000 271.590000 ;
      RECT 1007.500000 270.410000 1008.500000 271.590000 ;
      RECT 966.500000 270.410000 999.500000 271.590000 ;
      RECT 957.500000 270.410000 958.500000 271.590000 ;
      RECT 916.500000 270.410000 949.500000 271.590000 ;
      RECT 907.500000 270.410000 908.500000 271.590000 ;
      RECT 866.500000 270.410000 899.500000 271.590000 ;
      RECT 857.500000 270.410000 858.500000 271.590000 ;
      RECT 816.500000 270.410000 849.500000 271.590000 ;
      RECT 807.500000 270.410000 808.500000 271.590000 ;
      RECT 766.500000 270.410000 799.500000 271.590000 ;
      RECT 757.500000 270.410000 758.500000 271.590000 ;
      RECT 716.500000 270.410000 749.500000 271.590000 ;
      RECT 707.500000 270.410000 708.500000 271.590000 ;
      RECT 666.500000 270.410000 699.500000 271.590000 ;
      RECT 657.500000 270.410000 658.500000 271.590000 ;
      RECT 616.500000 270.410000 649.500000 271.590000 ;
      RECT 607.500000 270.410000 608.500000 271.590000 ;
      RECT 566.500000 270.410000 599.500000 271.590000 ;
      RECT 557.500000 270.410000 558.500000 271.590000 ;
      RECT 516.500000 270.410000 549.500000 271.590000 ;
      RECT 507.500000 270.410000 508.500000 271.590000 ;
      RECT 466.500000 270.410000 499.500000 271.590000 ;
      RECT 457.500000 270.410000 458.500000 271.590000 ;
      RECT 416.500000 270.410000 449.500000 271.590000 ;
      RECT 407.500000 270.410000 408.500000 271.590000 ;
      RECT 366.500000 270.410000 399.500000 271.590000 ;
      RECT 357.500000 270.410000 358.500000 271.590000 ;
      RECT 316.500000 270.410000 349.500000 271.590000 ;
      RECT 307.500000 270.410000 308.500000 271.590000 ;
      RECT 266.500000 270.410000 299.500000 271.590000 ;
      RECT 257.500000 270.410000 258.500000 271.590000 ;
      RECT 216.500000 270.410000 249.500000 271.590000 ;
      RECT 207.500000 270.410000 208.500000 271.590000 ;
      RECT 166.500000 270.410000 199.500000 271.590000 ;
      RECT 157.500000 270.410000 158.500000 271.590000 ;
      RECT 116.500000 270.410000 149.500000 271.590000 ;
      RECT 107.500000 270.410000 108.500000 271.590000 ;
      RECT 66.500000 270.410000 99.500000 271.590000 ;
      RECT 57.500000 270.410000 58.500000 271.590000 ;
      RECT 29.500000 270.410000 49.500000 271.590000 ;
      RECT 15.500000 270.410000 16.500000 271.590000 ;
      RECT 1157.500000 269.590000 1170.500000 270.410000 ;
      RECT 1107.500000 269.590000 1149.500000 270.410000 ;
      RECT 1057.500000 269.590000 1099.500000 270.410000 ;
      RECT 1007.500000 269.590000 1049.500000 270.410000 ;
      RECT 957.500000 269.590000 999.500000 270.410000 ;
      RECT 907.500000 269.590000 949.500000 270.410000 ;
      RECT 857.500000 269.590000 899.500000 270.410000 ;
      RECT 807.500000 269.590000 849.500000 270.410000 ;
      RECT 757.500000 269.590000 799.500000 270.410000 ;
      RECT 707.500000 269.590000 749.500000 270.410000 ;
      RECT 657.500000 269.590000 699.500000 270.410000 ;
      RECT 607.500000 269.590000 649.500000 270.410000 ;
      RECT 557.500000 269.590000 599.500000 270.410000 ;
      RECT 507.500000 269.590000 549.500000 270.410000 ;
      RECT 457.500000 269.590000 499.500000 270.410000 ;
      RECT 407.500000 269.590000 449.500000 270.410000 ;
      RECT 357.500000 269.590000 399.500000 270.410000 ;
      RECT 307.500000 269.590000 349.500000 270.410000 ;
      RECT 257.500000 269.590000 299.500000 270.410000 ;
      RECT 207.500000 269.590000 249.500000 270.410000 ;
      RECT 157.500000 269.590000 199.500000 270.410000 ;
      RECT 107.500000 269.590000 149.500000 270.410000 ;
      RECT 57.500000 269.590000 99.500000 270.410000 ;
      RECT 15.500000 269.590000 49.500000 270.410000 ;
      RECT 1183.500000 268.410000 1186.000000 271.590000 ;
      RECT 1169.500000 268.410000 1170.500000 269.590000 ;
      RECT 1116.500000 268.410000 1149.500000 269.590000 ;
      RECT 1107.500000 268.410000 1108.500000 269.590000 ;
      RECT 1066.500000 268.410000 1099.500000 269.590000 ;
      RECT 1057.500000 268.410000 1058.500000 269.590000 ;
      RECT 1016.500000 268.410000 1049.500000 269.590000 ;
      RECT 1007.500000 268.410000 1008.500000 269.590000 ;
      RECT 966.500000 268.410000 999.500000 269.590000 ;
      RECT 957.500000 268.410000 958.500000 269.590000 ;
      RECT 916.500000 268.410000 949.500000 269.590000 ;
      RECT 907.500000 268.410000 908.500000 269.590000 ;
      RECT 866.500000 268.410000 899.500000 269.590000 ;
      RECT 857.500000 268.410000 858.500000 269.590000 ;
      RECT 816.500000 268.410000 849.500000 269.590000 ;
      RECT 807.500000 268.410000 808.500000 269.590000 ;
      RECT 766.500000 268.410000 799.500000 269.590000 ;
      RECT 757.500000 268.410000 758.500000 269.590000 ;
      RECT 716.500000 268.410000 749.500000 269.590000 ;
      RECT 707.500000 268.410000 708.500000 269.590000 ;
      RECT 666.500000 268.410000 699.500000 269.590000 ;
      RECT 657.500000 268.410000 658.500000 269.590000 ;
      RECT 616.500000 268.410000 649.500000 269.590000 ;
      RECT 607.500000 268.410000 608.500000 269.590000 ;
      RECT 566.500000 268.410000 599.500000 269.590000 ;
      RECT 557.500000 268.410000 558.500000 269.590000 ;
      RECT 516.500000 268.410000 549.500000 269.590000 ;
      RECT 507.500000 268.410000 508.500000 269.590000 ;
      RECT 466.500000 268.410000 499.500000 269.590000 ;
      RECT 457.500000 268.410000 458.500000 269.590000 ;
      RECT 416.500000 268.410000 449.500000 269.590000 ;
      RECT 407.500000 268.410000 408.500000 269.590000 ;
      RECT 366.500000 268.410000 399.500000 269.590000 ;
      RECT 357.500000 268.410000 358.500000 269.590000 ;
      RECT 316.500000 268.410000 349.500000 269.590000 ;
      RECT 307.500000 268.410000 308.500000 269.590000 ;
      RECT 266.500000 268.410000 299.500000 269.590000 ;
      RECT 257.500000 268.410000 258.500000 269.590000 ;
      RECT 216.500000 268.410000 249.500000 269.590000 ;
      RECT 207.500000 268.410000 208.500000 269.590000 ;
      RECT 166.500000 268.410000 199.500000 269.590000 ;
      RECT 157.500000 268.410000 158.500000 269.590000 ;
      RECT 116.500000 268.410000 149.500000 269.590000 ;
      RECT 107.500000 268.410000 108.500000 269.590000 ;
      RECT 66.500000 268.410000 99.500000 269.590000 ;
      RECT 57.500000 268.410000 58.500000 269.590000 ;
      RECT 29.500000 268.410000 49.500000 269.590000 ;
      RECT 15.500000 268.410000 16.500000 269.590000 ;
      RECT 0.000000 268.410000 2.500000 271.590000 ;
      RECT 1169.500000 267.590000 1186.000000 268.410000 ;
      RECT 1116.500000 267.590000 1156.500000 268.410000 ;
      RECT 1066.500000 267.590000 1108.500000 268.410000 ;
      RECT 1016.500000 267.590000 1058.500000 268.410000 ;
      RECT 966.500000 267.590000 1008.500000 268.410000 ;
      RECT 916.500000 267.590000 958.500000 268.410000 ;
      RECT 866.500000 267.590000 908.500000 268.410000 ;
      RECT 816.500000 267.590000 858.500000 268.410000 ;
      RECT 766.500000 267.590000 808.500000 268.410000 ;
      RECT 716.500000 267.590000 758.500000 268.410000 ;
      RECT 666.500000 267.590000 708.500000 268.410000 ;
      RECT 616.500000 267.590000 658.500000 268.410000 ;
      RECT 566.500000 267.590000 608.500000 268.410000 ;
      RECT 516.500000 267.590000 558.500000 268.410000 ;
      RECT 466.500000 267.590000 508.500000 268.410000 ;
      RECT 416.500000 267.590000 458.500000 268.410000 ;
      RECT 366.500000 267.590000 408.500000 268.410000 ;
      RECT 316.500000 267.590000 358.500000 268.410000 ;
      RECT 266.500000 267.590000 308.500000 268.410000 ;
      RECT 216.500000 267.590000 258.500000 268.410000 ;
      RECT 166.500000 267.590000 208.500000 268.410000 ;
      RECT 116.500000 267.590000 158.500000 268.410000 ;
      RECT 66.500000 267.590000 108.500000 268.410000 ;
      RECT 29.500000 267.590000 58.500000 268.410000 ;
      RECT 0.000000 267.590000 16.500000 268.410000 ;
      RECT 1169.500000 266.410000 1170.500000 267.590000 ;
      RECT 1116.500000 266.410000 1149.500000 267.590000 ;
      RECT 1107.500000 266.410000 1108.500000 267.590000 ;
      RECT 1066.500000 266.410000 1099.500000 267.590000 ;
      RECT 1057.500000 266.410000 1058.500000 267.590000 ;
      RECT 1016.500000 266.410000 1049.500000 267.590000 ;
      RECT 1007.500000 266.410000 1008.500000 267.590000 ;
      RECT 966.500000 266.410000 999.500000 267.590000 ;
      RECT 957.500000 266.410000 958.500000 267.590000 ;
      RECT 916.500000 266.410000 949.500000 267.590000 ;
      RECT 907.500000 266.410000 908.500000 267.590000 ;
      RECT 866.500000 266.410000 899.500000 267.590000 ;
      RECT 857.500000 266.410000 858.500000 267.590000 ;
      RECT 816.500000 266.410000 849.500000 267.590000 ;
      RECT 807.500000 266.410000 808.500000 267.590000 ;
      RECT 766.500000 266.410000 799.500000 267.590000 ;
      RECT 757.500000 266.410000 758.500000 267.590000 ;
      RECT 716.500000 266.410000 749.500000 267.590000 ;
      RECT 707.500000 266.410000 708.500000 267.590000 ;
      RECT 666.500000 266.410000 699.500000 267.590000 ;
      RECT 657.500000 266.410000 658.500000 267.590000 ;
      RECT 616.500000 266.410000 649.500000 267.590000 ;
      RECT 607.500000 266.410000 608.500000 267.590000 ;
      RECT 566.500000 266.410000 599.500000 267.590000 ;
      RECT 557.500000 266.410000 558.500000 267.590000 ;
      RECT 516.500000 266.410000 549.500000 267.590000 ;
      RECT 507.500000 266.410000 508.500000 267.590000 ;
      RECT 466.500000 266.410000 499.500000 267.590000 ;
      RECT 457.500000 266.410000 458.500000 267.590000 ;
      RECT 416.500000 266.410000 449.500000 267.590000 ;
      RECT 407.500000 266.410000 408.500000 267.590000 ;
      RECT 366.500000 266.410000 399.500000 267.590000 ;
      RECT 357.500000 266.410000 358.500000 267.590000 ;
      RECT 316.500000 266.410000 349.500000 267.590000 ;
      RECT 307.500000 266.410000 308.500000 267.590000 ;
      RECT 266.500000 266.410000 299.500000 267.590000 ;
      RECT 257.500000 266.410000 258.500000 267.590000 ;
      RECT 216.500000 266.410000 249.500000 267.590000 ;
      RECT 207.500000 266.410000 208.500000 267.590000 ;
      RECT 166.500000 266.410000 199.500000 267.590000 ;
      RECT 157.500000 266.410000 158.500000 267.590000 ;
      RECT 116.500000 266.410000 149.500000 267.590000 ;
      RECT 107.500000 266.410000 108.500000 267.590000 ;
      RECT 66.500000 266.410000 99.500000 267.590000 ;
      RECT 57.500000 266.410000 58.500000 267.590000 ;
      RECT 29.500000 266.410000 49.500000 267.590000 ;
      RECT 15.500000 266.410000 16.500000 267.590000 ;
      RECT 1157.500000 265.590000 1170.500000 266.410000 ;
      RECT 1107.500000 265.590000 1149.500000 266.410000 ;
      RECT 1057.500000 265.590000 1099.500000 266.410000 ;
      RECT 1007.500000 265.590000 1049.500000 266.410000 ;
      RECT 957.500000 265.590000 999.500000 266.410000 ;
      RECT 907.500000 265.590000 949.500000 266.410000 ;
      RECT 857.500000 265.590000 899.500000 266.410000 ;
      RECT 807.500000 265.590000 849.500000 266.410000 ;
      RECT 757.500000 265.590000 799.500000 266.410000 ;
      RECT 707.500000 265.590000 749.500000 266.410000 ;
      RECT 657.500000 265.590000 699.500000 266.410000 ;
      RECT 607.500000 265.590000 649.500000 266.410000 ;
      RECT 557.500000 265.590000 599.500000 266.410000 ;
      RECT 507.500000 265.590000 549.500000 266.410000 ;
      RECT 457.500000 265.590000 499.500000 266.410000 ;
      RECT 407.500000 265.590000 449.500000 266.410000 ;
      RECT 357.500000 265.590000 399.500000 266.410000 ;
      RECT 307.500000 265.590000 349.500000 266.410000 ;
      RECT 257.500000 265.590000 299.500000 266.410000 ;
      RECT 207.500000 265.590000 249.500000 266.410000 ;
      RECT 157.500000 265.590000 199.500000 266.410000 ;
      RECT 107.500000 265.590000 149.500000 266.410000 ;
      RECT 57.500000 265.590000 99.500000 266.410000 ;
      RECT 15.500000 265.590000 49.500000 266.410000 ;
      RECT 1183.500000 264.410000 1186.000000 267.590000 ;
      RECT 1169.500000 264.410000 1170.500000 265.590000 ;
      RECT 1116.500000 264.410000 1149.500000 265.590000 ;
      RECT 1107.500000 264.410000 1108.500000 265.590000 ;
      RECT 1066.500000 264.410000 1099.500000 265.590000 ;
      RECT 1057.500000 264.410000 1058.500000 265.590000 ;
      RECT 1016.500000 264.410000 1049.500000 265.590000 ;
      RECT 1007.500000 264.410000 1008.500000 265.590000 ;
      RECT 966.500000 264.410000 999.500000 265.590000 ;
      RECT 957.500000 264.410000 958.500000 265.590000 ;
      RECT 916.500000 264.410000 949.500000 265.590000 ;
      RECT 907.500000 264.410000 908.500000 265.590000 ;
      RECT 866.500000 264.410000 899.500000 265.590000 ;
      RECT 857.500000 264.410000 858.500000 265.590000 ;
      RECT 816.500000 264.410000 849.500000 265.590000 ;
      RECT 807.500000 264.410000 808.500000 265.590000 ;
      RECT 766.500000 264.410000 799.500000 265.590000 ;
      RECT 757.500000 264.410000 758.500000 265.590000 ;
      RECT 716.500000 264.410000 749.500000 265.590000 ;
      RECT 707.500000 264.410000 708.500000 265.590000 ;
      RECT 666.500000 264.410000 699.500000 265.590000 ;
      RECT 657.500000 264.410000 658.500000 265.590000 ;
      RECT 616.500000 264.410000 649.500000 265.590000 ;
      RECT 607.500000 264.410000 608.500000 265.590000 ;
      RECT 566.500000 264.410000 599.500000 265.590000 ;
      RECT 557.500000 264.410000 558.500000 265.590000 ;
      RECT 516.500000 264.410000 549.500000 265.590000 ;
      RECT 507.500000 264.410000 508.500000 265.590000 ;
      RECT 466.500000 264.410000 499.500000 265.590000 ;
      RECT 457.500000 264.410000 458.500000 265.590000 ;
      RECT 416.500000 264.410000 449.500000 265.590000 ;
      RECT 407.500000 264.410000 408.500000 265.590000 ;
      RECT 366.500000 264.410000 399.500000 265.590000 ;
      RECT 357.500000 264.410000 358.500000 265.590000 ;
      RECT 316.500000 264.410000 349.500000 265.590000 ;
      RECT 307.500000 264.410000 308.500000 265.590000 ;
      RECT 266.500000 264.410000 299.500000 265.590000 ;
      RECT 257.500000 264.410000 258.500000 265.590000 ;
      RECT 216.500000 264.410000 249.500000 265.590000 ;
      RECT 207.500000 264.410000 208.500000 265.590000 ;
      RECT 166.500000 264.410000 199.500000 265.590000 ;
      RECT 157.500000 264.410000 158.500000 265.590000 ;
      RECT 116.500000 264.410000 149.500000 265.590000 ;
      RECT 107.500000 264.410000 108.500000 265.590000 ;
      RECT 66.500000 264.410000 99.500000 265.590000 ;
      RECT 57.500000 264.410000 58.500000 265.590000 ;
      RECT 29.500000 264.410000 49.500000 265.590000 ;
      RECT 15.500000 264.410000 16.500000 265.590000 ;
      RECT 0.000000 264.410000 2.500000 267.590000 ;
      RECT 1169.500000 263.590000 1186.000000 264.410000 ;
      RECT 1116.500000 263.590000 1156.500000 264.410000 ;
      RECT 1066.500000 263.590000 1108.500000 264.410000 ;
      RECT 1016.500000 263.590000 1058.500000 264.410000 ;
      RECT 966.500000 263.590000 1008.500000 264.410000 ;
      RECT 916.500000 263.590000 958.500000 264.410000 ;
      RECT 866.500000 263.590000 908.500000 264.410000 ;
      RECT 816.500000 263.590000 858.500000 264.410000 ;
      RECT 766.500000 263.590000 808.500000 264.410000 ;
      RECT 716.500000 263.590000 758.500000 264.410000 ;
      RECT 666.500000 263.590000 708.500000 264.410000 ;
      RECT 616.500000 263.590000 658.500000 264.410000 ;
      RECT 566.500000 263.590000 608.500000 264.410000 ;
      RECT 516.500000 263.590000 558.500000 264.410000 ;
      RECT 466.500000 263.590000 508.500000 264.410000 ;
      RECT 416.500000 263.590000 458.500000 264.410000 ;
      RECT 366.500000 263.590000 408.500000 264.410000 ;
      RECT 316.500000 263.590000 358.500000 264.410000 ;
      RECT 266.500000 263.590000 308.500000 264.410000 ;
      RECT 216.500000 263.590000 258.500000 264.410000 ;
      RECT 166.500000 263.590000 208.500000 264.410000 ;
      RECT 116.500000 263.590000 158.500000 264.410000 ;
      RECT 66.500000 263.590000 108.500000 264.410000 ;
      RECT 29.500000 263.590000 58.500000 264.410000 ;
      RECT 0.000000 263.590000 16.500000 264.410000 ;
      RECT 1169.500000 262.410000 1170.500000 263.590000 ;
      RECT 1116.500000 262.410000 1149.500000 263.590000 ;
      RECT 1107.500000 262.410000 1108.500000 263.590000 ;
      RECT 1066.500000 262.410000 1099.500000 263.590000 ;
      RECT 1057.500000 262.410000 1058.500000 263.590000 ;
      RECT 1016.500000 262.410000 1049.500000 263.590000 ;
      RECT 1007.500000 262.410000 1008.500000 263.590000 ;
      RECT 966.500000 262.410000 999.500000 263.590000 ;
      RECT 957.500000 262.410000 958.500000 263.590000 ;
      RECT 916.500000 262.410000 949.500000 263.590000 ;
      RECT 907.500000 262.410000 908.500000 263.590000 ;
      RECT 866.500000 262.410000 899.500000 263.590000 ;
      RECT 857.500000 262.410000 858.500000 263.590000 ;
      RECT 816.500000 262.410000 849.500000 263.590000 ;
      RECT 807.500000 262.410000 808.500000 263.590000 ;
      RECT 766.500000 262.410000 799.500000 263.590000 ;
      RECT 757.500000 262.410000 758.500000 263.590000 ;
      RECT 716.500000 262.410000 749.500000 263.590000 ;
      RECT 707.500000 262.410000 708.500000 263.590000 ;
      RECT 666.500000 262.410000 699.500000 263.590000 ;
      RECT 657.500000 262.410000 658.500000 263.590000 ;
      RECT 616.500000 262.410000 649.500000 263.590000 ;
      RECT 607.500000 262.410000 608.500000 263.590000 ;
      RECT 566.500000 262.410000 599.500000 263.590000 ;
      RECT 557.500000 262.410000 558.500000 263.590000 ;
      RECT 516.500000 262.410000 549.500000 263.590000 ;
      RECT 507.500000 262.410000 508.500000 263.590000 ;
      RECT 466.500000 262.410000 499.500000 263.590000 ;
      RECT 457.500000 262.410000 458.500000 263.590000 ;
      RECT 416.500000 262.410000 449.500000 263.590000 ;
      RECT 407.500000 262.410000 408.500000 263.590000 ;
      RECT 366.500000 262.410000 399.500000 263.590000 ;
      RECT 357.500000 262.410000 358.500000 263.590000 ;
      RECT 316.500000 262.410000 349.500000 263.590000 ;
      RECT 307.500000 262.410000 308.500000 263.590000 ;
      RECT 266.500000 262.410000 299.500000 263.590000 ;
      RECT 257.500000 262.410000 258.500000 263.590000 ;
      RECT 216.500000 262.410000 249.500000 263.590000 ;
      RECT 207.500000 262.410000 208.500000 263.590000 ;
      RECT 166.500000 262.410000 199.500000 263.590000 ;
      RECT 157.500000 262.410000 158.500000 263.590000 ;
      RECT 116.500000 262.410000 149.500000 263.590000 ;
      RECT 107.500000 262.410000 108.500000 263.590000 ;
      RECT 66.500000 262.410000 99.500000 263.590000 ;
      RECT 57.500000 262.410000 58.500000 263.590000 ;
      RECT 29.500000 262.410000 49.500000 263.590000 ;
      RECT 15.500000 262.410000 16.500000 263.590000 ;
      RECT 1157.500000 261.590000 1170.500000 262.410000 ;
      RECT 1107.500000 261.590000 1149.500000 262.410000 ;
      RECT 1057.500000 261.590000 1099.500000 262.410000 ;
      RECT 1007.500000 261.590000 1049.500000 262.410000 ;
      RECT 957.500000 261.590000 999.500000 262.410000 ;
      RECT 907.500000 261.590000 949.500000 262.410000 ;
      RECT 857.500000 261.590000 899.500000 262.410000 ;
      RECT 807.500000 261.590000 849.500000 262.410000 ;
      RECT 757.500000 261.590000 799.500000 262.410000 ;
      RECT 707.500000 261.590000 749.500000 262.410000 ;
      RECT 657.500000 261.590000 699.500000 262.410000 ;
      RECT 607.500000 261.590000 649.500000 262.410000 ;
      RECT 557.500000 261.590000 599.500000 262.410000 ;
      RECT 507.500000 261.590000 549.500000 262.410000 ;
      RECT 457.500000 261.590000 499.500000 262.410000 ;
      RECT 407.500000 261.590000 449.500000 262.410000 ;
      RECT 357.500000 261.590000 399.500000 262.410000 ;
      RECT 307.500000 261.590000 349.500000 262.410000 ;
      RECT 257.500000 261.590000 299.500000 262.410000 ;
      RECT 207.500000 261.590000 249.500000 262.410000 ;
      RECT 157.500000 261.590000 199.500000 262.410000 ;
      RECT 107.500000 261.590000 149.500000 262.410000 ;
      RECT 57.500000 261.590000 99.500000 262.410000 ;
      RECT 15.500000 261.590000 49.500000 262.410000 ;
      RECT 1183.500000 260.410000 1186.000000 263.590000 ;
      RECT 1169.500000 260.410000 1170.500000 261.590000 ;
      RECT 1116.500000 260.410000 1149.500000 261.590000 ;
      RECT 1107.500000 260.410000 1108.500000 261.590000 ;
      RECT 1066.500000 260.410000 1099.500000 261.590000 ;
      RECT 1057.500000 260.410000 1058.500000 261.590000 ;
      RECT 1016.500000 260.410000 1049.500000 261.590000 ;
      RECT 1007.500000 260.410000 1008.500000 261.590000 ;
      RECT 966.500000 260.410000 999.500000 261.590000 ;
      RECT 957.500000 260.410000 958.500000 261.590000 ;
      RECT 916.500000 260.410000 949.500000 261.590000 ;
      RECT 907.500000 260.410000 908.500000 261.590000 ;
      RECT 866.500000 260.410000 899.500000 261.590000 ;
      RECT 857.500000 260.410000 858.500000 261.590000 ;
      RECT 816.500000 260.410000 849.500000 261.590000 ;
      RECT 807.500000 260.410000 808.500000 261.590000 ;
      RECT 766.500000 260.410000 799.500000 261.590000 ;
      RECT 757.500000 260.410000 758.500000 261.590000 ;
      RECT 716.500000 260.410000 749.500000 261.590000 ;
      RECT 707.500000 260.410000 708.500000 261.590000 ;
      RECT 666.500000 260.410000 699.500000 261.590000 ;
      RECT 657.500000 260.410000 658.500000 261.590000 ;
      RECT 616.500000 260.410000 649.500000 261.590000 ;
      RECT 607.500000 260.410000 608.500000 261.590000 ;
      RECT 566.500000 260.410000 599.500000 261.590000 ;
      RECT 557.500000 260.410000 558.500000 261.590000 ;
      RECT 516.500000 260.410000 549.500000 261.590000 ;
      RECT 507.500000 260.410000 508.500000 261.590000 ;
      RECT 466.500000 260.410000 499.500000 261.590000 ;
      RECT 457.500000 260.410000 458.500000 261.590000 ;
      RECT 416.500000 260.410000 449.500000 261.590000 ;
      RECT 407.500000 260.410000 408.500000 261.590000 ;
      RECT 366.500000 260.410000 399.500000 261.590000 ;
      RECT 357.500000 260.410000 358.500000 261.590000 ;
      RECT 316.500000 260.410000 349.500000 261.590000 ;
      RECT 307.500000 260.410000 308.500000 261.590000 ;
      RECT 266.500000 260.410000 299.500000 261.590000 ;
      RECT 257.500000 260.410000 258.500000 261.590000 ;
      RECT 216.500000 260.410000 249.500000 261.590000 ;
      RECT 207.500000 260.410000 208.500000 261.590000 ;
      RECT 166.500000 260.410000 199.500000 261.590000 ;
      RECT 157.500000 260.410000 158.500000 261.590000 ;
      RECT 116.500000 260.410000 149.500000 261.590000 ;
      RECT 107.500000 260.410000 108.500000 261.590000 ;
      RECT 66.500000 260.410000 99.500000 261.590000 ;
      RECT 57.500000 260.410000 58.500000 261.590000 ;
      RECT 29.500000 260.410000 49.500000 261.590000 ;
      RECT 15.500000 260.410000 16.500000 261.590000 ;
      RECT 0.000000 260.410000 2.500000 263.590000 ;
      RECT 1169.500000 259.590000 1186.000000 260.410000 ;
      RECT 1116.500000 259.590000 1156.500000 260.410000 ;
      RECT 1169.500000 258.410000 1170.500000 259.590000 ;
      RECT 1116.500000 258.410000 1149.500000 259.590000 ;
      RECT 1066.500000 258.410000 1108.500000 260.410000 ;
      RECT 1016.500000 258.410000 1058.500000 260.410000 ;
      RECT 966.500000 258.410000 1008.500000 260.410000 ;
      RECT 916.500000 258.410000 958.500000 260.410000 ;
      RECT 866.500000 258.410000 908.500000 260.410000 ;
      RECT 816.500000 258.410000 858.500000 260.410000 ;
      RECT 766.500000 258.410000 808.500000 260.410000 ;
      RECT 716.500000 258.410000 758.500000 260.410000 ;
      RECT 666.500000 258.410000 708.500000 260.410000 ;
      RECT 616.500000 258.410000 658.500000 260.410000 ;
      RECT 566.500000 258.410000 608.500000 260.410000 ;
      RECT 516.500000 258.410000 558.500000 260.410000 ;
      RECT 466.500000 258.410000 508.500000 260.410000 ;
      RECT 416.500000 258.410000 458.500000 260.410000 ;
      RECT 366.500000 258.410000 408.500000 260.410000 ;
      RECT 316.500000 258.410000 358.500000 260.410000 ;
      RECT 266.500000 258.410000 308.500000 260.410000 ;
      RECT 216.500000 258.410000 258.500000 260.410000 ;
      RECT 166.500000 258.410000 208.500000 260.410000 ;
      RECT 116.500000 258.410000 158.500000 260.410000 ;
      RECT 66.500000 258.410000 108.500000 260.410000 ;
      RECT 29.500000 258.410000 58.500000 260.410000 ;
      RECT 0.000000 258.410000 16.500000 260.410000 ;
      RECT 1157.500000 257.590000 1170.500000 258.410000 ;
      RECT 1183.500000 256.410000 1186.000000 259.590000 ;
      RECT 1169.500000 256.410000 1170.500000 257.590000 ;
      RECT 0.000000 256.410000 1149.500000 258.410000 ;
      RECT 1169.500000 255.590000 1186.000000 256.410000 ;
      RECT 1169.500000 254.410000 1170.500000 255.590000 ;
      RECT 0.000000 254.410000 1156.500000 256.410000 ;
      RECT 0.000000 253.590000 1170.500000 254.410000 ;
      RECT 1183.500000 252.410000 1186.000000 255.590000 ;
      RECT 1169.500000 252.410000 1170.500000 253.590000 ;
      RECT 1169.500000 251.590000 1186.000000 252.410000 ;
      RECT 1169.500000 250.410000 1170.500000 251.590000 ;
      RECT 0.000000 250.410000 1156.500000 253.590000 ;
      RECT 0.000000 249.590000 1170.500000 250.410000 ;
      RECT 1183.500000 248.410000 1186.000000 251.590000 ;
      RECT 1169.500000 248.410000 1170.500000 249.590000 ;
      RECT 1169.500000 247.590000 1186.000000 248.410000 ;
      RECT 1169.500000 246.410000 1170.500000 247.590000 ;
      RECT 0.000000 246.410000 1156.500000 249.590000 ;
      RECT 0.000000 245.590000 1170.500000 246.410000 ;
      RECT 1183.500000 244.410000 1186.000000 247.590000 ;
      RECT 1169.500000 244.410000 1170.500000 245.590000 ;
      RECT 1169.500000 243.590000 1186.000000 244.410000 ;
      RECT 1169.500000 242.410000 1170.500000 243.590000 ;
      RECT 0.000000 242.410000 1156.500000 245.590000 ;
      RECT 0.000000 241.590000 1170.500000 242.410000 ;
      RECT 1183.500000 240.410000 1186.000000 243.590000 ;
      RECT 1169.500000 240.410000 1170.500000 241.590000 ;
      RECT 1169.500000 239.590000 1186.000000 240.410000 ;
      RECT 1169.500000 238.410000 1170.500000 239.590000 ;
      RECT 0.000000 238.410000 1156.500000 241.590000 ;
      RECT 0.000000 237.590000 1170.500000 238.410000 ;
      RECT 1183.500000 236.410000 1186.000000 239.590000 ;
      RECT 1169.500000 236.410000 1170.500000 237.590000 ;
      RECT 1169.500000 235.590000 1186.000000 236.410000 ;
      RECT 1169.500000 234.410000 1170.500000 235.590000 ;
      RECT 0.000000 234.410000 1156.500000 237.590000 ;
      RECT 0.000000 233.590000 1170.500000 234.410000 ;
      RECT 1183.500000 232.410000 1186.000000 235.590000 ;
      RECT 1169.500000 232.410000 1170.500000 233.590000 ;
      RECT 1169.500000 231.590000 1186.000000 232.410000 ;
      RECT 1169.500000 230.410000 1170.500000 231.590000 ;
      RECT 0.000000 230.410000 1156.500000 233.590000 ;
      RECT 0.000000 229.590000 1170.500000 230.410000 ;
      RECT 1183.500000 228.410000 1186.000000 231.590000 ;
      RECT 1169.500000 228.410000 1170.500000 229.590000 ;
      RECT 1169.500000 227.590000 1186.000000 228.410000 ;
      RECT 1169.500000 226.410000 1170.500000 227.590000 ;
      RECT 0.000000 226.410000 1156.500000 229.590000 ;
      RECT 0.000000 225.590000 1170.500000 226.410000 ;
      RECT 1183.500000 224.410000 1186.000000 227.590000 ;
      RECT 1169.500000 224.410000 1170.500000 225.590000 ;
      RECT 1169.500000 223.590000 1186.000000 224.410000 ;
      RECT 1169.500000 222.410000 1170.500000 223.590000 ;
      RECT 0.000000 222.410000 1156.500000 225.590000 ;
      RECT 0.000000 221.590000 1170.500000 222.410000 ;
      RECT 1183.500000 220.410000 1186.000000 223.590000 ;
      RECT 1169.500000 220.410000 1170.500000 221.590000 ;
      RECT 1169.500000 219.590000 1186.000000 220.410000 ;
      RECT 1169.500000 218.410000 1170.500000 219.590000 ;
      RECT 0.000000 218.410000 1156.500000 221.590000 ;
      RECT 0.000000 217.590000 1170.500000 218.410000 ;
      RECT 1183.500000 216.410000 1186.000000 219.590000 ;
      RECT 1169.500000 216.410000 1170.500000 217.590000 ;
      RECT 1169.500000 215.590000 1186.000000 216.410000 ;
      RECT 1169.500000 214.410000 1170.500000 215.590000 ;
      RECT 0.000000 214.410000 1156.500000 217.590000 ;
      RECT 0.000000 213.590000 1170.500000 214.410000 ;
      RECT 1183.500000 212.410000 1186.000000 215.590000 ;
      RECT 1169.500000 212.410000 1170.500000 213.590000 ;
      RECT 1169.500000 211.590000 1186.000000 212.410000 ;
      RECT 1169.500000 210.410000 1170.500000 211.590000 ;
      RECT 0.000000 210.410000 1156.500000 213.590000 ;
      RECT 0.000000 209.590000 1170.500000 210.410000 ;
      RECT 1183.500000 208.410000 1186.000000 211.590000 ;
      RECT 1169.500000 208.410000 1170.500000 209.590000 ;
      RECT 1169.500000 207.590000 1186.000000 208.410000 ;
      RECT 1169.500000 206.410000 1170.500000 207.590000 ;
      RECT 0.000000 206.410000 1156.500000 209.590000 ;
      RECT 0.000000 205.590000 1170.500000 206.410000 ;
      RECT 1183.500000 204.410000 1186.000000 207.590000 ;
      RECT 1169.500000 204.410000 1170.500000 205.590000 ;
      RECT 1169.500000 203.590000 1186.000000 204.410000 ;
      RECT 1169.500000 202.410000 1170.500000 203.590000 ;
      RECT 0.000000 202.410000 1156.500000 205.590000 ;
      RECT 0.000000 201.590000 1170.500000 202.410000 ;
      RECT 1183.500000 200.410000 1186.000000 203.590000 ;
      RECT 1169.500000 200.410000 1170.500000 201.590000 ;
      RECT 1169.500000 199.590000 1186.000000 200.410000 ;
      RECT 1169.500000 198.410000 1170.500000 199.590000 ;
      RECT 0.000000 198.410000 1156.500000 201.590000 ;
      RECT 0.000000 197.590000 1170.500000 198.410000 ;
      RECT 1183.500000 196.410000 1186.000000 199.590000 ;
      RECT 1169.500000 196.410000 1170.500000 197.590000 ;
      RECT 1169.500000 195.590000 1186.000000 196.410000 ;
      RECT 1169.500000 194.410000 1170.500000 195.590000 ;
      RECT 0.000000 194.410000 1156.500000 197.590000 ;
      RECT 0.000000 193.590000 1170.500000 194.410000 ;
      RECT 1183.500000 192.410000 1186.000000 195.590000 ;
      RECT 1169.500000 192.410000 1170.500000 193.590000 ;
      RECT 1169.500000 191.590000 1186.000000 192.410000 ;
      RECT 1169.500000 190.410000 1170.500000 191.590000 ;
      RECT 0.000000 190.410000 1156.500000 193.590000 ;
      RECT 0.000000 189.590000 1170.500000 190.410000 ;
      RECT 1183.500000 188.410000 1186.000000 191.590000 ;
      RECT 1169.500000 188.410000 1170.500000 189.590000 ;
      RECT 1169.500000 187.590000 1186.000000 188.410000 ;
      RECT 1169.500000 186.410000 1170.500000 187.590000 ;
      RECT 0.000000 186.410000 1156.500000 189.590000 ;
      RECT 0.000000 185.590000 1170.500000 186.410000 ;
      RECT 1183.500000 184.410000 1186.000000 187.590000 ;
      RECT 1169.500000 184.410000 1170.500000 185.590000 ;
      RECT 1169.500000 183.590000 1186.000000 184.410000 ;
      RECT 1169.500000 182.410000 1170.500000 183.590000 ;
      RECT 0.000000 182.410000 1156.500000 185.590000 ;
      RECT 0.000000 181.590000 1170.500000 182.410000 ;
      RECT 1183.500000 180.410000 1186.000000 183.590000 ;
      RECT 1169.500000 180.410000 1170.500000 181.590000 ;
      RECT 1169.500000 179.590000 1186.000000 180.410000 ;
      RECT 1169.500000 178.410000 1170.500000 179.590000 ;
      RECT 0.000000 178.410000 1156.500000 181.590000 ;
      RECT 0.000000 177.590000 1170.500000 178.410000 ;
      RECT 1183.500000 176.410000 1186.000000 179.590000 ;
      RECT 1169.500000 176.410000 1170.500000 177.590000 ;
      RECT 1169.500000 175.590000 1186.000000 176.410000 ;
      RECT 1169.500000 174.410000 1170.500000 175.590000 ;
      RECT 0.000000 174.410000 1156.500000 177.590000 ;
      RECT 0.000000 173.590000 1170.500000 174.410000 ;
      RECT 1183.500000 172.410000 1186.000000 175.590000 ;
      RECT 1169.500000 172.410000 1170.500000 173.590000 ;
      RECT 1169.500000 171.590000 1186.000000 172.410000 ;
      RECT 1169.500000 170.410000 1170.500000 171.590000 ;
      RECT 0.000000 170.410000 1156.500000 173.590000 ;
      RECT 0.000000 169.590000 1170.500000 170.410000 ;
      RECT 1183.500000 168.410000 1186.000000 171.590000 ;
      RECT 1169.500000 168.410000 1170.500000 169.590000 ;
      RECT 1169.500000 167.590000 1186.000000 168.410000 ;
      RECT 1169.500000 166.410000 1170.500000 167.590000 ;
      RECT 0.000000 166.410000 1156.500000 169.590000 ;
      RECT 0.000000 165.590000 1170.500000 166.410000 ;
      RECT 1183.500000 164.410000 1186.000000 167.590000 ;
      RECT 1169.500000 164.410000 1170.500000 165.590000 ;
      RECT 1169.500000 163.590000 1186.000000 164.410000 ;
      RECT 1169.500000 162.410000 1170.500000 163.590000 ;
      RECT 0.000000 162.410000 1156.500000 165.590000 ;
      RECT 0.000000 161.590000 1170.500000 162.410000 ;
      RECT 1183.500000 160.410000 1186.000000 163.590000 ;
      RECT 1169.500000 160.410000 1170.500000 161.590000 ;
      RECT 1169.500000 159.590000 1186.000000 160.410000 ;
      RECT 1169.500000 158.410000 1170.500000 159.590000 ;
      RECT 0.000000 158.410000 1156.500000 161.590000 ;
      RECT 0.000000 157.590000 1170.500000 158.410000 ;
      RECT 1183.500000 156.410000 1186.000000 159.590000 ;
      RECT 1169.500000 156.410000 1170.500000 157.590000 ;
      RECT 1169.500000 155.590000 1186.000000 156.410000 ;
      RECT 1169.500000 154.410000 1170.500000 155.590000 ;
      RECT 0.000000 154.410000 1156.500000 157.590000 ;
      RECT 0.000000 153.590000 1170.500000 154.410000 ;
      RECT 1183.500000 152.410000 1186.000000 155.590000 ;
      RECT 1169.500000 152.410000 1170.500000 153.590000 ;
      RECT 1169.500000 151.590000 1186.000000 152.410000 ;
      RECT 1169.500000 150.410000 1170.500000 151.590000 ;
      RECT 0.000000 150.410000 1156.500000 153.590000 ;
      RECT 0.000000 149.590000 1170.500000 150.410000 ;
      RECT 1183.500000 148.410000 1186.000000 151.590000 ;
      RECT 1169.500000 148.410000 1170.500000 149.590000 ;
      RECT 1169.500000 147.590000 1186.000000 148.410000 ;
      RECT 1169.500000 146.410000 1170.500000 147.590000 ;
      RECT 0.000000 146.410000 1156.500000 149.590000 ;
      RECT 0.000000 145.590000 1170.500000 146.410000 ;
      RECT 1183.500000 144.410000 1186.000000 147.590000 ;
      RECT 1169.500000 144.410000 1170.500000 145.590000 ;
      RECT 1169.500000 143.590000 1186.000000 144.410000 ;
      RECT 1169.500000 142.410000 1170.500000 143.590000 ;
      RECT 0.000000 142.410000 1156.500000 145.590000 ;
      RECT 0.000000 141.590000 1170.500000 142.410000 ;
      RECT 1183.500000 140.410000 1186.000000 143.590000 ;
      RECT 1169.500000 140.410000 1170.500000 141.590000 ;
      RECT 1169.500000 139.590000 1186.000000 140.410000 ;
      RECT 1169.500000 138.410000 1170.500000 139.590000 ;
      RECT 0.000000 138.410000 1156.500000 141.590000 ;
      RECT 0.000000 137.590000 1170.500000 138.410000 ;
      RECT 1183.500000 136.410000 1186.000000 139.590000 ;
      RECT 1169.500000 136.410000 1170.500000 137.590000 ;
      RECT 1169.500000 135.590000 1186.000000 136.410000 ;
      RECT 0.000000 135.590000 1156.500000 137.590000 ;
      RECT 1169.500000 134.410000 1170.500000 135.590000 ;
      RECT 1157.500000 133.590000 1170.500000 134.410000 ;
      RECT 1183.500000 132.410000 1186.000000 135.590000 ;
      RECT 1169.500000 132.410000 1170.500000 133.590000 ;
      RECT 0.000000 132.410000 1149.500000 135.590000 ;
      RECT 1169.500000 131.590000 1186.000000 132.410000 ;
      RECT 1169.500000 130.410000 1170.500000 131.590000 ;
      RECT 0.000000 130.410000 1156.500000 132.410000 ;
      RECT 0.000000 129.590000 1170.500000 130.410000 ;
      RECT 1183.500000 128.410000 1186.000000 131.590000 ;
      RECT 1169.500000 128.410000 1170.500000 129.590000 ;
      RECT 1169.500000 127.590000 1186.000000 128.410000 ;
      RECT 1169.500000 126.410000 1170.500000 127.590000 ;
      RECT 0.000000 126.410000 1156.500000 129.590000 ;
      RECT 0.000000 125.590000 1170.500000 126.410000 ;
      RECT 1183.500000 124.410000 1186.000000 127.590000 ;
      RECT 1169.500000 124.410000 1170.500000 125.590000 ;
      RECT 1169.500000 123.590000 1186.000000 124.410000 ;
      RECT 1169.500000 122.410000 1170.500000 123.590000 ;
      RECT 0.000000 122.410000 1156.500000 125.590000 ;
      RECT 0.000000 121.590000 1170.500000 122.410000 ;
      RECT 1183.500000 120.410000 1186.000000 123.590000 ;
      RECT 1169.500000 120.410000 1170.500000 121.590000 ;
      RECT 1169.500000 119.590000 1186.000000 120.410000 ;
      RECT 1169.500000 118.410000 1170.500000 119.590000 ;
      RECT 0.000000 118.410000 1156.500000 121.590000 ;
      RECT 0.000000 117.590000 1170.500000 118.410000 ;
      RECT 1183.500000 116.410000 1186.000000 119.590000 ;
      RECT 1169.500000 116.410000 1170.500000 117.590000 ;
      RECT 1169.500000 115.590000 1186.000000 116.410000 ;
      RECT 1169.500000 114.410000 1170.500000 115.590000 ;
      RECT 0.000000 114.410000 1156.500000 117.590000 ;
      RECT 0.000000 113.590000 1170.500000 114.410000 ;
      RECT 1183.500000 112.410000 1186.000000 115.590000 ;
      RECT 1169.500000 112.410000 1170.500000 113.590000 ;
      RECT 1169.500000 111.590000 1186.000000 112.410000 ;
      RECT 1169.500000 110.410000 1170.500000 111.590000 ;
      RECT 0.000000 110.410000 1156.500000 113.590000 ;
      RECT 0.000000 109.590000 1170.500000 110.410000 ;
      RECT 1183.500000 108.410000 1186.000000 111.590000 ;
      RECT 1169.500000 108.410000 1170.500000 109.590000 ;
      RECT 1169.500000 107.590000 1186.000000 108.410000 ;
      RECT 1169.500000 106.410000 1170.500000 107.590000 ;
      RECT 0.000000 106.410000 1156.500000 109.590000 ;
      RECT 0.000000 105.590000 1170.500000 106.410000 ;
      RECT 1183.500000 104.410000 1186.000000 107.590000 ;
      RECT 1169.500000 104.410000 1170.500000 105.590000 ;
      RECT 1169.500000 103.590000 1186.000000 104.410000 ;
      RECT 1169.500000 102.410000 1170.500000 103.590000 ;
      RECT 0.000000 102.410000 1156.500000 105.590000 ;
      RECT 0.000000 101.590000 1170.500000 102.410000 ;
      RECT 1183.500000 100.410000 1186.000000 103.590000 ;
      RECT 1169.500000 100.410000 1170.500000 101.590000 ;
      RECT 1169.500000 99.590000 1186.000000 100.410000 ;
      RECT 1169.500000 98.410000 1170.500000 99.590000 ;
      RECT 0.000000 98.410000 1156.500000 101.590000 ;
      RECT 0.000000 97.590000 1170.500000 98.410000 ;
      RECT 1183.500000 96.410000 1186.000000 99.590000 ;
      RECT 1169.500000 96.410000 1170.500000 97.590000 ;
      RECT 1169.500000 95.590000 1186.000000 96.410000 ;
      RECT 1169.500000 94.410000 1170.500000 95.590000 ;
      RECT 0.000000 94.410000 1156.500000 97.590000 ;
      RECT 0.000000 93.590000 1170.500000 94.410000 ;
      RECT 1183.500000 92.410000 1186.000000 95.590000 ;
      RECT 1169.500000 92.410000 1170.500000 93.590000 ;
      RECT 1169.500000 91.590000 1186.000000 92.410000 ;
      RECT 1169.500000 90.410000 1170.500000 91.590000 ;
      RECT 0.000000 90.410000 1156.500000 93.590000 ;
      RECT 0.000000 89.590000 1170.500000 90.410000 ;
      RECT 1183.500000 88.410000 1186.000000 91.590000 ;
      RECT 1169.500000 88.410000 1170.500000 89.590000 ;
      RECT 1169.500000 87.590000 1186.000000 88.410000 ;
      RECT 1169.500000 86.410000 1170.500000 87.590000 ;
      RECT 0.000000 86.410000 1156.500000 89.590000 ;
      RECT 0.000000 85.590000 1170.500000 86.410000 ;
      RECT 1183.500000 84.410000 1186.000000 87.590000 ;
      RECT 1169.500000 84.410000 1170.500000 85.590000 ;
      RECT 1169.500000 83.590000 1186.000000 84.410000 ;
      RECT 1169.500000 82.410000 1170.500000 83.590000 ;
      RECT 0.000000 82.410000 1156.500000 85.590000 ;
      RECT 0.000000 81.590000 1170.500000 82.410000 ;
      RECT 1183.500000 80.410000 1186.000000 83.590000 ;
      RECT 1169.500000 80.410000 1170.500000 81.590000 ;
      RECT 1169.500000 79.590000 1186.000000 80.410000 ;
      RECT 1169.500000 78.410000 1170.500000 79.590000 ;
      RECT 0.000000 78.410000 1156.500000 81.590000 ;
      RECT 0.000000 77.590000 1170.500000 78.410000 ;
      RECT 1183.500000 76.410000 1186.000000 79.590000 ;
      RECT 1169.500000 76.410000 1170.500000 77.590000 ;
      RECT 1169.500000 75.590000 1186.000000 76.410000 ;
      RECT 1169.500000 74.410000 1170.500000 75.590000 ;
      RECT 0.000000 74.410000 1156.500000 77.590000 ;
      RECT 0.000000 73.590000 1170.500000 74.410000 ;
      RECT 1183.500000 72.410000 1186.000000 75.590000 ;
      RECT 1169.500000 72.410000 1170.500000 73.590000 ;
      RECT 1169.500000 71.590000 1186.000000 72.410000 ;
      RECT 1169.500000 70.410000 1170.500000 71.590000 ;
      RECT 0.000000 70.410000 1156.500000 73.590000 ;
      RECT 0.000000 69.590000 1170.500000 70.410000 ;
      RECT 1183.500000 68.410000 1186.000000 71.590000 ;
      RECT 1169.500000 68.410000 1170.500000 69.590000 ;
      RECT 1169.500000 67.590000 1186.000000 68.410000 ;
      RECT 1169.500000 66.410000 1170.500000 67.590000 ;
      RECT 0.000000 66.410000 1156.500000 69.590000 ;
      RECT 0.000000 65.590000 1170.500000 66.410000 ;
      RECT 1183.500000 64.410000 1186.000000 67.590000 ;
      RECT 1169.500000 64.410000 1170.500000 65.590000 ;
      RECT 1169.500000 63.590000 1186.000000 64.410000 ;
      RECT 1169.500000 62.410000 1170.500000 63.590000 ;
      RECT 0.000000 62.410000 1156.500000 65.590000 ;
      RECT 0.000000 61.590000 1170.500000 62.410000 ;
      RECT 1183.500000 60.410000 1186.000000 63.590000 ;
      RECT 1169.500000 60.410000 1170.500000 61.590000 ;
      RECT 1169.500000 59.590000 1186.000000 60.410000 ;
      RECT 1169.500000 58.410000 1170.500000 59.590000 ;
      RECT 0.000000 58.410000 1156.500000 61.590000 ;
      RECT 0.000000 57.590000 1170.500000 58.410000 ;
      RECT 1183.500000 56.410000 1186.000000 59.590000 ;
      RECT 1169.500000 56.410000 1170.500000 57.590000 ;
      RECT 1169.500000 55.590000 1186.000000 56.410000 ;
      RECT 1169.500000 54.410000 1170.500000 55.590000 ;
      RECT 0.000000 54.410000 1156.500000 57.590000 ;
      RECT 0.000000 53.590000 1170.500000 54.410000 ;
      RECT 1183.500000 52.410000 1186.000000 55.590000 ;
      RECT 1169.500000 52.410000 1170.500000 53.590000 ;
      RECT 1169.500000 51.590000 1186.000000 52.410000 ;
      RECT 1169.500000 50.410000 1170.500000 51.590000 ;
      RECT 0.000000 50.410000 1156.500000 53.590000 ;
      RECT 0.000000 49.590000 1170.500000 50.410000 ;
      RECT 1183.500000 48.410000 1186.000000 51.590000 ;
      RECT 1169.500000 48.410000 1170.500000 49.590000 ;
      RECT 1169.500000 47.590000 1186.000000 48.410000 ;
      RECT 1169.500000 46.410000 1170.500000 47.590000 ;
      RECT 0.000000 46.410000 1156.500000 49.590000 ;
      RECT 0.000000 45.590000 1170.500000 46.410000 ;
      RECT 1183.500000 44.410000 1186.000000 47.590000 ;
      RECT 1169.500000 44.410000 1170.500000 45.590000 ;
      RECT 1169.500000 43.590000 1186.000000 44.410000 ;
      RECT 1169.500000 42.410000 1170.500000 43.590000 ;
      RECT 0.000000 42.410000 1156.500000 45.590000 ;
      RECT 0.000000 41.590000 1170.500000 42.410000 ;
      RECT 1183.500000 40.410000 1186.000000 43.590000 ;
      RECT 1169.500000 40.410000 1170.500000 41.590000 ;
      RECT 1169.500000 39.590000 1186.000000 40.410000 ;
      RECT 1169.500000 38.410000 1170.500000 39.590000 ;
      RECT 0.000000 38.410000 1156.500000 41.590000 ;
      RECT 0.000000 37.590000 1170.500000 38.410000 ;
      RECT 1183.500000 36.410000 1186.000000 39.590000 ;
      RECT 1169.500000 36.410000 1170.500000 37.590000 ;
      RECT 1169.500000 35.590000 1186.000000 36.410000 ;
      RECT 1169.500000 34.410000 1170.500000 35.590000 ;
      RECT 0.000000 34.410000 1156.500000 37.590000 ;
      RECT 0.000000 33.590000 1170.500000 34.410000 ;
      RECT 1183.500000 32.410000 1186.000000 35.590000 ;
      RECT 1169.500000 32.410000 1170.500000 33.590000 ;
      RECT 1169.500000 31.590000 1186.000000 32.410000 ;
      RECT 1169.500000 30.410000 1170.500000 31.590000 ;
      RECT 0.000000 30.410000 1156.500000 33.590000 ;
      RECT 0.000000 29.590000 1170.500000 30.410000 ;
      RECT 1183.500000 28.410000 1186.000000 31.590000 ;
      RECT 1169.500000 28.410000 1170.500000 29.590000 ;
      RECT 1169.500000 27.590000 1186.000000 28.410000 ;
      RECT 1169.500000 26.410000 1170.500000 27.590000 ;
      RECT 0.000000 26.410000 1156.500000 29.590000 ;
      RECT 0.000000 25.590000 1170.500000 26.410000 ;
      RECT 1183.500000 24.410000 1186.000000 27.590000 ;
      RECT 1169.500000 24.410000 1170.500000 25.590000 ;
      RECT 1169.500000 23.590000 1186.000000 24.410000 ;
      RECT 1169.500000 22.410000 1170.500000 23.590000 ;
      RECT 0.000000 22.410000 1156.500000 25.590000 ;
      RECT 0.000000 21.590000 1170.500000 22.410000 ;
      RECT 1183.500000 20.410000 1186.000000 23.590000 ;
      RECT 1169.500000 20.410000 1170.500000 21.590000 ;
      RECT 1169.500000 19.590000 1186.000000 20.410000 ;
      RECT 1169.500000 18.410000 1170.500000 19.590000 ;
      RECT 0.000000 18.410000 1156.500000 21.590000 ;
      RECT 0.000000 17.590000 1170.500000 18.410000 ;
      RECT 1183.500000 16.410000 1186.000000 19.590000 ;
      RECT 1166.500000 16.410000 1170.500000 17.590000 ;
      RECT 1166.500000 15.590000 1186.000000 16.410000 ;
      RECT 1166.500000 14.410000 1170.500000 15.590000 ;
      RECT 0.000000 14.410000 1158.500000 17.590000 ;
      RECT 0.000000 13.590000 1170.500000 14.410000 ;
      RECT 1183.500000 12.410000 1186.000000 15.590000 ;
      RECT 1166.500000 12.410000 1170.500000 13.590000 ;
      RECT 1166.500000 11.590000 1186.000000 12.410000 ;
      RECT 1166.500000 10.410000 1170.500000 11.590000 ;
      RECT 0.000000 10.410000 1158.500000 13.590000 ;
      RECT 0.000000 9.590000 1170.500000 10.410000 ;
      RECT 1183.500000 8.410000 1186.000000 11.590000 ;
      RECT 1166.500000 8.410000 1170.500000 9.590000 ;
      RECT 1166.500000 7.590000 1186.000000 8.410000 ;
      RECT 1116.500000 7.590000 1158.500000 9.590000 ;
      RECT 1066.500000 7.590000 1108.500000 9.590000 ;
      RECT 1016.500000 7.590000 1058.500000 9.590000 ;
      RECT 966.500000 7.590000 1008.500000 9.590000 ;
      RECT 916.500000 7.590000 958.500000 9.590000 ;
      RECT 866.500000 7.590000 908.500000 9.590000 ;
      RECT 816.500000 7.590000 858.500000 9.590000 ;
      RECT 766.500000 7.590000 808.500000 9.590000 ;
      RECT 716.500000 7.590000 758.500000 9.590000 ;
      RECT 666.500000 7.590000 708.500000 9.590000 ;
      RECT 616.500000 7.590000 658.500000 9.590000 ;
      RECT 566.500000 7.590000 608.500000 9.590000 ;
      RECT 516.500000 7.590000 558.500000 9.590000 ;
      RECT 466.500000 7.590000 508.500000 9.590000 ;
      RECT 416.500000 7.590000 458.500000 9.590000 ;
      RECT 366.500000 7.590000 408.500000 9.590000 ;
      RECT 316.500000 7.590000 358.500000 9.590000 ;
      RECT 266.500000 7.590000 308.500000 9.590000 ;
      RECT 216.500000 7.590000 258.500000 9.590000 ;
      RECT 166.500000 7.590000 208.500000 9.590000 ;
      RECT 116.500000 7.590000 158.500000 9.590000 ;
      RECT 66.500000 7.590000 108.500000 9.590000 ;
      RECT 0.000000 7.590000 58.500000 9.590000 ;
      RECT 1166.500000 6.410000 1170.500000 7.590000 ;
      RECT 1157.500000 6.410000 1158.500000 7.590000 ;
      RECT 1116.500000 6.410000 1149.500000 7.590000 ;
      RECT 1107.500000 6.410000 1108.500000 7.590000 ;
      RECT 1066.500000 6.410000 1099.500000 7.590000 ;
      RECT 1057.500000 6.410000 1058.500000 7.590000 ;
      RECT 1016.500000 6.410000 1049.500000 7.590000 ;
      RECT 1007.500000 6.410000 1008.500000 7.590000 ;
      RECT 966.500000 6.410000 999.500000 7.590000 ;
      RECT 957.500000 6.410000 958.500000 7.590000 ;
      RECT 916.500000 6.410000 949.500000 7.590000 ;
      RECT 907.500000 6.410000 908.500000 7.590000 ;
      RECT 866.500000 6.410000 899.500000 7.590000 ;
      RECT 857.500000 6.410000 858.500000 7.590000 ;
      RECT 816.500000 6.410000 849.500000 7.590000 ;
      RECT 807.500000 6.410000 808.500000 7.590000 ;
      RECT 766.500000 6.410000 799.500000 7.590000 ;
      RECT 757.500000 6.410000 758.500000 7.590000 ;
      RECT 716.500000 6.410000 749.500000 7.590000 ;
      RECT 707.500000 6.410000 708.500000 7.590000 ;
      RECT 666.500000 6.410000 699.500000 7.590000 ;
      RECT 657.500000 6.410000 658.500000 7.590000 ;
      RECT 616.500000 6.410000 649.500000 7.590000 ;
      RECT 607.500000 6.410000 608.500000 7.590000 ;
      RECT 566.500000 6.410000 599.500000 7.590000 ;
      RECT 557.500000 6.410000 558.500000 7.590000 ;
      RECT 516.500000 6.410000 549.500000 7.590000 ;
      RECT 507.500000 6.410000 508.500000 7.590000 ;
      RECT 466.500000 6.410000 499.500000 7.590000 ;
      RECT 457.500000 6.410000 458.500000 7.590000 ;
      RECT 416.500000 6.410000 449.500000 7.590000 ;
      RECT 407.500000 6.410000 408.500000 7.590000 ;
      RECT 366.500000 6.410000 399.500000 7.590000 ;
      RECT 357.500000 6.410000 358.500000 7.590000 ;
      RECT 316.500000 6.410000 349.500000 7.590000 ;
      RECT 307.500000 6.410000 308.500000 7.590000 ;
      RECT 266.500000 6.410000 299.500000 7.590000 ;
      RECT 257.500000 6.410000 258.500000 7.590000 ;
      RECT 216.500000 6.410000 249.500000 7.590000 ;
      RECT 207.500000 6.410000 208.500000 7.590000 ;
      RECT 166.500000 6.410000 199.500000 7.590000 ;
      RECT 157.500000 6.410000 158.500000 7.590000 ;
      RECT 116.500000 6.410000 149.500000 7.590000 ;
      RECT 107.500000 6.410000 108.500000 7.590000 ;
      RECT 66.500000 6.410000 99.500000 7.590000 ;
      RECT 57.500000 6.410000 58.500000 7.590000 ;
      RECT 1157.500000 5.590000 1170.500000 6.410000 ;
      RECT 1107.500000 5.590000 1149.500000 6.410000 ;
      RECT 1057.500000 5.590000 1099.500000 6.410000 ;
      RECT 1007.500000 5.590000 1049.500000 6.410000 ;
      RECT 957.500000 5.590000 999.500000 6.410000 ;
      RECT 907.500000 5.590000 949.500000 6.410000 ;
      RECT 857.500000 5.590000 899.500000 6.410000 ;
      RECT 807.500000 5.590000 849.500000 6.410000 ;
      RECT 757.500000 5.590000 799.500000 6.410000 ;
      RECT 707.500000 5.590000 749.500000 6.410000 ;
      RECT 657.500000 5.590000 699.500000 6.410000 ;
      RECT 607.500000 5.590000 649.500000 6.410000 ;
      RECT 557.500000 5.590000 599.500000 6.410000 ;
      RECT 507.500000 5.590000 549.500000 6.410000 ;
      RECT 457.500000 5.590000 499.500000 6.410000 ;
      RECT 407.500000 5.590000 449.500000 6.410000 ;
      RECT 357.500000 5.590000 399.500000 6.410000 ;
      RECT 307.500000 5.590000 349.500000 6.410000 ;
      RECT 257.500000 5.590000 299.500000 6.410000 ;
      RECT 207.500000 5.590000 249.500000 6.410000 ;
      RECT 157.500000 5.590000 199.500000 6.410000 ;
      RECT 107.500000 5.590000 149.500000 6.410000 ;
      RECT 57.500000 5.590000 99.500000 6.410000 ;
      RECT 1183.500000 4.410000 1186.000000 7.590000 ;
      RECT 1166.500000 4.410000 1170.500000 5.590000 ;
      RECT 1157.500000 4.410000 1158.500000 5.590000 ;
      RECT 1116.500000 4.410000 1149.500000 5.590000 ;
      RECT 1107.500000 4.410000 1108.500000 5.590000 ;
      RECT 1066.500000 4.410000 1099.500000 5.590000 ;
      RECT 1057.500000 4.410000 1058.500000 5.590000 ;
      RECT 1016.500000 4.410000 1049.500000 5.590000 ;
      RECT 1007.500000 4.410000 1008.500000 5.590000 ;
      RECT 966.500000 4.410000 999.500000 5.590000 ;
      RECT 957.500000 4.410000 958.500000 5.590000 ;
      RECT 916.500000 4.410000 949.500000 5.590000 ;
      RECT 907.500000 4.410000 908.500000 5.590000 ;
      RECT 866.500000 4.410000 899.500000 5.590000 ;
      RECT 857.500000 4.410000 858.500000 5.590000 ;
      RECT 816.500000 4.410000 849.500000 5.590000 ;
      RECT 807.500000 4.410000 808.500000 5.590000 ;
      RECT 766.500000 4.410000 799.500000 5.590000 ;
      RECT 757.500000 4.410000 758.500000 5.590000 ;
      RECT 716.500000 4.410000 749.500000 5.590000 ;
      RECT 707.500000 4.410000 708.500000 5.590000 ;
      RECT 666.500000 4.410000 699.500000 5.590000 ;
      RECT 657.500000 4.410000 658.500000 5.590000 ;
      RECT 616.500000 4.410000 649.500000 5.590000 ;
      RECT 607.500000 4.410000 608.500000 5.590000 ;
      RECT 566.500000 4.410000 599.500000 5.590000 ;
      RECT 557.500000 4.410000 558.500000 5.590000 ;
      RECT 516.500000 4.410000 549.500000 5.590000 ;
      RECT 507.500000 4.410000 508.500000 5.590000 ;
      RECT 466.500000 4.410000 499.500000 5.590000 ;
      RECT 457.500000 4.410000 458.500000 5.590000 ;
      RECT 416.500000 4.410000 449.500000 5.590000 ;
      RECT 407.500000 4.410000 408.500000 5.590000 ;
      RECT 366.500000 4.410000 399.500000 5.590000 ;
      RECT 357.500000 4.410000 358.500000 5.590000 ;
      RECT 316.500000 4.410000 349.500000 5.590000 ;
      RECT 307.500000 4.410000 308.500000 5.590000 ;
      RECT 266.500000 4.410000 299.500000 5.590000 ;
      RECT 257.500000 4.410000 258.500000 5.590000 ;
      RECT 216.500000 4.410000 249.500000 5.590000 ;
      RECT 207.500000 4.410000 208.500000 5.590000 ;
      RECT 166.500000 4.410000 199.500000 5.590000 ;
      RECT 157.500000 4.410000 158.500000 5.590000 ;
      RECT 116.500000 4.410000 149.500000 5.590000 ;
      RECT 107.500000 4.410000 108.500000 5.590000 ;
      RECT 66.500000 4.410000 99.500000 5.590000 ;
      RECT 57.500000 4.410000 58.500000 5.590000 ;
      RECT 15.500000 4.410000 49.500000 7.590000 ;
      RECT 0.000000 4.410000 2.500000 7.590000 ;
      RECT 1116.500000 3.590000 1158.500000 4.410000 ;
      RECT 1066.500000 3.590000 1108.500000 4.410000 ;
      RECT 1016.500000 3.590000 1058.500000 4.410000 ;
      RECT 966.500000 3.590000 1008.500000 4.410000 ;
      RECT 916.500000 3.590000 958.500000 4.410000 ;
      RECT 866.500000 3.590000 908.500000 4.410000 ;
      RECT 816.500000 3.590000 858.500000 4.410000 ;
      RECT 766.500000 3.590000 808.500000 4.410000 ;
      RECT 716.500000 3.590000 758.500000 4.410000 ;
      RECT 666.500000 3.590000 708.500000 4.410000 ;
      RECT 616.500000 3.590000 658.500000 4.410000 ;
      RECT 566.500000 3.590000 608.500000 4.410000 ;
      RECT 516.500000 3.590000 558.500000 4.410000 ;
      RECT 466.500000 3.590000 508.500000 4.410000 ;
      RECT 416.500000 3.590000 458.500000 4.410000 ;
      RECT 366.500000 3.590000 408.500000 4.410000 ;
      RECT 316.500000 3.590000 358.500000 4.410000 ;
      RECT 266.500000 3.590000 308.500000 4.410000 ;
      RECT 216.500000 3.590000 258.500000 4.410000 ;
      RECT 166.500000 3.590000 208.500000 4.410000 ;
      RECT 116.500000 3.590000 158.500000 4.410000 ;
      RECT 66.500000 3.590000 108.500000 4.410000 ;
      RECT 0.000000 3.590000 58.500000 4.410000 ;
      RECT 1166.500000 2.410000 1186.000000 4.410000 ;
      RECT 1157.500000 2.410000 1158.500000 3.590000 ;
      RECT 1116.500000 2.410000 1149.500000 3.590000 ;
      RECT 1107.500000 2.410000 1108.500000 3.590000 ;
      RECT 1066.500000 2.410000 1099.500000 3.590000 ;
      RECT 1057.500000 2.410000 1058.500000 3.590000 ;
      RECT 1016.500000 2.410000 1049.500000 3.590000 ;
      RECT 1007.500000 2.410000 1008.500000 3.590000 ;
      RECT 966.500000 2.410000 999.500000 3.590000 ;
      RECT 957.500000 2.410000 958.500000 3.590000 ;
      RECT 916.500000 2.410000 949.500000 3.590000 ;
      RECT 907.500000 2.410000 908.500000 3.590000 ;
      RECT 866.500000 2.410000 899.500000 3.590000 ;
      RECT 857.500000 2.410000 858.500000 3.590000 ;
      RECT 816.500000 2.410000 849.500000 3.590000 ;
      RECT 807.500000 2.410000 808.500000 3.590000 ;
      RECT 766.500000 2.410000 799.500000 3.590000 ;
      RECT 757.500000 2.410000 758.500000 3.590000 ;
      RECT 716.500000 2.410000 749.500000 3.590000 ;
      RECT 707.500000 2.410000 708.500000 3.590000 ;
      RECT 666.500000 2.410000 699.500000 3.590000 ;
      RECT 657.500000 2.410000 658.500000 3.590000 ;
      RECT 616.500000 2.410000 649.500000 3.590000 ;
      RECT 607.500000 2.410000 608.500000 3.590000 ;
      RECT 566.500000 2.410000 599.500000 3.590000 ;
      RECT 557.500000 2.410000 558.500000 3.590000 ;
      RECT 516.500000 2.410000 549.500000 3.590000 ;
      RECT 507.500000 2.410000 508.500000 3.590000 ;
      RECT 466.500000 2.410000 499.500000 3.590000 ;
      RECT 457.500000 2.410000 458.500000 3.590000 ;
      RECT 416.500000 2.410000 449.500000 3.590000 ;
      RECT 407.500000 2.410000 408.500000 3.590000 ;
      RECT 366.500000 2.410000 399.500000 3.590000 ;
      RECT 357.500000 2.410000 358.500000 3.590000 ;
      RECT 316.500000 2.410000 349.500000 3.590000 ;
      RECT 307.500000 2.410000 308.500000 3.590000 ;
      RECT 266.500000 2.410000 299.500000 3.590000 ;
      RECT 257.500000 2.410000 258.500000 3.590000 ;
      RECT 216.500000 2.410000 249.500000 3.590000 ;
      RECT 207.500000 2.410000 208.500000 3.590000 ;
      RECT 166.500000 2.410000 199.500000 3.590000 ;
      RECT 157.500000 2.410000 158.500000 3.590000 ;
      RECT 116.500000 2.410000 149.500000 3.590000 ;
      RECT 107.500000 2.410000 108.500000 3.590000 ;
      RECT 66.500000 2.410000 99.500000 3.590000 ;
      RECT 57.500000 2.410000 58.500000 3.590000 ;
      RECT 1157.500000 0.410000 1186.000000 2.410000 ;
      RECT 1107.500000 0.410000 1149.500000 2.410000 ;
      RECT 1057.500000 0.410000 1099.500000 2.410000 ;
      RECT 1007.500000 0.410000 1049.500000 2.410000 ;
      RECT 957.500000 0.410000 999.500000 2.410000 ;
      RECT 907.500000 0.410000 949.500000 2.410000 ;
      RECT 857.500000 0.410000 899.500000 2.410000 ;
      RECT 807.500000 0.410000 849.500000 2.410000 ;
      RECT 757.500000 0.410000 799.500000 2.410000 ;
      RECT 707.500000 0.410000 749.500000 2.410000 ;
      RECT 657.500000 0.410000 699.500000 2.410000 ;
      RECT 607.500000 0.410000 649.500000 2.410000 ;
      RECT 557.500000 0.410000 599.500000 2.410000 ;
      RECT 507.500000 0.410000 549.500000 2.410000 ;
      RECT 457.500000 0.410000 499.500000 2.410000 ;
      RECT 407.500000 0.410000 449.500000 2.410000 ;
      RECT 357.500000 0.410000 399.500000 2.410000 ;
      RECT 307.500000 0.410000 349.500000 2.410000 ;
      RECT 257.500000 0.410000 299.500000 2.410000 ;
      RECT 207.500000 0.410000 249.500000 2.410000 ;
      RECT 157.500000 0.410000 199.500000 2.410000 ;
      RECT 107.500000 0.410000 149.500000 2.410000 ;
      RECT 57.500000 0.410000 99.500000 2.410000 ;
      RECT 0.000000 0.410000 49.500000 3.590000 ;
      RECT 0.000000 0.000000 1186.000000 0.410000 ;
  END
END MCU

END LIBRARY
